
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"c9",x"01"),
     1 => (x"cf",x"03",x"87",x"cc"),
     2 => (x"87",x"fd",x"00",x"87"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"36",x"27",x"4f",x"00"),
     5 => (x"4f",x"00",x"00",x"00"),
     6 => (x"0e",x"1e",x"18",x"0e"),
     7 => (x"00",x"00",x"44",x"27"),
     8 => (x"48",x"26",x"0f",x"00"),
     9 => (x"08",x"26",x"80",x"ff"),
    10 => (x"c0",x"c0",x"c2",x"4f"),
    11 => (x"05",x"38",x"27",x"4e"),
    12 => (x"00",x"0f",x"00",x"00"),
    13 => (x"f0",x"c1",x"87",x"fd"),
    14 => (x"43",x"27",x"4e",x"c0"),
    15 => (x"0f",x"00",x"00",x"00"),
    16 => (x"4f",x"87",x"fd",x"00"),
    17 => (x"0e",x"1e",x"18",x"0e"),
    18 => (x"80",x"ff",x"48",x"26"),
    19 => (x"1e",x"4f",x"08",x"26"),
    20 => (x"ff",x"1e",x"1e",x"72"),
    21 => (x"48",x"6a",x"4a",x"c0"),
    22 => (x"c4",x"98",x"c0",x"c4"),
    23 => (x"02",x"6e",x"58",x"a6"),
    24 => (x"cc",x"87",x"f3",x"ff"),
    25 => (x"66",x"cc",x"7a",x"66"),
    26 => (x"4a",x"26",x"26",x"48"),
    27 => (x"5e",x"0e",x"4f",x"26"),
    28 => (x"5d",x"5c",x"5b",x"5a"),
    29 => (x"4b",x"66",x"d4",x"0e"),
    30 => (x"4c",x"13",x"4d",x"c0"),
    31 => (x"c0",x"02",x"9c",x"74"),
    32 => (x"4a",x"74",x"87",x"d6"),
    33 => (x"4f",x"27",x"1e",x"72"),
    34 => (x"0f",x"00",x"00",x"00"),
    35 => (x"85",x"c1",x"86",x"c4"),
    36 => (x"9c",x"74",x"4c",x"13"),
    37 => (x"87",x"ea",x"ff",x"05"),
    38 => (x"4d",x"26",x"48",x"75"),
    39 => (x"4b",x"26",x"4c",x"26"),
    40 => (x"4f",x"26",x"4a",x"26"),
    41 => (x"5b",x"5a",x"5e",x"0e"),
    42 => (x"c8",x"0e",x"5d",x"5c"),
    43 => (x"66",x"e0",x"c0",x"8e"),
    44 => (x"4c",x"66",x"dc",x"4d"),
    45 => (x"00",x"16",x"48",x"27"),
    46 => (x"49",x"76",x"4b",x"00"),
    47 => (x"00",x"0e",x"90",x"27"),
    48 => (x"a6",x"c4",x"79",x"00"),
    49 => (x"c0",x"79",x"c0",x"49"),
    50 => (x"c0",x"03",x"ac",x"b7"),
    51 => (x"ed",x"c0",x"87",x"cd"),
    52 => (x"00",x"4f",x"27",x"1e"),
    53 => (x"c4",x"0f",x"00",x"00"),
    54 => (x"74",x"8c",x"0c",x"86"),
    55 => (x"c6",x"c0",x"05",x"9c"),
    56 => (x"53",x"f0",x"c0",x"87"),
    57 => (x"74",x"87",x"f6",x"c0"),
    58 => (x"f0",x"c0",x"02",x"9c"),
    59 => (x"72",x"49",x"74",x"87"),
    60 => (x"66",x"e8",x"c0",x"1e"),
    61 => (x"04",x"da",x"27",x"4a"),
    62 => (x"26",x"0f",x"00",x"00"),
    63 => (x"72",x"4a",x"71",x"4a"),
    64 => (x"12",x"82",x"6e",x"4a"),
    65 => (x"72",x"49",x"74",x"53"),
    66 => (x"66",x"e8",x"c0",x"1e"),
    67 => (x"04",x"da",x"27",x"4a"),
    68 => (x"26",x"0f",x"00",x"00"),
    69 => (x"74",x"4c",x"70",x"4a"),
    70 => (x"d0",x"ff",x"05",x"9c"),
    71 => (x"16",x"48",x"27",x"87"),
    72 => (x"ab",x"b7",x"00",x"00"),
    73 => (x"87",x"d8",x"c0",x"02"),
    74 => (x"6b",x"97",x"8b",x"c1"),
    75 => (x"48",x"66",x"c4",x"55"),
    76 => (x"a6",x"c8",x"80",x"c1"),
    77 => (x"16",x"48",x"27",x"58"),
    78 => (x"ab",x"b7",x"00",x"00"),
    79 => (x"87",x"e8",x"ff",x"05"),
    80 => (x"66",x"c4",x"55",x"c0"),
    81 => (x"26",x"86",x"c8",x"48"),
    82 => (x"26",x"4c",x"26",x"4d"),
    83 => (x"26",x"4a",x"26",x"4b"),
    84 => (x"5a",x"5e",x"0e",x"4f"),
    85 => (x"0e",x"5d",x"5c",x"5b"),
    86 => (x"76",x"4c",x"c0",x"1e"),
    87 => (x"dc",x"79",x"c0",x"49"),
    88 => (x"66",x"d8",x"4b",x"a6"),
    89 => (x"48",x"66",x"d8",x"4a"),
    90 => (x"a6",x"dc",x"80",x"c1"),
    91 => (x"c1",x"4d",x"12",x"58"),
    92 => (x"c0",x"c0",x"c0",x"c0"),
    93 => (x"b7",x"c0",x"c4",x"95"),
    94 => (x"9d",x"75",x"4d",x"95"),
    95 => (x"87",x"d2",x"c4",x"02"),
    96 => (x"d7",x"c3",x"02",x"6e"),
    97 => (x"c0",x"49",x"76",x"87"),
    98 => (x"c1",x"4a",x"75",x"79"),
    99 => (x"c2",x"02",x"ad",x"e3"),
   100 => (x"e4",x"c1",x"87",x"dd"),
   101 => (x"d8",x"c0",x"02",x"aa"),
   102 => (x"aa",x"ec",x"c1",x"87"),
   103 => (x"87",x"c8",x"c2",x"02"),
   104 => (x"02",x"aa",x"f3",x"c1"),
   105 => (x"c1",x"87",x"e8",x"c1"),
   106 => (x"c0",x"02",x"aa",x"f8"),
   107 => (x"d3",x"c2",x"87",x"f2"),
   108 => (x"27",x"1e",x"ca",x"87"),
   109 => (x"00",x"00",x"16",x"98"),
   110 => (x"73",x"83",x"c4",x"1e"),
   111 => (x"6a",x"8a",x"c4",x"4a"),
   112 => (x"00",x"a4",x"27",x"1e"),
   113 => (x"cc",x"0f",x"00",x"00"),
   114 => (x"74",x"4a",x"70",x"86"),
   115 => (x"27",x"84",x"72",x"4c"),
   116 => (x"00",x"00",x"16",x"98"),
   117 => (x"00",x"6e",x"27",x"1e"),
   118 => (x"c4",x"0f",x"00",x"00"),
   119 => (x"87",x"d4",x"c2",x"86"),
   120 => (x"98",x"27",x"1e",x"d0"),
   121 => (x"1e",x"00",x"00",x"16"),
   122 => (x"4a",x"73",x"83",x"c4"),
   123 => (x"1e",x"6a",x"8a",x"c4"),
   124 => (x"00",x"00",x"a4",x"27"),
   125 => (x"86",x"cc",x"0f",x"00"),
   126 => (x"4c",x"74",x"4a",x"70"),
   127 => (x"98",x"27",x"84",x"72"),
   128 => (x"1e",x"00",x"00",x"16"),
   129 => (x"00",x"00",x"6e",x"27"),
   130 => (x"86",x"c4",x"0f",x"00"),
   131 => (x"c4",x"87",x"e5",x"c1"),
   132 => (x"c4",x"4a",x"73",x"83"),
   133 => (x"27",x"1e",x"6a",x"8a"),
   134 => (x"00",x"00",x"00",x"6e"),
   135 => (x"70",x"86",x"c4",x"0f"),
   136 => (x"72",x"4c",x"74",x"4a"),
   137 => (x"87",x"cc",x"c1",x"84"),
   138 => (x"79",x"c1",x"49",x"76"),
   139 => (x"c4",x"87",x"c5",x"c1"),
   140 => (x"c4",x"4a",x"73",x"83"),
   141 => (x"27",x"1e",x"6a",x"8a"),
   142 => (x"00",x"00",x"00",x"4f"),
   143 => (x"c1",x"86",x"c4",x"0f"),
   144 => (x"87",x"f0",x"c0",x"84"),
   145 => (x"27",x"1e",x"e5",x"c0"),
   146 => (x"00",x"00",x"00",x"4f"),
   147 => (x"75",x"86",x"c4",x"0f"),
   148 => (x"00",x"4f",x"27",x"1e"),
   149 => (x"c4",x"0f",x"00",x"00"),
   150 => (x"87",x"d8",x"c0",x"86"),
   151 => (x"05",x"ad",x"e5",x"c0"),
   152 => (x"76",x"87",x"c7",x"c0"),
   153 => (x"c0",x"79",x"c1",x"49"),
   154 => (x"1e",x"75",x"87",x"ca"),
   155 => (x"00",x"00",x"4f",x"27"),
   156 => (x"86",x"c4",x"0f",x"00"),
   157 => (x"d8",x"4a",x"66",x"d8"),
   158 => (x"80",x"c1",x"48",x"66"),
   159 => (x"12",x"58",x"a6",x"dc"),
   160 => (x"c0",x"c0",x"c1",x"4d"),
   161 => (x"c4",x"95",x"c0",x"c0"),
   162 => (x"4d",x"95",x"b7",x"c0"),
   163 => (x"fb",x"05",x"9d",x"75"),
   164 => (x"48",x"74",x"87",x"ee"),
   165 => (x"26",x"4d",x"26",x"26"),
   166 => (x"26",x"4b",x"26",x"4c"),
   167 => (x"0e",x"4f",x"26",x"4a"),
   168 => (x"0e",x"5b",x"5a",x"5e"),
   169 => (x"cc",x"4b",x"66",x"d0"),
   170 => (x"66",x"cc",x"7b",x"66"),
   171 => (x"04",x"c6",x"27",x"1e"),
   172 => (x"c4",x"0f",x"00",x"00"),
   173 => (x"72",x"4a",x"70",x"86"),
   174 => (x"c2",x"c0",x"05",x"9a"),
   175 => (x"cc",x"7b",x"c3",x"87"),
   176 => (x"66",x"cc",x"4a",x"66"),
   177 => (x"a9",x"b7",x"c0",x"49"),
   178 => (x"87",x"df",x"c0",x"02"),
   179 => (x"02",x"aa",x"b7",x"c1"),
   180 => (x"c2",x"87",x"dd",x"c0"),
   181 => (x"c0",x"02",x"aa",x"b7"),
   182 => (x"b7",x"c3",x"87",x"ef"),
   183 => (x"ef",x"c0",x"02",x"aa"),
   184 => (x"aa",x"b7",x"c4",x"87"),
   185 => (x"87",x"e6",x"c0",x"02"),
   186 => (x"c0",x"87",x"e5",x"c0"),
   187 => (x"87",x"e0",x"c0",x"7b"),
   188 => (x"00",x"16",x"c0",x"27"),
   189 => (x"c1",x"49",x"bf",x"00"),
   190 => (x"06",x"a9",x"b7",x"e4"),
   191 => (x"c0",x"87",x"c5",x"c0"),
   192 => (x"87",x"cc",x"c0",x"7b"),
   193 => (x"c7",x"c0",x"7b",x"c3"),
   194 => (x"c0",x"7b",x"c1",x"87"),
   195 => (x"7b",x"c2",x"87",x"c2"),
   196 => (x"4a",x"26",x"4b",x"26"),
   197 => (x"72",x"1e",x"4f",x"26"),
   198 => (x"4a",x"66",x"c8",x"1e"),
   199 => (x"66",x"cc",x"82",x"c2"),
   200 => (x"d0",x"80",x"72",x"48"),
   201 => (x"79",x"70",x"49",x"66"),
   202 => (x"4f",x"26",x"4a",x"26"),
   203 => (x"5b",x"5a",x"5e",x"0e"),
   204 => (x"dc",x"0e",x"5d",x"5c"),
   205 => (x"85",x"c5",x"4d",x"66"),
   206 => (x"92",x"c4",x"4a",x"75"),
   207 => (x"66",x"d4",x"4a",x"72"),
   208 => (x"66",x"e0",x"c0",x"82"),
   209 => (x"c4",x"4b",x"72",x"7a"),
   210 => (x"c1",x"7b",x"6a",x"83"),
   211 => (x"7a",x"75",x"82",x"f8"),
   212 => (x"4a",x"75",x"4c",x"75"),
   213 => (x"b7",x"72",x"82",x"c1"),
   214 => (x"e1",x"c0",x"01",x"ad"),
   215 => (x"c3",x"4b",x"75",x"87"),
   216 => (x"4b",x"73",x"93",x"c8"),
   217 => (x"74",x"83",x"66",x"d8"),
   218 => (x"72",x"92",x"c4",x"4a"),
   219 => (x"75",x"82",x"73",x"4a"),
   220 => (x"75",x"84",x"c1",x"7a"),
   221 => (x"72",x"82",x"c1",x"4a"),
   222 => (x"ff",x"06",x"ac",x"b7"),
   223 => (x"4c",x"75",x"87",x"df"),
   224 => (x"74",x"94",x"c8",x"c3"),
   225 => (x"84",x"66",x"d8",x"4c"),
   226 => (x"92",x"c4",x"4a",x"75"),
   227 => (x"83",x"72",x"4b",x"74"),
   228 => (x"48",x"6b",x"8b",x"c4"),
   229 => (x"7b",x"70",x"80",x"c1"),
   230 => (x"72",x"4b",x"66",x"d4"),
   231 => (x"e0",x"fe",x"c0",x"83"),
   232 => (x"74",x"4a",x"72",x"84"),
   233 => (x"27",x"7a",x"6b",x"82"),
   234 => (x"00",x"00",x"16",x"c0"),
   235 => (x"26",x"79",x"c5",x"49"),
   236 => (x"26",x"4c",x"26",x"4d"),
   237 => (x"26",x"4a",x"26",x"4b"),
   238 => (x"5a",x"5e",x"0e",x"4f"),
   239 => (x"97",x"0e",x"5c",x"5b"),
   240 => (x"74",x"4c",x"66",x"d0"),
   241 => (x"c0",x"c0",x"c1",x"4b"),
   242 => (x"c4",x"93",x"c0",x"c0"),
   243 => (x"4b",x"93",x"b7",x"c0"),
   244 => (x"4a",x"66",x"d4",x"97"),
   245 => (x"c0",x"c0",x"c0",x"c1"),
   246 => (x"c0",x"c4",x"92",x"c0"),
   247 => (x"72",x"4a",x"92",x"b7"),
   248 => (x"c0",x"02",x"ab",x"b7"),
   249 => (x"48",x"c0",x"87",x"c5"),
   250 => (x"27",x"87",x"ca",x"c0"),
   251 => (x"00",x"00",x"16",x"c8"),
   252 => (x"c1",x"51",x"74",x"49"),
   253 => (x"26",x"4c",x"26",x"48"),
   254 => (x"26",x"4a",x"26",x"4b"),
   255 => (x"5a",x"5e",x"0e",x"4f"),
   256 => (x"1e",x"0e",x"5c",x"5b"),
   257 => (x"c2",x"4c",x"6e",x"97"),
   258 => (x"4a",x"66",x"d8",x"4b"),
   259 => (x"82",x"73",x"82",x"c1"),
   260 => (x"c1",x"4a",x"6a",x"97"),
   261 => (x"c0",x"c0",x"c0",x"c0"),
   262 => (x"b7",x"c0",x"c4",x"92"),
   263 => (x"1e",x"72",x"4a",x"92"),
   264 => (x"73",x"4a",x"66",x"d8"),
   265 => (x"4a",x"6a",x"97",x"82"),
   266 => (x"c0",x"c0",x"c0",x"c1"),
   267 => (x"c0",x"c4",x"92",x"c0"),
   268 => (x"72",x"4a",x"92",x"b7"),
   269 => (x"03",x"b9",x"27",x"1e"),
   270 => (x"c8",x"0f",x"00",x"00"),
   271 => (x"72",x"4a",x"70",x"86"),
   272 => (x"c5",x"c0",x"05",x"9a"),
   273 => (x"4c",x"c1",x"c1",x"87"),
   274 => (x"b7",x"c2",x"83",x"c1"),
   275 => (x"f8",x"fe",x"06",x"ab"),
   276 => (x"c1",x"4a",x"74",x"87"),
   277 => (x"c0",x"c0",x"c0",x"c0"),
   278 => (x"b7",x"c0",x"c4",x"92"),
   279 => (x"d7",x"c1",x"4a",x"92"),
   280 => (x"c0",x"04",x"aa",x"b7"),
   281 => (x"4a",x"74",x"87",x"d7"),
   282 => (x"c0",x"c0",x"c0",x"c1"),
   283 => (x"c0",x"c4",x"92",x"c0"),
   284 => (x"c1",x"4a",x"92",x"b7"),
   285 => (x"03",x"aa",x"b7",x"da"),
   286 => (x"c7",x"87",x"c2",x"c0"),
   287 => (x"c1",x"4a",x"74",x"4b"),
   288 => (x"c0",x"c0",x"c0",x"c0"),
   289 => (x"b7",x"c0",x"c4",x"92"),
   290 => (x"d2",x"c1",x"4a",x"92"),
   291 => (x"c0",x"05",x"aa",x"b7"),
   292 => (x"48",x"c1",x"87",x"c5"),
   293 => (x"d4",x"87",x"e6",x"c0"),
   294 => (x"66",x"d8",x"4a",x"66"),
   295 => (x"05",x"24",x"27",x"49"),
   296 => (x"70",x"0f",x"00",x"00"),
   297 => (x"aa",x"b7",x"c0",x"4a"),
   298 => (x"87",x"cf",x"c0",x"06"),
   299 => (x"80",x"c7",x"48",x"73"),
   300 => (x"00",x"16",x"c4",x"27"),
   301 => (x"48",x"c1",x"58",x"00"),
   302 => (x"c0",x"87",x"c2",x"c0"),
   303 => (x"4c",x"26",x"26",x"48"),
   304 => (x"4a",x"26",x"4b",x"26"),
   305 => (x"c4",x"1e",x"4f",x"26"),
   306 => (x"b7",x"c2",x"49",x"66"),
   307 => (x"c5",x"c0",x"05",x"a9"),
   308 => (x"c0",x"48",x"c1",x"87"),
   309 => (x"48",x"c0",x"87",x"c2"),
   310 => (x"73",x"1e",x"4f",x"26"),
   311 => (x"02",x"9a",x"72",x"1e"),
   312 => (x"48",x"c0",x"87",x"d9"),
   313 => (x"a9",x"72",x"4b",x"c1"),
   314 => (x"83",x"73",x"82",x"01"),
   315 => (x"a9",x"72",x"87",x"f8"),
   316 => (x"80",x"73",x"89",x"03"),
   317 => (x"2b",x"2a",x"c1",x"07"),
   318 => (x"26",x"87",x"f3",x"05"),
   319 => (x"1e",x"4f",x"26",x"4b"),
   320 => (x"4d",x"c0",x"1e",x"75"),
   321 => (x"ff",x"04",x"a1",x"71"),
   322 => (x"bd",x"81",x"c1",x"b9"),
   323 => (x"04",x"a2",x"72",x"07"),
   324 => (x"82",x"c1",x"ba",x"ff"),
   325 => (x"87",x"c2",x"07",x"bd"),
   326 => (x"ff",x"05",x"9d",x"75"),
   327 => (x"07",x"80",x"c1",x"b8"),
   328 => (x"4f",x"26",x"4d",x"25"),
   329 => (x"11",x"48",x"12",x"1e"),
   330 => (x"88",x"87",x"c4",x"02"),
   331 => (x"26",x"87",x"f6",x"02"),
   332 => (x"c8",x"ff",x"1e",x"4f"),
   333 => (x"4f",x"26",x"48",x"bf"),
   334 => (x"5b",x"5a",x"5e",x"0e"),
   335 => (x"d0",x"0e",x"5d",x"5c"),
   336 => (x"4c",x"66",x"c4",x"8e"),
   337 => (x"00",x"16",x"bc",x"27"),
   338 => (x"c0",x"27",x"49",x"00"),
   339 => (x"79",x"00",x"00",x"3e"),
   340 => (x"00",x"16",x"b8",x"27"),
   341 => (x"f0",x"27",x"49",x"00"),
   342 => (x"79",x"00",x"00",x"3e"),
   343 => (x"00",x"3e",x"f0",x"27"),
   344 => (x"c0",x"27",x"49",x"00"),
   345 => (x"79",x"00",x"00",x"3e"),
   346 => (x"00",x"3e",x"f4",x"27"),
   347 => (x"79",x"c0",x"49",x"00"),
   348 => (x"00",x"3e",x"f8",x"27"),
   349 => (x"79",x"c2",x"49",x"00"),
   350 => (x"00",x"3e",x"fc",x"27"),
   351 => (x"e8",x"c0",x"49",x"00"),
   352 => (x"3f",x"00",x"27",x"79"),
   353 => (x"27",x"49",x"00",x"00"),
   354 => (x"00",x"00",x"10",x"1a"),
   355 => (x"20",x"1e",x"72",x"48"),
   356 => (x"20",x"41",x"20",x"41"),
   357 => (x"20",x"41",x"20",x"41"),
   358 => (x"20",x"41",x"20",x"41"),
   359 => (x"10",x"51",x"10",x"41"),
   360 => (x"26",x"51",x"10",x"51"),
   361 => (x"3f",x"20",x"27",x"4a"),
   362 => (x"27",x"49",x"00",x"00"),
   363 => (x"00",x"00",x"10",x"39"),
   364 => (x"20",x"1e",x"72",x"48"),
   365 => (x"20",x"41",x"20",x"41"),
   366 => (x"20",x"41",x"20",x"41"),
   367 => (x"20",x"41",x"20",x"41"),
   368 => (x"10",x"51",x"10",x"41"),
   369 => (x"26",x"51",x"10",x"51"),
   370 => (x"1d",x"f4",x"27",x"4a"),
   371 => (x"ca",x"49",x"00",x"00"),
   372 => (x"10",x"58",x"27",x"79"),
   373 => (x"27",x"1e",x"00",x"00"),
   374 => (x"00",x"00",x"01",x"51"),
   375 => (x"27",x"86",x"c4",x"0f"),
   376 => (x"00",x"00",x"10",x"5a"),
   377 => (x"01",x"51",x"27",x"1e"),
   378 => (x"c4",x"0f",x"00",x"00"),
   379 => (x"10",x"8a",x"27",x"86"),
   380 => (x"27",x"1e",x"00",x"00"),
   381 => (x"00",x"00",x"01",x"51"),
   382 => (x"27",x"86",x"c4",x"0f"),
   383 => (x"00",x"00",x"16",x"40"),
   384 => (x"df",x"c0",x"02",x"bf"),
   385 => (x"0e",x"a1",x"27",x"87"),
   386 => (x"27",x"1e",x"00",x"00"),
   387 => (x"00",x"00",x"01",x"51"),
   388 => (x"27",x"86",x"c4",x"0f"),
   389 => (x"00",x"00",x"0e",x"cd"),
   390 => (x"01",x"51",x"27",x"1e"),
   391 => (x"c4",x"0f",x"00",x"00"),
   392 => (x"87",x"dc",x"c0",x"86"),
   393 => (x"00",x"0e",x"cf",x"27"),
   394 => (x"51",x"27",x"1e",x"00"),
   395 => (x"0f",x"00",x"00",x"01"),
   396 => (x"fe",x"27",x"86",x"c4"),
   397 => (x"1e",x"00",x"00",x"0e"),
   398 => (x"00",x"01",x"51",x"27"),
   399 => (x"86",x"c4",x"0f",x"00"),
   400 => (x"00",x"16",x"44",x"27"),
   401 => (x"27",x"1e",x"bf",x"00"),
   402 => (x"00",x"00",x"10",x"8c"),
   403 => (x"01",x"51",x"27",x"1e"),
   404 => (x"c8",x"0f",x"00",x"00"),
   405 => (x"05",x"31",x"27",x"86"),
   406 => (x"27",x"0f",x"00",x"00"),
   407 => (x"00",x"00",x"3e",x"ac"),
   408 => (x"27",x"4d",x"c1",x"58"),
   409 => (x"00",x"00",x"16",x"44"),
   410 => (x"b7",x"c0",x"49",x"bf"),
   411 => (x"f9",x"c6",x"06",x"a9"),
   412 => (x"0e",x"7c",x"27",x"87"),
   413 => (x"27",x"0f",x"00",x"00"),
   414 => (x"00",x"00",x"0e",x"3b"),
   415 => (x"c2",x"49",x"76",x"0f"),
   416 => (x"27",x"4c",x"c3",x"79"),
   417 => (x"00",x"00",x"3f",x"40"),
   418 => (x"0f",x"1f",x"27",x"49"),
   419 => (x"72",x"48",x"00",x"00"),
   420 => (x"20",x"41",x"20",x"1e"),
   421 => (x"20",x"41",x"20",x"41"),
   422 => (x"20",x"41",x"20",x"41"),
   423 => (x"10",x"41",x"20",x"41"),
   424 => (x"10",x"51",x"10",x"51"),
   425 => (x"c8",x"4a",x"26",x"51"),
   426 => (x"79",x"c1",x"49",x"a6"),
   427 => (x"00",x"3f",x"40",x"27"),
   428 => (x"20",x"27",x"1e",x"00"),
   429 => (x"1e",x"00",x"00",x"3f"),
   430 => (x"00",x"03",x"fd",x"27"),
   431 => (x"86",x"c8",x"0f",x"00"),
   432 => (x"9a",x"72",x"4a",x"70"),
   433 => (x"87",x"c5",x"c0",x"05"),
   434 => (x"c2",x"c0",x"4a",x"c1"),
   435 => (x"27",x"4a",x"c0",x"87"),
   436 => (x"00",x"00",x"16",x"c4"),
   437 => (x"6e",x"79",x"72",x"49"),
   438 => (x"a9",x"b7",x"74",x"49"),
   439 => (x"87",x"ed",x"c0",x"03"),
   440 => (x"92",x"c5",x"4a",x"6e"),
   441 => (x"88",x"74",x"48",x"72"),
   442 => (x"cc",x"58",x"a6",x"d0"),
   443 => (x"1e",x"72",x"4a",x"a6"),
   444 => (x"66",x"c8",x"1e",x"74"),
   445 => (x"03",x"16",x"27",x"1e"),
   446 => (x"cc",x"0f",x"00",x"00"),
   447 => (x"c1",x"48",x"6e",x"86"),
   448 => (x"58",x"a6",x"c4",x"80"),
   449 => (x"b7",x"74",x"49",x"6e"),
   450 => (x"d3",x"ff",x"04",x"a9"),
   451 => (x"1e",x"66",x"cc",x"87"),
   452 => (x"27",x"1e",x"66",x"c4"),
   453 => (x"00",x"00",x"17",x"98"),
   454 => (x"16",x"d0",x"27",x"1e"),
   455 => (x"27",x"1e",x"00",x"00"),
   456 => (x"00",x"00",x"03",x"2c"),
   457 => (x"27",x"86",x"d0",x"0f"),
   458 => (x"00",x"00",x"16",x"b8"),
   459 => (x"1c",x"27",x"1e",x"bf"),
   460 => (x"0f",x"00",x"00",x"0d"),
   461 => (x"a6",x"c4",x"86",x"c4"),
   462 => (x"51",x"c1",x"c1",x"49"),
   463 => (x"00",x"16",x"c9",x"27"),
   464 => (x"4a",x"bf",x"97",x"00"),
   465 => (x"c0",x"c0",x"c0",x"c1"),
   466 => (x"c0",x"c4",x"92",x"c0"),
   467 => (x"c1",x"4a",x"92",x"b7"),
   468 => (x"04",x"aa",x"b7",x"c1"),
   469 => (x"c1",x"87",x"d8",x"c2"),
   470 => (x"c8",x"97",x"1e",x"c3"),
   471 => (x"c0",x"c1",x"4a",x"66"),
   472 => (x"92",x"c0",x"c0",x"c0"),
   473 => (x"92",x"b7",x"c0",x"c4"),
   474 => (x"27",x"1e",x"72",x"4a"),
   475 => (x"00",x"00",x"03",x"b9"),
   476 => (x"70",x"86",x"c8",x"0f"),
   477 => (x"49",x"66",x"c8",x"4a"),
   478 => (x"05",x"a9",x"b7",x"72"),
   479 => (x"c8",x"87",x"fd",x"c0"),
   480 => (x"1e",x"72",x"4a",x"a6"),
   481 => (x"9f",x"27",x"1e",x"c0"),
   482 => (x"0f",x"00",x"00",x"02"),
   483 => (x"40",x"27",x"86",x"c8"),
   484 => (x"49",x"00",x"00",x"3f"),
   485 => (x"00",x"0f",x"00",x"27"),
   486 => (x"1e",x"72",x"48",x"00"),
   487 => (x"41",x"20",x"41",x"20"),
   488 => (x"41",x"20",x"41",x"20"),
   489 => (x"41",x"20",x"41",x"20"),
   490 => (x"51",x"10",x"41",x"20"),
   491 => (x"51",x"10",x"51",x"10"),
   492 => (x"4c",x"75",x"4a",x"26"),
   493 => (x"00",x"16",x"c0",x"27"),
   494 => (x"79",x"75",x"49",x"00"),
   495 => (x"48",x"66",x"c4",x"97"),
   496 => (x"a6",x"c4",x"80",x"c1"),
   497 => (x"c4",x"97",x"50",x"08"),
   498 => (x"c0",x"c1",x"4b",x"66"),
   499 => (x"93",x"c0",x"c0",x"c0"),
   500 => (x"93",x"b7",x"c0",x"c4"),
   501 => (x"16",x"c9",x"27",x"4b"),
   502 => (x"bf",x"97",x"00",x"00"),
   503 => (x"c0",x"c0",x"c1",x"4a"),
   504 => (x"c4",x"92",x"c0",x"c0"),
   505 => (x"4a",x"92",x"b7",x"c0"),
   506 => (x"06",x"ab",x"b7",x"72"),
   507 => (x"6e",x"87",x"e8",x"fd"),
   508 => (x"72",x"49",x"74",x"94"),
   509 => (x"4a",x"66",x"d0",x"1e"),
   510 => (x"00",x"04",x"da",x"27"),
   511 => (x"4a",x"26",x"0f",x"00"),
   512 => (x"a6",x"c4",x"48",x"70"),
   513 => (x"cc",x"4a",x"74",x"58"),
   514 => (x"92",x"c7",x"8a",x"66"),
   515 => (x"8c",x"6e",x"4c",x"72"),
   516 => (x"1e",x"72",x"4a",x"76"),
   517 => (x"00",x"0d",x"b7",x"27"),
   518 => (x"86",x"c4",x"0f",x"00"),
   519 => (x"44",x"27",x"85",x"c1"),
   520 => (x"bf",x"00",x"00",x"16"),
   521 => (x"f9",x"06",x"ad",x"b7"),
   522 => (x"31",x"27",x"87",x"c7"),
   523 => (x"0f",x"00",x"00",x"05"),
   524 => (x"00",x"3e",x"b0",x"27"),
   525 => (x"b9",x"27",x"58",x"00"),
   526 => (x"1e",x"00",x"00",x"10"),
   527 => (x"00",x"01",x"51",x"27"),
   528 => (x"86",x"c4",x"0f",x"00"),
   529 => (x"00",x"10",x"c9",x"27"),
   530 => (x"51",x"27",x"1e",x"00"),
   531 => (x"0f",x"00",x"00",x"01"),
   532 => (x"cb",x"27",x"86",x"c4"),
   533 => (x"1e",x"00",x"00",x"10"),
   534 => (x"00",x"01",x"51",x"27"),
   535 => (x"86",x"c4",x"0f",x"00"),
   536 => (x"00",x"11",x"01",x"27"),
   537 => (x"51",x"27",x"1e",x"00"),
   538 => (x"0f",x"00",x"00",x"01"),
   539 => (x"c0",x"27",x"86",x"c4"),
   540 => (x"bf",x"00",x"00",x"16"),
   541 => (x"11",x"03",x"27",x"1e"),
   542 => (x"27",x"1e",x"00",x"00"),
   543 => (x"00",x"00",x"01",x"51"),
   544 => (x"c5",x"86",x"c8",x"0f"),
   545 => (x"11",x"1c",x"27",x"1e"),
   546 => (x"27",x"1e",x"00",x"00"),
   547 => (x"00",x"00",x"01",x"51"),
   548 => (x"27",x"86",x"c8",x"0f"),
   549 => (x"00",x"00",x"16",x"c4"),
   550 => (x"35",x"27",x"1e",x"bf"),
   551 => (x"1e",x"00",x"00",x"11"),
   552 => (x"00",x"01",x"51",x"27"),
   553 => (x"86",x"c8",x"0f",x"00"),
   554 => (x"4e",x"27",x"1e",x"c1"),
   555 => (x"1e",x"00",x"00",x"11"),
   556 => (x"00",x"01",x"51",x"27"),
   557 => (x"86",x"c8",x"0f",x"00"),
   558 => (x"00",x"16",x"c8",x"27"),
   559 => (x"4a",x"bf",x"97",x"00"),
   560 => (x"c0",x"c0",x"c0",x"c1"),
   561 => (x"c0",x"c4",x"92",x"c0"),
   562 => (x"72",x"4a",x"92",x"b7"),
   563 => (x"11",x"67",x"27",x"1e"),
   564 => (x"27",x"1e",x"00",x"00"),
   565 => (x"00",x"00",x"01",x"51"),
   566 => (x"c1",x"86",x"c8",x"0f"),
   567 => (x"80",x"27",x"1e",x"c1"),
   568 => (x"1e",x"00",x"00",x"11"),
   569 => (x"00",x"01",x"51",x"27"),
   570 => (x"86",x"c8",x"0f",x"00"),
   571 => (x"00",x"16",x"c9",x"27"),
   572 => (x"4a",x"bf",x"97",x"00"),
   573 => (x"c0",x"c0",x"c0",x"c1"),
   574 => (x"c0",x"c4",x"92",x"c0"),
   575 => (x"72",x"4a",x"92",x"b7"),
   576 => (x"11",x"99",x"27",x"1e"),
   577 => (x"27",x"1e",x"00",x"00"),
   578 => (x"00",x"00",x"01",x"51"),
   579 => (x"c1",x"86",x"c8",x"0f"),
   580 => (x"b2",x"27",x"1e",x"c2"),
   581 => (x"1e",x"00",x"00",x"11"),
   582 => (x"00",x"01",x"51",x"27"),
   583 => (x"86",x"c8",x"0f",x"00"),
   584 => (x"00",x"16",x"f0",x"27"),
   585 => (x"27",x"1e",x"bf",x"00"),
   586 => (x"00",x"00",x"11",x"cb"),
   587 => (x"01",x"51",x"27",x"1e"),
   588 => (x"c8",x"0f",x"00",x"00"),
   589 => (x"27",x"1e",x"c7",x"86"),
   590 => (x"00",x"00",x"11",x"e4"),
   591 => (x"01",x"51",x"27",x"1e"),
   592 => (x"c8",x"0f",x"00",x"00"),
   593 => (x"1d",x"f4",x"27",x"86"),
   594 => (x"1e",x"bf",x"00",x"00"),
   595 => (x"00",x"11",x"fd",x"27"),
   596 => (x"51",x"27",x"1e",x"00"),
   597 => (x"0f",x"00",x"00",x"01"),
   598 => (x"16",x"27",x"86",x"c8"),
   599 => (x"1e",x"00",x"00",x"12"),
   600 => (x"00",x"01",x"51",x"27"),
   601 => (x"86",x"c4",x"0f",x"00"),
   602 => (x"00",x"12",x"40",x"27"),
   603 => (x"51",x"27",x"1e",x"00"),
   604 => (x"0f",x"00",x"00",x"01"),
   605 => (x"b8",x"27",x"86",x"c4"),
   606 => (x"bf",x"00",x"00",x"16"),
   607 => (x"4c",x"27",x"1e",x"bf"),
   608 => (x"1e",x"00",x"00",x"12"),
   609 => (x"00",x"01",x"51",x"27"),
   610 => (x"86",x"c8",x"0f",x"00"),
   611 => (x"00",x"12",x"65",x"27"),
   612 => (x"51",x"27",x"1e",x"00"),
   613 => (x"0f",x"00",x"00",x"01"),
   614 => (x"b8",x"27",x"86",x"c4"),
   615 => (x"bf",x"00",x"00",x"16"),
   616 => (x"6a",x"82",x"c4",x"4a"),
   617 => (x"12",x"96",x"27",x"1e"),
   618 => (x"27",x"1e",x"00",x"00"),
   619 => (x"00",x"00",x"01",x"51"),
   620 => (x"c0",x"86",x"c8",x"0f"),
   621 => (x"12",x"af",x"27",x"1e"),
   622 => (x"27",x"1e",x"00",x"00"),
   623 => (x"00",x"00",x"01",x"51"),
   624 => (x"27",x"86",x"c8",x"0f"),
   625 => (x"00",x"00",x"16",x"b8"),
   626 => (x"82",x"c8",x"4a",x"bf"),
   627 => (x"c8",x"27",x"1e",x"6a"),
   628 => (x"1e",x"00",x"00",x"12"),
   629 => (x"00",x"01",x"51",x"27"),
   630 => (x"86",x"c8",x"0f",x"00"),
   631 => (x"e1",x"27",x"1e",x"c2"),
   632 => (x"1e",x"00",x"00",x"12"),
   633 => (x"00",x"01",x"51",x"27"),
   634 => (x"86",x"c8",x"0f",x"00"),
   635 => (x"00",x"16",x"b8",x"27"),
   636 => (x"cc",x"4a",x"bf",x"00"),
   637 => (x"27",x"1e",x"6a",x"82"),
   638 => (x"00",x"00",x"12",x"fa"),
   639 => (x"01",x"51",x"27",x"1e"),
   640 => (x"c8",x"0f",x"00",x"00"),
   641 => (x"27",x"1e",x"d1",x"86"),
   642 => (x"00",x"00",x"13",x"13"),
   643 => (x"01",x"51",x"27",x"1e"),
   644 => (x"c8",x"0f",x"00",x"00"),
   645 => (x"16",x"b8",x"27",x"86"),
   646 => (x"4a",x"bf",x"00",x"00"),
   647 => (x"1e",x"72",x"82",x"d0"),
   648 => (x"00",x"13",x"2c",x"27"),
   649 => (x"51",x"27",x"1e",x"00"),
   650 => (x"0f",x"00",x"00",x"01"),
   651 => (x"45",x"27",x"86",x"c8"),
   652 => (x"1e",x"00",x"00",x"13"),
   653 => (x"00",x"01",x"51",x"27"),
   654 => (x"86",x"c4",x"0f",x"00"),
   655 => (x"00",x"13",x"7a",x"27"),
   656 => (x"51",x"27",x"1e",x"00"),
   657 => (x"0f",x"00",x"00",x"01"),
   658 => (x"bc",x"27",x"86",x"c4"),
   659 => (x"bf",x"00",x"00",x"16"),
   660 => (x"8b",x"27",x"1e",x"bf"),
   661 => (x"1e",x"00",x"00",x"13"),
   662 => (x"00",x"01",x"51",x"27"),
   663 => (x"86",x"c8",x"0f",x"00"),
   664 => (x"00",x"13",x"a4",x"27"),
   665 => (x"51",x"27",x"1e",x"00"),
   666 => (x"0f",x"00",x"00",x"01"),
   667 => (x"bc",x"27",x"86",x"c4"),
   668 => (x"bf",x"00",x"00",x"16"),
   669 => (x"6a",x"82",x"c4",x"4a"),
   670 => (x"13",x"e4",x"27",x"1e"),
   671 => (x"27",x"1e",x"00",x"00"),
   672 => (x"00",x"00",x"01",x"51"),
   673 => (x"c0",x"86",x"c8",x"0f"),
   674 => (x"13",x"fd",x"27",x"1e"),
   675 => (x"27",x"1e",x"00",x"00"),
   676 => (x"00",x"00",x"01",x"51"),
   677 => (x"27",x"86",x"c8",x"0f"),
   678 => (x"00",x"00",x"16",x"bc"),
   679 => (x"82",x"c8",x"4a",x"bf"),
   680 => (x"16",x"27",x"1e",x"6a"),
   681 => (x"1e",x"00",x"00",x"14"),
   682 => (x"00",x"01",x"51",x"27"),
   683 => (x"86",x"c8",x"0f",x"00"),
   684 => (x"2f",x"27",x"1e",x"c1"),
   685 => (x"1e",x"00",x"00",x"14"),
   686 => (x"00",x"01",x"51",x"27"),
   687 => (x"86",x"c8",x"0f",x"00"),
   688 => (x"00",x"16",x"bc",x"27"),
   689 => (x"cc",x"4a",x"bf",x"00"),
   690 => (x"27",x"1e",x"6a",x"82"),
   691 => (x"00",x"00",x"14",x"48"),
   692 => (x"01",x"51",x"27",x"1e"),
   693 => (x"c8",x"0f",x"00",x"00"),
   694 => (x"27",x"1e",x"d2",x"86"),
   695 => (x"00",x"00",x"14",x"61"),
   696 => (x"01",x"51",x"27",x"1e"),
   697 => (x"c8",x"0f",x"00",x"00"),
   698 => (x"16",x"bc",x"27",x"86"),
   699 => (x"4a",x"bf",x"00",x"00"),
   700 => (x"1e",x"72",x"82",x"d0"),
   701 => (x"00",x"14",x"7a",x"27"),
   702 => (x"51",x"27",x"1e",x"00"),
   703 => (x"0f",x"00",x"00",x"01"),
   704 => (x"93",x"27",x"86",x"c8"),
   705 => (x"1e",x"00",x"00",x"14"),
   706 => (x"00",x"01",x"51",x"27"),
   707 => (x"86",x"c4",x"0f",x"00"),
   708 => (x"c8",x"27",x"1e",x"6e"),
   709 => (x"1e",x"00",x"00",x"14"),
   710 => (x"00",x"01",x"51",x"27"),
   711 => (x"86",x"c8",x"0f",x"00"),
   712 => (x"e1",x"27",x"1e",x"c5"),
   713 => (x"1e",x"00",x"00",x"14"),
   714 => (x"00",x"01",x"51",x"27"),
   715 => (x"86",x"c8",x"0f",x"00"),
   716 => (x"fa",x"27",x"1e",x"74"),
   717 => (x"1e",x"00",x"00",x"14"),
   718 => (x"00",x"01",x"51",x"27"),
   719 => (x"86",x"c8",x"0f",x"00"),
   720 => (x"13",x"27",x"1e",x"cd"),
   721 => (x"1e",x"00",x"00",x"15"),
   722 => (x"00",x"01",x"51",x"27"),
   723 => (x"86",x"c8",x"0f",x"00"),
   724 => (x"27",x"1e",x"66",x"cc"),
   725 => (x"00",x"00",x"15",x"2c"),
   726 => (x"01",x"51",x"27",x"1e"),
   727 => (x"c8",x"0f",x"00",x"00"),
   728 => (x"27",x"1e",x"c7",x"86"),
   729 => (x"00",x"00",x"15",x"45"),
   730 => (x"01",x"51",x"27",x"1e"),
   731 => (x"c8",x"0f",x"00",x"00"),
   732 => (x"1e",x"66",x"c8",x"86"),
   733 => (x"00",x"15",x"5e",x"27"),
   734 => (x"51",x"27",x"1e",x"00"),
   735 => (x"0f",x"00",x"00",x"01"),
   736 => (x"1e",x"c1",x"86",x"c8"),
   737 => (x"00",x"15",x"77",x"27"),
   738 => (x"51",x"27",x"1e",x"00"),
   739 => (x"0f",x"00",x"00",x"01"),
   740 => (x"20",x"27",x"86",x"c8"),
   741 => (x"1e",x"00",x"00",x"3f"),
   742 => (x"00",x"15",x"90",x"27"),
   743 => (x"51",x"27",x"1e",x"00"),
   744 => (x"0f",x"00",x"00",x"01"),
   745 => (x"a9",x"27",x"86",x"c8"),
   746 => (x"1e",x"00",x"00",x"15"),
   747 => (x"00",x"01",x"51",x"27"),
   748 => (x"86",x"c4",x"0f",x"00"),
   749 => (x"00",x"3f",x"40",x"27"),
   750 => (x"de",x"27",x"1e",x"00"),
   751 => (x"1e",x"00",x"00",x"15"),
   752 => (x"00",x"01",x"51",x"27"),
   753 => (x"86",x"c8",x"0f",x"00"),
   754 => (x"00",x"15",x"f7",x"27"),
   755 => (x"51",x"27",x"1e",x"00"),
   756 => (x"0f",x"00",x"00",x"01"),
   757 => (x"2c",x"27",x"86",x"c4"),
   758 => (x"1e",x"00",x"00",x"16"),
   759 => (x"00",x"01",x"51",x"27"),
   760 => (x"86",x"c4",x"0f",x"00"),
   761 => (x"00",x"3e",x"ac",x"27"),
   762 => (x"27",x"4a",x"bf",x"00"),
   763 => (x"00",x"00",x"3e",x"a8"),
   764 => (x"b0",x"27",x"8a",x"bf"),
   765 => (x"49",x"00",x"00",x"3e"),
   766 => (x"1e",x"72",x"79",x"72"),
   767 => (x"00",x"16",x"2e",x"27"),
   768 => (x"51",x"27",x"1e",x"00"),
   769 => (x"0f",x"00",x"00",x"01"),
   770 => (x"b0",x"27",x"86",x"c8"),
   771 => (x"bf",x"00",x"00",x"3e"),
   772 => (x"b7",x"f8",x"c1",x"49"),
   773 => (x"ea",x"c0",x"03",x"a9"),
   774 => (x"0f",x"3e",x"27",x"87"),
   775 => (x"27",x"1e",x"00",x"00"),
   776 => (x"00",x"00",x"01",x"51"),
   777 => (x"27",x"86",x"c4",x"0f"),
   778 => (x"00",x"00",x"0f",x"74"),
   779 => (x"01",x"51",x"27",x"1e"),
   780 => (x"c4",x"0f",x"00",x"00"),
   781 => (x"0f",x"94",x"27",x"86"),
   782 => (x"27",x"1e",x"00",x"00"),
   783 => (x"00",x"00",x"01",x"51"),
   784 => (x"27",x"86",x"c4",x"0f"),
   785 => (x"00",x"00",x"3e",x"b0"),
   786 => (x"4b",x"72",x"4a",x"bf"),
   787 => (x"73",x"93",x"e8",x"cf"),
   788 => (x"27",x"1e",x"72",x"49"),
   789 => (x"00",x"00",x"16",x"44"),
   790 => (x"da",x"27",x"4a",x"bf"),
   791 => (x"0f",x"00",x"00",x"04"),
   792 => (x"48",x"70",x"4a",x"26"),
   793 => (x"00",x"3e",x"b8",x"27"),
   794 => (x"44",x"27",x"58",x"00"),
   795 => (x"bf",x"00",x"00",x"16"),
   796 => (x"cf",x"4c",x"73",x"4b"),
   797 => (x"49",x"74",x"94",x"e8"),
   798 => (x"4a",x"72",x"1e",x"72"),
   799 => (x"00",x"04",x"da",x"27"),
   800 => (x"4a",x"26",x"0f",x"00"),
   801 => (x"bc",x"27",x"48",x"70"),
   802 => (x"58",x"00",x"00",x"3e"),
   803 => (x"73",x"93",x"f9",x"c8"),
   804 => (x"72",x"1e",x"72",x"49"),
   805 => (x"04",x"da",x"27",x"4a"),
   806 => (x"26",x"0f",x"00",x"00"),
   807 => (x"27",x"48",x"70",x"4a"),
   808 => (x"00",x"00",x"3e",x"c0"),
   809 => (x"0f",x"96",x"27",x"58"),
   810 => (x"27",x"1e",x"00",x"00"),
   811 => (x"00",x"00",x"01",x"51"),
   812 => (x"27",x"86",x"c4",x"0f"),
   813 => (x"00",x"00",x"3e",x"b4"),
   814 => (x"c3",x"27",x"1e",x"bf"),
   815 => (x"1e",x"00",x"00",x"0f"),
   816 => (x"00",x"01",x"51",x"27"),
   817 => (x"86",x"c8",x"0f",x"00"),
   818 => (x"00",x"0f",x"c8",x"27"),
   819 => (x"51",x"27",x"1e",x"00"),
   820 => (x"0f",x"00",x"00",x"01"),
   821 => (x"b8",x"27",x"86",x"c4"),
   822 => (x"bf",x"00",x"00",x"3e"),
   823 => (x"0f",x"f5",x"27",x"1e"),
   824 => (x"27",x"1e",x"00",x"00"),
   825 => (x"00",x"00",x"01",x"51"),
   826 => (x"27",x"86",x"c8",x"0f"),
   827 => (x"00",x"00",x"3e",x"bc"),
   828 => (x"fa",x"27",x"1e",x"bf"),
   829 => (x"1e",x"00",x"00",x"0f"),
   830 => (x"00",x"01",x"51",x"27"),
   831 => (x"86",x"c8",x"0f",x"00"),
   832 => (x"00",x"10",x"18",x"27"),
   833 => (x"51",x"27",x"1e",x"00"),
   834 => (x"0f",x"00",x"00",x"01"),
   835 => (x"48",x"c0",x"86",x"c4"),
   836 => (x"4d",x"26",x"86",x"d0"),
   837 => (x"4b",x"26",x"4c",x"26"),
   838 => (x"4f",x"26",x"4a",x"26"),
   839 => (x"5b",x"5a",x"5e",x"0e"),
   840 => (x"d4",x"0e",x"5d",x"5c"),
   841 => (x"72",x"4a",x"bf",x"66"),
   842 => (x"16",x"b8",x"27",x"4d"),
   843 => (x"48",x"bf",x"00",x"00"),
   844 => (x"f0",x"c0",x"1e",x"72"),
   845 => (x"42",x"20",x"49",x"a2"),
   846 => (x"f9",x"05",x"a9",x"72"),
   847 => (x"d4",x"4a",x"26",x"87"),
   848 => (x"84",x"cc",x"4c",x"66"),
   849 => (x"4b",x"72",x"7c",x"c5"),
   850 => (x"7b",x"6c",x"83",x"cc"),
   851 => (x"7a",x"bf",x"66",x"d4"),
   852 => (x"03",x"27",x"1e",x"72"),
   853 => (x"0f",x"00",x"00",x"0e"),
   854 => (x"82",x"c4",x"86",x"c4"),
   855 => (x"c0",x"05",x"9a",x"6a"),
   856 => (x"4b",x"75",x"87",x"f4"),
   857 => (x"4a",x"75",x"83",x"c8"),
   858 => (x"7a",x"c6",x"82",x"cc"),
   859 => (x"66",x"d8",x"1e",x"73"),
   860 => (x"6b",x"83",x"c8",x"4b"),
   861 => (x"02",x"9f",x"27",x"1e"),
   862 => (x"c8",x"0f",x"00",x"00"),
   863 => (x"16",x"b8",x"27",x"86"),
   864 => (x"bf",x"bf",x"00",x"00"),
   865 => (x"ca",x"1e",x"72",x"7d"),
   866 => (x"27",x"1e",x"6a",x"1e"),
   867 => (x"00",x"00",x"03",x"16"),
   868 => (x"c0",x"86",x"cc",x"0f"),
   869 => (x"66",x"d4",x"87",x"d7"),
   870 => (x"66",x"d4",x"4a",x"bf"),
   871 => (x"1e",x"72",x"48",x"49"),
   872 => (x"4a",x"a1",x"f0",x"c0"),
   873 => (x"aa",x"71",x"41",x"20"),
   874 => (x"26",x"87",x"f9",x"05"),
   875 => (x"26",x"4d",x"26",x"4a"),
   876 => (x"26",x"4b",x"26",x"4c"),
   877 => (x"0e",x"4f",x"26",x"4a"),
   878 => (x"5c",x"5b",x"5a",x"5e"),
   879 => (x"6e",x"1e",x"0e",x"5d"),
   880 => (x"4c",x"66",x"d8",x"4d"),
   881 => (x"83",x"ca",x"4b",x"6c"),
   882 => (x"00",x"16",x"c8",x"27"),
   883 => (x"4a",x"bf",x"97",x"00"),
   884 => (x"c0",x"c0",x"c0",x"c1"),
   885 => (x"c0",x"c4",x"92",x"c0"),
   886 => (x"c1",x"4a",x"92",x"b7"),
   887 => (x"05",x"aa",x"b7",x"c1"),
   888 => (x"c1",x"87",x"cf",x"c0"),
   889 => (x"27",x"48",x"73",x"8b"),
   890 => (x"00",x"00",x"16",x"c0"),
   891 => (x"7c",x"70",x"88",x"bf"),
   892 => (x"9d",x"75",x"4d",x"c0"),
   893 => (x"87",x"d0",x"ff",x"05"),
   894 => (x"26",x"4d",x"26",x"26"),
   895 => (x"26",x"4b",x"26",x"4c"),
   896 => (x"1e",x"4f",x"26",x"4a"),
   897 => (x"b8",x"27",x"1e",x"72"),
   898 => (x"bf",x"00",x"00",x"16"),
   899 => (x"87",x"cb",x"c0",x"02"),
   900 => (x"27",x"49",x"66",x"c8"),
   901 => (x"00",x"00",x"16",x"b8"),
   902 => (x"27",x"79",x"bf",x"bf"),
   903 => (x"00",x"00",x"16",x"b8"),
   904 => (x"82",x"cc",x"4a",x"bf"),
   905 => (x"c0",x"27",x"1e",x"72"),
   906 => (x"bf",x"00",x"00",x"16"),
   907 => (x"27",x"1e",x"ca",x"1e"),
   908 => (x"00",x"00",x"03",x"16"),
   909 => (x"26",x"86",x"cc",x"0f"),
   910 => (x"1e",x"4f",x"26",x"4a"),
   911 => (x"c8",x"27",x"1e",x"72"),
   912 => (x"97",x"00",x"00",x"16"),
   913 => (x"c0",x"c1",x"4a",x"bf"),
   914 => (x"92",x"c0",x"c0",x"c0"),
   915 => (x"92",x"b7",x"c0",x"c4"),
   916 => (x"b7",x"c1",x"c1",x"4a"),
   917 => (x"c5",x"c0",x"02",x"aa"),
   918 => (x"c0",x"4a",x"c0",x"87"),
   919 => (x"4a",x"c1",x"87",x"c2"),
   920 => (x"00",x"16",x"c4",x"27"),
   921 => (x"72",x"48",x"bf",x"00"),
   922 => (x"16",x"c8",x"27",x"b0"),
   923 => (x"27",x"58",x"00",x"00"),
   924 => (x"00",x"00",x"16",x"c9"),
   925 => (x"51",x"c2",x"c1",x"49"),
   926 => (x"4f",x"26",x"4a",x"26"),
   927 => (x"16",x"c8",x"27",x"1e"),
   928 => (x"c1",x"49",x"00",x"00"),
   929 => (x"c4",x"27",x"51",x"c1"),
   930 => (x"49",x"00",x"00",x"16"),
   931 => (x"4f",x"26",x"79",x"c0"),
   932 => (x"33",x"32",x"31",x"30"),
   933 => (x"37",x"36",x"35",x"34"),
   934 => (x"42",x"41",x"39",x"38"),
   935 => (x"46",x"45",x"44",x"43"),
   936 => (x"6f",x"72",x"50",x"00"),
   937 => (x"6d",x"61",x"72",x"67"),
   938 => (x"6d",x"6f",x"63",x"20"),
   939 => (x"65",x"6c",x"69",x"70"),
   940 => (x"69",x"77",x"20",x"64"),
   941 => (x"27",x"20",x"68",x"74"),
   942 => (x"69",x"67",x"65",x"72"),
   943 => (x"72",x"65",x"74",x"73"),
   944 => (x"74",x"61",x"20",x"27"),
   945 => (x"62",x"69",x"72",x"74"),
   946 => (x"0a",x"65",x"74",x"75"),
   947 => (x"50",x"00",x"0a",x"00"),
   948 => (x"72",x"67",x"6f",x"72"),
   949 => (x"63",x"20",x"6d",x"61"),
   950 => (x"69",x"70",x"6d",x"6f"),
   951 => (x"20",x"64",x"65",x"6c"),
   952 => (x"68",x"74",x"69",x"77"),
   953 => (x"20",x"74",x"75",x"6f"),
   954 => (x"67",x"65",x"72",x"27"),
   955 => (x"65",x"74",x"73",x"69"),
   956 => (x"61",x"20",x"27",x"72"),
   957 => (x"69",x"72",x"74",x"74"),
   958 => (x"65",x"74",x"75",x"62"),
   959 => (x"00",x"0a",x"00",x"0a"),
   960 => (x"59",x"52",x"48",x"44"),
   961 => (x"4e",x"4f",x"54",x"53"),
   962 => (x"52",x"50",x"20",x"45"),
   963 => (x"41",x"52",x"47",x"4f"),
   964 => (x"33",x"20",x"2c",x"4d"),
   965 => (x"20",x"44",x"52",x"27"),
   966 => (x"49",x"52",x"54",x"53"),
   967 => (x"44",x"00",x"47",x"4e"),
   968 => (x"53",x"59",x"52",x"48"),
   969 => (x"45",x"4e",x"4f",x"54"),
   970 => (x"4f",x"52",x"50",x"20"),
   971 => (x"4d",x"41",x"52",x"47"),
   972 => (x"27",x"32",x"20",x"2c"),
   973 => (x"53",x"20",x"44",x"4e"),
   974 => (x"4e",x"49",x"52",x"54"),
   975 => (x"65",x"4d",x"00",x"47"),
   976 => (x"72",x"75",x"73",x"61"),
   977 => (x"74",x"20",x"64",x"65"),
   978 => (x"20",x"65",x"6d",x"69"),
   979 => (x"20",x"6f",x"6f",x"74"),
   980 => (x"6c",x"61",x"6d",x"73"),
   981 => (x"6f",x"74",x"20",x"6c"),
   982 => (x"74",x"62",x"6f",x"20"),
   983 => (x"20",x"6e",x"69",x"61"),
   984 => (x"6e",x"61",x"65",x"6d"),
   985 => (x"66",x"67",x"6e",x"69"),
   986 => (x"72",x"20",x"6c",x"75"),
   987 => (x"6c",x"75",x"73",x"65"),
   988 => (x"00",x"0a",x"73",x"74"),
   989 => (x"61",x"65",x"6c",x"50"),
   990 => (x"69",x"20",x"65",x"73"),
   991 => (x"65",x"72",x"63",x"6e"),
   992 => (x"20",x"65",x"73",x"61"),
   993 => (x"62",x"6d",x"75",x"6e"),
   994 => (x"6f",x"20",x"72",x"65"),
   995 => (x"75",x"72",x"20",x"66"),
   996 => (x"00",x"0a",x"73",x"6e"),
   997 => (x"69",x"4d",x"00",x"0a"),
   998 => (x"73",x"6f",x"72",x"63"),
   999 => (x"6e",x"6f",x"63",x"65"),
  1000 => (x"66",x"20",x"73",x"64"),
  1001 => (x"6f",x"20",x"72",x"6f"),
  1002 => (x"72",x"20",x"65",x"6e"),
  1003 => (x"74",x"20",x"6e",x"75"),
  1004 => (x"75",x"6f",x"72",x"68"),
  1005 => (x"44",x"20",x"68",x"67"),
  1006 => (x"73",x"79",x"72",x"68"),
  1007 => (x"65",x"6e",x"6f",x"74"),
  1008 => (x"25",x"00",x"20",x"3a"),
  1009 => (x"00",x"0a",x"20",x"64"),
  1010 => (x"79",x"72",x"68",x"44"),
  1011 => (x"6e",x"6f",x"74",x"73"),
  1012 => (x"70",x"20",x"73",x"65"),
  1013 => (x"53",x"20",x"72",x"65"),
  1014 => (x"6e",x"6f",x"63",x"65"),
  1015 => (x"20",x"20",x"3a",x"64"),
  1016 => (x"20",x"20",x"20",x"20"),
  1017 => (x"20",x"20",x"20",x"20"),
  1018 => (x"20",x"20",x"20",x"20"),
  1019 => (x"20",x"20",x"20",x"20"),
  1020 => (x"20",x"20",x"20",x"20"),
  1021 => (x"20",x"64",x"25",x"00"),
  1022 => (x"41",x"56",x"00",x"0a"),
  1023 => (x"49",x"4d",x"20",x"58"),
  1024 => (x"72",x"20",x"53",x"50"),
  1025 => (x"6e",x"69",x"74",x"61"),
  1026 => (x"20",x"2a",x"20",x"67"),
  1027 => (x"30",x"30",x"30",x"31"),
  1028 => (x"25",x"20",x"3d",x"20"),
  1029 => (x"00",x"0a",x"20",x"64"),
  1030 => (x"48",x"44",x"00",x"0a"),
  1031 => (x"54",x"53",x"59",x"52"),
  1032 => (x"20",x"45",x"4e",x"4f"),
  1033 => (x"47",x"4f",x"52",x"50"),
  1034 => (x"2c",x"4d",x"41",x"52"),
  1035 => (x"4d",x"4f",x"53",x"20"),
  1036 => (x"54",x"53",x"20",x"45"),
  1037 => (x"47",x"4e",x"49",x"52"),
  1038 => (x"52",x"48",x"44",x"00"),
  1039 => (x"4f",x"54",x"53",x"59"),
  1040 => (x"50",x"20",x"45",x"4e"),
  1041 => (x"52",x"47",x"4f",x"52"),
  1042 => (x"20",x"2c",x"4d",x"41"),
  1043 => (x"54",x"53",x"27",x"31"),
  1044 => (x"52",x"54",x"53",x"20"),
  1045 => (x"00",x"47",x"4e",x"49"),
  1046 => (x"68",x"44",x"00",x"0a"),
  1047 => (x"74",x"73",x"79",x"72"),
  1048 => (x"20",x"65",x"6e",x"6f"),
  1049 => (x"63",x"6e",x"65",x"42"),
  1050 => (x"72",x"61",x"6d",x"68"),
  1051 => (x"56",x"20",x"2c",x"6b"),
  1052 => (x"69",x"73",x"72",x"65"),
  1053 => (x"32",x"20",x"6e",x"6f"),
  1054 => (x"28",x"20",x"31",x"2e"),
  1055 => (x"67",x"6e",x"61",x"4c"),
  1056 => (x"65",x"67",x"61",x"75"),
  1057 => (x"29",x"43",x"20",x"3a"),
  1058 => (x"00",x"0a",x"00",x"0a"),
  1059 => (x"63",x"65",x"78",x"45"),
  1060 => (x"6f",x"69",x"74",x"75"),
  1061 => (x"74",x"73",x"20",x"6e"),
  1062 => (x"73",x"74",x"72",x"61"),
  1063 => (x"64",x"25",x"20",x"2c"),
  1064 => (x"6e",x"75",x"72",x"20"),
  1065 => (x"68",x"74",x"20",x"73"),
  1066 => (x"67",x"75",x"6f",x"72"),
  1067 => (x"68",x"44",x"20",x"68"),
  1068 => (x"74",x"73",x"79",x"72"),
  1069 => (x"0a",x"65",x"6e",x"6f"),
  1070 => (x"65",x"78",x"45",x"00"),
  1071 => (x"69",x"74",x"75",x"63"),
  1072 => (x"65",x"20",x"6e",x"6f"),
  1073 => (x"0a",x"73",x"64",x"6e"),
  1074 => (x"46",x"00",x"0a",x"00"),
  1075 => (x"6c",x"61",x"6e",x"69"),
  1076 => (x"6c",x"61",x"76",x"20"),
  1077 => (x"20",x"73",x"65",x"75"),
  1078 => (x"74",x"20",x"66",x"6f"),
  1079 => (x"76",x"20",x"65",x"68"),
  1080 => (x"61",x"69",x"72",x"61"),
  1081 => (x"73",x"65",x"6c",x"62"),
  1082 => (x"65",x"73",x"75",x"20"),
  1083 => (x"6e",x"69",x"20",x"64"),
  1084 => (x"65",x"68",x"74",x"20"),
  1085 => (x"6e",x"65",x"62",x"20"),
  1086 => (x"61",x"6d",x"68",x"63"),
  1087 => (x"0a",x"3a",x"6b",x"72"),
  1088 => (x"49",x"00",x"0a",x"00"),
  1089 => (x"47",x"5f",x"74",x"6e"),
  1090 => (x"3a",x"62",x"6f",x"6c"),
  1091 => (x"20",x"20",x"20",x"20"),
  1092 => (x"20",x"20",x"20",x"20"),
  1093 => (x"20",x"20",x"20",x"20"),
  1094 => (x"00",x"0a",x"64",x"25"),
  1095 => (x"20",x"20",x"20",x"20"),
  1096 => (x"20",x"20",x"20",x"20"),
  1097 => (x"75",x"6f",x"68",x"73"),
  1098 => (x"62",x"20",x"64",x"6c"),
  1099 => (x"20",x"20",x"3a",x"65"),
  1100 => (x"0a",x"64",x"25",x"20"),
  1101 => (x"6f",x"6f",x"42",x"00"),
  1102 => (x"6c",x"47",x"5f",x"6c"),
  1103 => (x"20",x"3a",x"62",x"6f"),
  1104 => (x"20",x"20",x"20",x"20"),
  1105 => (x"20",x"20",x"20",x"20"),
  1106 => (x"64",x"25",x"20",x"20"),
  1107 => (x"20",x"20",x"00",x"0a"),
  1108 => (x"20",x"20",x"20",x"20"),
  1109 => (x"68",x"73",x"20",x"20"),
  1110 => (x"64",x"6c",x"75",x"6f"),
  1111 => (x"3a",x"65",x"62",x"20"),
  1112 => (x"25",x"20",x"20",x"20"),
  1113 => (x"43",x"00",x"0a",x"64"),
  1114 => (x"5f",x"31",x"5f",x"68"),
  1115 => (x"62",x"6f",x"6c",x"47"),
  1116 => (x"20",x"20",x"20",x"3a"),
  1117 => (x"20",x"20",x"20",x"20"),
  1118 => (x"20",x"20",x"20",x"20"),
  1119 => (x"00",x"0a",x"63",x"25"),
  1120 => (x"20",x"20",x"20",x"20"),
  1121 => (x"20",x"20",x"20",x"20"),
  1122 => (x"75",x"6f",x"68",x"73"),
  1123 => (x"62",x"20",x"64",x"6c"),
  1124 => (x"20",x"20",x"3a",x"65"),
  1125 => (x"0a",x"63",x"25",x"20"),
  1126 => (x"5f",x"68",x"43",x"00"),
  1127 => (x"6c",x"47",x"5f",x"32"),
  1128 => (x"20",x"3a",x"62",x"6f"),
  1129 => (x"20",x"20",x"20",x"20"),
  1130 => (x"20",x"20",x"20",x"20"),
  1131 => (x"63",x"25",x"20",x"20"),
  1132 => (x"20",x"20",x"00",x"0a"),
  1133 => (x"20",x"20",x"20",x"20"),
  1134 => (x"68",x"73",x"20",x"20"),
  1135 => (x"64",x"6c",x"75",x"6f"),
  1136 => (x"3a",x"65",x"62",x"20"),
  1137 => (x"25",x"20",x"20",x"20"),
  1138 => (x"41",x"00",x"0a",x"63"),
  1139 => (x"31",x"5f",x"72",x"72"),
  1140 => (x"6f",x"6c",x"47",x"5f"),
  1141 => (x"5d",x"38",x"5b",x"62"),
  1142 => (x"20",x"20",x"20",x"3a"),
  1143 => (x"20",x"20",x"20",x"20"),
  1144 => (x"00",x"0a",x"64",x"25"),
  1145 => (x"20",x"20",x"20",x"20"),
  1146 => (x"20",x"20",x"20",x"20"),
  1147 => (x"75",x"6f",x"68",x"73"),
  1148 => (x"62",x"20",x"64",x"6c"),
  1149 => (x"20",x"20",x"3a",x"65"),
  1150 => (x"0a",x"64",x"25",x"20"),
  1151 => (x"72",x"72",x"41",x"00"),
  1152 => (x"47",x"5f",x"32",x"5f"),
  1153 => (x"5b",x"62",x"6f",x"6c"),
  1154 => (x"37",x"5b",x"5d",x"38"),
  1155 => (x"20",x"20",x"3a",x"5d"),
  1156 => (x"64",x"25",x"20",x"20"),
  1157 => (x"20",x"20",x"00",x"0a"),
  1158 => (x"20",x"20",x"20",x"20"),
  1159 => (x"68",x"73",x"20",x"20"),
  1160 => (x"64",x"6c",x"75",x"6f"),
  1161 => (x"3a",x"65",x"62",x"20"),
  1162 => (x"4e",x"20",x"20",x"20"),
  1163 => (x"65",x"62",x"6d",x"75"),
  1164 => (x"66",x"4f",x"5f",x"72"),
  1165 => (x"6e",x"75",x"52",x"5f"),
  1166 => (x"20",x"2b",x"20",x"73"),
  1167 => (x"00",x"0a",x"30",x"31"),
  1168 => (x"5f",x"72",x"74",x"50"),
  1169 => (x"62",x"6f",x"6c",x"47"),
  1170 => (x"00",x"0a",x"3e",x"2d"),
  1171 => (x"74",x"50",x"20",x"20"),
  1172 => (x"6f",x"43",x"5f",x"72"),
  1173 => (x"20",x"3a",x"70",x"6d"),
  1174 => (x"20",x"20",x"20",x"20"),
  1175 => (x"20",x"20",x"20",x"20"),
  1176 => (x"0a",x"64",x"25",x"20"),
  1177 => (x"20",x"20",x"20",x"00"),
  1178 => (x"20",x"20",x"20",x"20"),
  1179 => (x"6f",x"68",x"73",x"20"),
  1180 => (x"20",x"64",x"6c",x"75"),
  1181 => (x"20",x"3a",x"65",x"62"),
  1182 => (x"69",x"28",x"20",x"20"),
  1183 => (x"65",x"6c",x"70",x"6d"),
  1184 => (x"74",x"6e",x"65",x"6d"),
  1185 => (x"6f",x"69",x"74",x"61"),
  1186 => (x"65",x"64",x"2d",x"6e"),
  1187 => (x"64",x"6e",x"65",x"70"),
  1188 => (x"29",x"74",x"6e",x"65"),
  1189 => (x"20",x"20",x"00",x"0a"),
  1190 => (x"63",x"73",x"69",x"44"),
  1191 => (x"20",x"20",x"3a",x"72"),
  1192 => (x"20",x"20",x"20",x"20"),
  1193 => (x"20",x"20",x"20",x"20"),
  1194 => (x"25",x"20",x"20",x"20"),
  1195 => (x"20",x"00",x"0a",x"64"),
  1196 => (x"20",x"20",x"20",x"20"),
  1197 => (x"73",x"20",x"20",x"20"),
  1198 => (x"6c",x"75",x"6f",x"68"),
  1199 => (x"65",x"62",x"20",x"64"),
  1200 => (x"20",x"20",x"20",x"3a"),
  1201 => (x"00",x"0a",x"64",x"25"),
  1202 => (x"6e",x"45",x"20",x"20"),
  1203 => (x"43",x"5f",x"6d",x"75"),
  1204 => (x"3a",x"70",x"6d",x"6f"),
  1205 => (x"20",x"20",x"20",x"20"),
  1206 => (x"20",x"20",x"20",x"20"),
  1207 => (x"0a",x"64",x"25",x"20"),
  1208 => (x"20",x"20",x"20",x"00"),
  1209 => (x"20",x"20",x"20",x"20"),
  1210 => (x"6f",x"68",x"73",x"20"),
  1211 => (x"20",x"64",x"6c",x"75"),
  1212 => (x"20",x"3a",x"65",x"62"),
  1213 => (x"64",x"25",x"20",x"20"),
  1214 => (x"20",x"20",x"00",x"0a"),
  1215 => (x"5f",x"74",x"6e",x"49"),
  1216 => (x"70",x"6d",x"6f",x"43"),
  1217 => (x"20",x"20",x"20",x"3a"),
  1218 => (x"20",x"20",x"20",x"20"),
  1219 => (x"25",x"20",x"20",x"20"),
  1220 => (x"20",x"00",x"0a",x"64"),
  1221 => (x"20",x"20",x"20",x"20"),
  1222 => (x"73",x"20",x"20",x"20"),
  1223 => (x"6c",x"75",x"6f",x"68"),
  1224 => (x"65",x"62",x"20",x"64"),
  1225 => (x"20",x"20",x"20",x"3a"),
  1226 => (x"00",x"0a",x"64",x"25"),
  1227 => (x"74",x"53",x"20",x"20"),
  1228 => (x"6f",x"43",x"5f",x"72"),
  1229 => (x"20",x"3a",x"70",x"6d"),
  1230 => (x"20",x"20",x"20",x"20"),
  1231 => (x"20",x"20",x"20",x"20"),
  1232 => (x"0a",x"73",x"25",x"20"),
  1233 => (x"20",x"20",x"20",x"00"),
  1234 => (x"20",x"20",x"20",x"20"),
  1235 => (x"6f",x"68",x"73",x"20"),
  1236 => (x"20",x"64",x"6c",x"75"),
  1237 => (x"20",x"3a",x"65",x"62"),
  1238 => (x"48",x"44",x"20",x"20"),
  1239 => (x"54",x"53",x"59",x"52"),
  1240 => (x"20",x"45",x"4e",x"4f"),
  1241 => (x"47",x"4f",x"52",x"50"),
  1242 => (x"2c",x"4d",x"41",x"52"),
  1243 => (x"4d",x"4f",x"53",x"20"),
  1244 => (x"54",x"53",x"20",x"45"),
  1245 => (x"47",x"4e",x"49",x"52"),
  1246 => (x"65",x"4e",x"00",x"0a"),
  1247 => (x"50",x"5f",x"74",x"78"),
  1248 => (x"47",x"5f",x"72",x"74"),
  1249 => (x"2d",x"62",x"6f",x"6c"),
  1250 => (x"20",x"00",x"0a",x"3e"),
  1251 => (x"72",x"74",x"50",x"20"),
  1252 => (x"6d",x"6f",x"43",x"5f"),
  1253 => (x"20",x"20",x"3a",x"70"),
  1254 => (x"20",x"20",x"20",x"20"),
  1255 => (x"20",x"20",x"20",x"20"),
  1256 => (x"00",x"0a",x"64",x"25"),
  1257 => (x"20",x"20",x"20",x"20"),
  1258 => (x"20",x"20",x"20",x"20"),
  1259 => (x"75",x"6f",x"68",x"73"),
  1260 => (x"62",x"20",x"64",x"6c"),
  1261 => (x"20",x"20",x"3a",x"65"),
  1262 => (x"6d",x"69",x"28",x"20"),
  1263 => (x"6d",x"65",x"6c",x"70"),
  1264 => (x"61",x"74",x"6e",x"65"),
  1265 => (x"6e",x"6f",x"69",x"74"),
  1266 => (x"70",x"65",x"64",x"2d"),
  1267 => (x"65",x"64",x"6e",x"65"),
  1268 => (x"2c",x"29",x"74",x"6e"),
  1269 => (x"6d",x"61",x"73",x"20"),
  1270 => (x"73",x"61",x"20",x"65"),
  1271 => (x"6f",x"62",x"61",x"20"),
  1272 => (x"00",x"0a",x"65",x"76"),
  1273 => (x"69",x"44",x"20",x"20"),
  1274 => (x"3a",x"72",x"63",x"73"),
  1275 => (x"20",x"20",x"20",x"20"),
  1276 => (x"20",x"20",x"20",x"20"),
  1277 => (x"20",x"20",x"20",x"20"),
  1278 => (x"0a",x"64",x"25",x"20"),
  1279 => (x"20",x"20",x"20",x"00"),
  1280 => (x"20",x"20",x"20",x"20"),
  1281 => (x"6f",x"68",x"73",x"20"),
  1282 => (x"20",x"64",x"6c",x"75"),
  1283 => (x"20",x"3a",x"65",x"62"),
  1284 => (x"64",x"25",x"20",x"20"),
  1285 => (x"20",x"20",x"00",x"0a"),
  1286 => (x"6d",x"75",x"6e",x"45"),
  1287 => (x"6d",x"6f",x"43",x"5f"),
  1288 => (x"20",x"20",x"3a",x"70"),
  1289 => (x"20",x"20",x"20",x"20"),
  1290 => (x"25",x"20",x"20",x"20"),
  1291 => (x"20",x"00",x"0a",x"64"),
  1292 => (x"20",x"20",x"20",x"20"),
  1293 => (x"73",x"20",x"20",x"20"),
  1294 => (x"6c",x"75",x"6f",x"68"),
  1295 => (x"65",x"62",x"20",x"64"),
  1296 => (x"20",x"20",x"20",x"3a"),
  1297 => (x"00",x"0a",x"64",x"25"),
  1298 => (x"6e",x"49",x"20",x"20"),
  1299 => (x"6f",x"43",x"5f",x"74"),
  1300 => (x"20",x"3a",x"70",x"6d"),
  1301 => (x"20",x"20",x"20",x"20"),
  1302 => (x"20",x"20",x"20",x"20"),
  1303 => (x"0a",x"64",x"25",x"20"),
  1304 => (x"20",x"20",x"20",x"00"),
  1305 => (x"20",x"20",x"20",x"20"),
  1306 => (x"6f",x"68",x"73",x"20"),
  1307 => (x"20",x"64",x"6c",x"75"),
  1308 => (x"20",x"3a",x"65",x"62"),
  1309 => (x"64",x"25",x"20",x"20"),
  1310 => (x"20",x"20",x"00",x"0a"),
  1311 => (x"5f",x"72",x"74",x"53"),
  1312 => (x"70",x"6d",x"6f",x"43"),
  1313 => (x"20",x"20",x"20",x"3a"),
  1314 => (x"20",x"20",x"20",x"20"),
  1315 => (x"25",x"20",x"20",x"20"),
  1316 => (x"20",x"00",x"0a",x"73"),
  1317 => (x"20",x"20",x"20",x"20"),
  1318 => (x"73",x"20",x"20",x"20"),
  1319 => (x"6c",x"75",x"6f",x"68"),
  1320 => (x"65",x"62",x"20",x"64"),
  1321 => (x"20",x"20",x"20",x"3a"),
  1322 => (x"59",x"52",x"48",x"44"),
  1323 => (x"4e",x"4f",x"54",x"53"),
  1324 => (x"52",x"50",x"20",x"45"),
  1325 => (x"41",x"52",x"47",x"4f"),
  1326 => (x"53",x"20",x"2c",x"4d"),
  1327 => (x"20",x"45",x"4d",x"4f"),
  1328 => (x"49",x"52",x"54",x"53"),
  1329 => (x"00",x"0a",x"47",x"4e"),
  1330 => (x"5f",x"74",x"6e",x"49"),
  1331 => (x"6f",x"4c",x"5f",x"31"),
  1332 => (x"20",x"20",x"3a",x"63"),
  1333 => (x"20",x"20",x"20",x"20"),
  1334 => (x"20",x"20",x"20",x"20"),
  1335 => (x"0a",x"64",x"25",x"20"),
  1336 => (x"20",x"20",x"20",x"00"),
  1337 => (x"20",x"20",x"20",x"20"),
  1338 => (x"6f",x"68",x"73",x"20"),
  1339 => (x"20",x"64",x"6c",x"75"),
  1340 => (x"20",x"3a",x"65",x"62"),
  1341 => (x"64",x"25",x"20",x"20"),
  1342 => (x"6e",x"49",x"00",x"0a"),
  1343 => (x"5f",x"32",x"5f",x"74"),
  1344 => (x"3a",x"63",x"6f",x"4c"),
  1345 => (x"20",x"20",x"20",x"20"),
  1346 => (x"20",x"20",x"20",x"20"),
  1347 => (x"25",x"20",x"20",x"20"),
  1348 => (x"20",x"00",x"0a",x"64"),
  1349 => (x"20",x"20",x"20",x"20"),
  1350 => (x"73",x"20",x"20",x"20"),
  1351 => (x"6c",x"75",x"6f",x"68"),
  1352 => (x"65",x"62",x"20",x"64"),
  1353 => (x"20",x"20",x"20",x"3a"),
  1354 => (x"00",x"0a",x"64",x"25"),
  1355 => (x"5f",x"74",x"6e",x"49"),
  1356 => (x"6f",x"4c",x"5f",x"33"),
  1357 => (x"20",x"20",x"3a",x"63"),
  1358 => (x"20",x"20",x"20",x"20"),
  1359 => (x"20",x"20",x"20",x"20"),
  1360 => (x"0a",x"64",x"25",x"20"),
  1361 => (x"20",x"20",x"20",x"00"),
  1362 => (x"20",x"20",x"20",x"20"),
  1363 => (x"6f",x"68",x"73",x"20"),
  1364 => (x"20",x"64",x"6c",x"75"),
  1365 => (x"20",x"3a",x"65",x"62"),
  1366 => (x"64",x"25",x"20",x"20"),
  1367 => (x"6e",x"45",x"00",x"0a"),
  1368 => (x"4c",x"5f",x"6d",x"75"),
  1369 => (x"20",x"3a",x"63",x"6f"),
  1370 => (x"20",x"20",x"20",x"20"),
  1371 => (x"20",x"20",x"20",x"20"),
  1372 => (x"25",x"20",x"20",x"20"),
  1373 => (x"20",x"00",x"0a",x"64"),
  1374 => (x"20",x"20",x"20",x"20"),
  1375 => (x"73",x"20",x"20",x"20"),
  1376 => (x"6c",x"75",x"6f",x"68"),
  1377 => (x"65",x"62",x"20",x"64"),
  1378 => (x"20",x"20",x"20",x"3a"),
  1379 => (x"00",x"0a",x"64",x"25"),
  1380 => (x"5f",x"72",x"74",x"53"),
  1381 => (x"6f",x"4c",x"5f",x"31"),
  1382 => (x"20",x"20",x"3a",x"63"),
  1383 => (x"20",x"20",x"20",x"20"),
  1384 => (x"20",x"20",x"20",x"20"),
  1385 => (x"0a",x"73",x"25",x"20"),
  1386 => (x"20",x"20",x"20",x"00"),
  1387 => (x"20",x"20",x"20",x"20"),
  1388 => (x"6f",x"68",x"73",x"20"),
  1389 => (x"20",x"64",x"6c",x"75"),
  1390 => (x"20",x"3a",x"65",x"62"),
  1391 => (x"48",x"44",x"20",x"20"),
  1392 => (x"54",x"53",x"59",x"52"),
  1393 => (x"20",x"45",x"4e",x"4f"),
  1394 => (x"47",x"4f",x"52",x"50"),
  1395 => (x"2c",x"4d",x"41",x"52"),
  1396 => (x"53",x"27",x"31",x"20"),
  1397 => (x"54",x"53",x"20",x"54"),
  1398 => (x"47",x"4e",x"49",x"52"),
  1399 => (x"74",x"53",x"00",x"0a"),
  1400 => (x"5f",x"32",x"5f",x"72"),
  1401 => (x"3a",x"63",x"6f",x"4c"),
  1402 => (x"20",x"20",x"20",x"20"),
  1403 => (x"20",x"20",x"20",x"20"),
  1404 => (x"25",x"20",x"20",x"20"),
  1405 => (x"20",x"00",x"0a",x"73"),
  1406 => (x"20",x"20",x"20",x"20"),
  1407 => (x"73",x"20",x"20",x"20"),
  1408 => (x"6c",x"75",x"6f",x"68"),
  1409 => (x"65",x"62",x"20",x"64"),
  1410 => (x"20",x"20",x"20",x"3a"),
  1411 => (x"59",x"52",x"48",x"44"),
  1412 => (x"4e",x"4f",x"54",x"53"),
  1413 => (x"52",x"50",x"20",x"45"),
  1414 => (x"41",x"52",x"47",x"4f"),
  1415 => (x"32",x"20",x"2c",x"4d"),
  1416 => (x"20",x"44",x"4e",x"27"),
  1417 => (x"49",x"52",x"54",x"53"),
  1418 => (x"00",x"0a",x"47",x"4e"),
  1419 => (x"73",x"55",x"00",x"0a"),
  1420 => (x"74",x"20",x"72",x"65"),
  1421 => (x"3a",x"65",x"6d",x"69"),
  1422 => (x"0a",x"64",x"25",x"20"),
  1423 => (x"00",x"00",x"00",x"00"),
  1424 => (x"00",x"00",x"00",x"00"),
  1425 => (x"00",x"00",x"61",x"a8"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
