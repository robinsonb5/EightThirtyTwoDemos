
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"d4",x"01"),
     1 => (x"18",x"0e",x"87",x"d7"),
     2 => (x"3e",x"27",x"0e",x"1e"),
     3 => (x"0f",x"00",x"00",x"00"),
     4 => (x"80",x"ff",x"48",x"26"),
     5 => (x"27",x"4f",x"08",x"26"),
     6 => (x"00",x"00",x"00",x"23"),
     7 => (x"00",x"30",x"27",x"4f"),
     8 => (x"c2",x"4f",x"00",x"00"),
     9 => (x"27",x"4e",x"c0",x"c0"),
    10 => (x"00",x"00",x"04",x"fe"),
    11 => (x"87",x"fd",x"00",x"0f"),
    12 => (x"4e",x"c0",x"f0",x"c1"),
    13 => (x"00",x"00",x"3d",x"27"),
    14 => (x"fd",x"00",x"0f",x"00"),
    15 => (x"1e",x"4f",x"4f",x"87"),
    16 => (x"ff",x"1e",x"1e",x"72"),
    17 => (x"48",x"6a",x"4a",x"c0"),
    18 => (x"c4",x"98",x"c0",x"c4"),
    19 => (x"02",x"6e",x"58",x"a6"),
    20 => (x"cc",x"87",x"f3",x"ff"),
    21 => (x"66",x"cc",x"7a",x"66"),
    22 => (x"4a",x"26",x"26",x"48"),
    23 => (x"5e",x"0e",x"4f",x"26"),
    24 => (x"5d",x"5c",x"5b",x"5a"),
    25 => (x"4b",x"66",x"d4",x"0e"),
    26 => (x"4c",x"13",x"4d",x"c0"),
    27 => (x"c0",x"02",x"9c",x"74"),
    28 => (x"4a",x"74",x"87",x"d6"),
    29 => (x"3f",x"27",x"1e",x"72"),
    30 => (x"0f",x"00",x"00",x"00"),
    31 => (x"85",x"c1",x"86",x"c4"),
    32 => (x"9c",x"74",x"4c",x"13"),
    33 => (x"87",x"ea",x"ff",x"05"),
    34 => (x"4d",x"26",x"48",x"75"),
    35 => (x"4b",x"26",x"4c",x"26"),
    36 => (x"4f",x"26",x"4a",x"26"),
    37 => (x"5b",x"5a",x"5e",x"0e"),
    38 => (x"1e",x"0e",x"5d",x"5c"),
    39 => (x"76",x"4d",x"66",x"d8"),
    40 => (x"c0",x"79",x"c0",x"49"),
    41 => (x"c0",x"03",x"ad",x"b7"),
    42 => (x"ed",x"c0",x"87",x"cd"),
    43 => (x"00",x"3f",x"27",x"1e"),
    44 => (x"c4",x"0f",x"00",x"00"),
    45 => (x"75",x"8d",x"0d",x"86"),
    46 => (x"c2",x"c1",x"02",x"9d"),
    47 => (x"75",x"4c",x"c0",x"87"),
    48 => (x"2a",x"b7",x"dc",x"4a"),
    49 => (x"9b",x"cf",x"4b",x"72"),
    50 => (x"9b",x"73",x"35",x"c4"),
    51 => (x"87",x"c4",x"c0",x"02"),
    52 => (x"79",x"c1",x"49",x"76"),
    53 => (x"06",x"ab",x"b7",x"c9"),
    54 => (x"c0",x"87",x"c6",x"c0"),
    55 => (x"c3",x"c0",x"83",x"f7"),
    56 => (x"83",x"f0",x"c0",x"87"),
    57 => (x"ca",x"c0",x"02",x"6e"),
    58 => (x"27",x"1e",x"73",x"87"),
    59 => (x"00",x"00",x"00",x"3f"),
    60 => (x"c1",x"86",x"c4",x"0f"),
    61 => (x"ac",x"b7",x"c8",x"84"),
    62 => (x"87",x"c3",x"ff",x"04"),
    63 => (x"c0",x"87",x"cb",x"c0"),
    64 => (x"3f",x"27",x"1e",x"f0"),
    65 => (x"0f",x"00",x"00",x"00"),
    66 => (x"48",x"c0",x"86",x"c4"),
    67 => (x"26",x"4d",x"26",x"26"),
    68 => (x"26",x"4b",x"26",x"4c"),
    69 => (x"0e",x"4f",x"26",x"4a"),
    70 => (x"5c",x"5b",x"5a",x"5e"),
    71 => (x"c0",x"1e",x"0e",x"5d"),
    72 => (x"c0",x"49",x"76",x"4c"),
    73 => (x"4b",x"a6",x"dc",x"79"),
    74 => (x"d8",x"4a",x"66",x"d8"),
    75 => (x"80",x"c1",x"48",x"66"),
    76 => (x"12",x"58",x"a6",x"dc"),
    77 => (x"c0",x"c0",x"c1",x"4d"),
    78 => (x"c4",x"95",x"c0",x"c0"),
    79 => (x"4d",x"95",x"b7",x"c0"),
    80 => (x"c4",x"02",x"9d",x"75"),
    81 => (x"02",x"6e",x"87",x"d2"),
    82 => (x"76",x"87",x"d7",x"c3"),
    83 => (x"75",x"79",x"c0",x"49"),
    84 => (x"ad",x"e3",x"c1",x"4a"),
    85 => (x"87",x"dd",x"c2",x"02"),
    86 => (x"02",x"aa",x"e4",x"c1"),
    87 => (x"c1",x"87",x"d8",x"c0"),
    88 => (x"c2",x"02",x"aa",x"ec"),
    89 => (x"f3",x"c1",x"87",x"c8"),
    90 => (x"e8",x"c1",x"02",x"aa"),
    91 => (x"aa",x"f8",x"c1",x"87"),
    92 => (x"87",x"f2",x"c0",x"02"),
    93 => (x"ca",x"87",x"d3",x"c2"),
    94 => (x"16",x"50",x"27",x"1e"),
    95 => (x"c4",x"1e",x"00",x"00"),
    96 => (x"c4",x"4a",x"73",x"83"),
    97 => (x"27",x"1e",x"6a",x"8a"),
    98 => (x"00",x"00",x"00",x"94"),
    99 => (x"70",x"86",x"cc",x"0f"),
   100 => (x"72",x"4c",x"74",x"4a"),
   101 => (x"16",x"50",x"27",x"84"),
   102 => (x"27",x"1e",x"00",x"00"),
   103 => (x"00",x"00",x"00",x"5e"),
   104 => (x"c2",x"86",x"c4",x"0f"),
   105 => (x"1e",x"d0",x"87",x"d4"),
   106 => (x"00",x"16",x"50",x"27"),
   107 => (x"83",x"c4",x"1e",x"00"),
   108 => (x"8a",x"c4",x"4a",x"73"),
   109 => (x"94",x"27",x"1e",x"6a"),
   110 => (x"0f",x"00",x"00",x"00"),
   111 => (x"4a",x"70",x"86",x"cc"),
   112 => (x"84",x"72",x"4c",x"74"),
   113 => (x"00",x"16",x"50",x"27"),
   114 => (x"5e",x"27",x"1e",x"00"),
   115 => (x"0f",x"00",x"00",x"00"),
   116 => (x"e5",x"c1",x"86",x"c4"),
   117 => (x"73",x"83",x"c4",x"87"),
   118 => (x"6a",x"8a",x"c4",x"4a"),
   119 => (x"00",x"5e",x"27",x"1e"),
   120 => (x"c4",x"0f",x"00",x"00"),
   121 => (x"74",x"4a",x"70",x"86"),
   122 => (x"c1",x"84",x"72",x"4c"),
   123 => (x"49",x"76",x"87",x"cc"),
   124 => (x"c5",x"c1",x"79",x"c1"),
   125 => (x"73",x"83",x"c4",x"87"),
   126 => (x"6a",x"8a",x"c4",x"4a"),
   127 => (x"00",x"3f",x"27",x"1e"),
   128 => (x"c4",x"0f",x"00",x"00"),
   129 => (x"c0",x"84",x"c1",x"86"),
   130 => (x"e5",x"c0",x"87",x"f0"),
   131 => (x"00",x"3f",x"27",x"1e"),
   132 => (x"c4",x"0f",x"00",x"00"),
   133 => (x"27",x"1e",x"75",x"86"),
   134 => (x"00",x"00",x"00",x"3f"),
   135 => (x"c0",x"86",x"c4",x"0f"),
   136 => (x"e5",x"c0",x"87",x"d8"),
   137 => (x"c7",x"c0",x"05",x"ad"),
   138 => (x"c1",x"49",x"76",x"87"),
   139 => (x"87",x"ca",x"c0",x"79"),
   140 => (x"3f",x"27",x"1e",x"75"),
   141 => (x"0f",x"00",x"00",x"00"),
   142 => (x"66",x"d8",x"86",x"c4"),
   143 => (x"48",x"66",x"d8",x"4a"),
   144 => (x"a6",x"dc",x"80",x"c1"),
   145 => (x"c1",x"4d",x"12",x"58"),
   146 => (x"c0",x"c0",x"c0",x"c0"),
   147 => (x"b7",x"c0",x"c4",x"95"),
   148 => (x"9d",x"75",x"4d",x"95"),
   149 => (x"87",x"ee",x"fb",x"05"),
   150 => (x"26",x"26",x"48",x"74"),
   151 => (x"26",x"4c",x"26",x"4d"),
   152 => (x"26",x"4a",x"26",x"4b"),
   153 => (x"5a",x"5e",x"0e",x"4f"),
   154 => (x"66",x"d0",x"0e",x"5b"),
   155 => (x"7b",x"66",x"cc",x"4b"),
   156 => (x"27",x"1e",x"66",x"cc"),
   157 => (x"00",x"00",x"04",x"8c"),
   158 => (x"70",x"86",x"c4",x"0f"),
   159 => (x"05",x"9a",x"72",x"4a"),
   160 => (x"c3",x"87",x"c2",x"c0"),
   161 => (x"4a",x"66",x"cc",x"7b"),
   162 => (x"c0",x"49",x"66",x"cc"),
   163 => (x"c0",x"02",x"a9",x"b7"),
   164 => (x"b7",x"c1",x"87",x"df"),
   165 => (x"dd",x"c0",x"02",x"aa"),
   166 => (x"aa",x"b7",x"c2",x"87"),
   167 => (x"87",x"ef",x"c0",x"02"),
   168 => (x"02",x"aa",x"b7",x"c3"),
   169 => (x"c4",x"87",x"ef",x"c0"),
   170 => (x"c0",x"02",x"aa",x"b7"),
   171 => (x"e5",x"c0",x"87",x"e6"),
   172 => (x"c0",x"7b",x"c0",x"87"),
   173 => (x"78",x"27",x"87",x"e0"),
   174 => (x"bf",x"00",x"00",x"16"),
   175 => (x"b7",x"e4",x"c1",x"49"),
   176 => (x"c5",x"c0",x"06",x"a9"),
   177 => (x"c0",x"7b",x"c0",x"87"),
   178 => (x"7b",x"c3",x"87",x"cc"),
   179 => (x"c1",x"87",x"c7",x"c0"),
   180 => (x"87",x"c2",x"c0",x"7b"),
   181 => (x"4b",x"26",x"7b",x"c2"),
   182 => (x"4f",x"26",x"4a",x"26"),
   183 => (x"c8",x"1e",x"72",x"1e"),
   184 => (x"82",x"c2",x"4a",x"66"),
   185 => (x"72",x"48",x"66",x"cc"),
   186 => (x"49",x"66",x"d0",x"80"),
   187 => (x"4a",x"26",x"79",x"70"),
   188 => (x"5e",x"0e",x"4f",x"26"),
   189 => (x"5d",x"5c",x"5b",x"5a"),
   190 => (x"4d",x"66",x"dc",x"0e"),
   191 => (x"4a",x"75",x"85",x"c5"),
   192 => (x"4a",x"72",x"92",x"c4"),
   193 => (x"c0",x"82",x"66",x"d4"),
   194 => (x"72",x"7a",x"66",x"e0"),
   195 => (x"6a",x"83",x"c4",x"4b"),
   196 => (x"82",x"f8",x"c1",x"7b"),
   197 => (x"4c",x"75",x"7a",x"75"),
   198 => (x"82",x"c1",x"4a",x"75"),
   199 => (x"01",x"ad",x"b7",x"72"),
   200 => (x"75",x"87",x"e1",x"c0"),
   201 => (x"93",x"c8",x"c3",x"4b"),
   202 => (x"66",x"d8",x"4b",x"73"),
   203 => (x"c4",x"4a",x"74",x"83"),
   204 => (x"73",x"4a",x"72",x"92"),
   205 => (x"c1",x"7a",x"75",x"82"),
   206 => (x"c1",x"4a",x"75",x"84"),
   207 => (x"ac",x"b7",x"72",x"82"),
   208 => (x"87",x"df",x"ff",x"06"),
   209 => (x"c8",x"c3",x"4c",x"75"),
   210 => (x"d8",x"4c",x"74",x"94"),
   211 => (x"4a",x"75",x"84",x"66"),
   212 => (x"4b",x"74",x"92",x"c4"),
   213 => (x"8b",x"c4",x"83",x"72"),
   214 => (x"80",x"c1",x"48",x"6b"),
   215 => (x"66",x"d4",x"7b",x"70"),
   216 => (x"c0",x"83",x"72",x"4b"),
   217 => (x"72",x"84",x"e0",x"fe"),
   218 => (x"6b",x"82",x"74",x"4a"),
   219 => (x"16",x"78",x"27",x"7a"),
   220 => (x"c5",x"49",x"00",x"00"),
   221 => (x"26",x"4d",x"26",x"79"),
   222 => (x"26",x"4b",x"26",x"4c"),
   223 => (x"0e",x"4f",x"26",x"4a"),
   224 => (x"5c",x"5b",x"5a",x"5e"),
   225 => (x"66",x"d0",x"97",x"0e"),
   226 => (x"c1",x"4b",x"74",x"4c"),
   227 => (x"c0",x"c0",x"c0",x"c0"),
   228 => (x"b7",x"c0",x"c4",x"93"),
   229 => (x"d4",x"97",x"4b",x"93"),
   230 => (x"c0",x"c1",x"4a",x"66"),
   231 => (x"92",x"c0",x"c0",x"c0"),
   232 => (x"92",x"b7",x"c0",x"c4"),
   233 => (x"ab",x"b7",x"72",x"4a"),
   234 => (x"87",x"c5",x"c0",x"02"),
   235 => (x"ca",x"c0",x"48",x"c0"),
   236 => (x"16",x"80",x"27",x"87"),
   237 => (x"74",x"49",x"00",x"00"),
   238 => (x"26",x"48",x"c1",x"51"),
   239 => (x"26",x"4b",x"26",x"4c"),
   240 => (x"0e",x"4f",x"26",x"4a"),
   241 => (x"5c",x"5b",x"5a",x"5e"),
   242 => (x"6e",x"97",x"1e",x"0e"),
   243 => (x"d8",x"4b",x"c2",x"4c"),
   244 => (x"82",x"c1",x"4a",x"66"),
   245 => (x"6a",x"97",x"82",x"73"),
   246 => (x"c0",x"c0",x"c1",x"4a"),
   247 => (x"c4",x"92",x"c0",x"c0"),
   248 => (x"4a",x"92",x"b7",x"c0"),
   249 => (x"66",x"d8",x"1e",x"72"),
   250 => (x"97",x"82",x"73",x"4a"),
   251 => (x"c0",x"c1",x"4a",x"6a"),
   252 => (x"92",x"c0",x"c0",x"c0"),
   253 => (x"92",x"b7",x"c0",x"c4"),
   254 => (x"27",x"1e",x"72",x"4a"),
   255 => (x"00",x"00",x"03",x"7f"),
   256 => (x"70",x"86",x"c8",x"0f"),
   257 => (x"05",x"9a",x"72",x"4a"),
   258 => (x"c1",x"87",x"c5",x"c0"),
   259 => (x"83",x"c1",x"4c",x"c1"),
   260 => (x"06",x"ab",x"b7",x"c2"),
   261 => (x"74",x"87",x"f8",x"fe"),
   262 => (x"c0",x"c0",x"c1",x"4a"),
   263 => (x"c4",x"92",x"c0",x"c0"),
   264 => (x"4a",x"92",x"b7",x"c0"),
   265 => (x"aa",x"b7",x"d7",x"c1"),
   266 => (x"87",x"d7",x"c0",x"04"),
   267 => (x"c0",x"c1",x"4a",x"74"),
   268 => (x"92",x"c0",x"c0",x"c0"),
   269 => (x"92",x"b7",x"c0",x"c4"),
   270 => (x"b7",x"da",x"c1",x"4a"),
   271 => (x"c2",x"c0",x"03",x"aa"),
   272 => (x"74",x"4b",x"c7",x"87"),
   273 => (x"c0",x"c0",x"c1",x"4a"),
   274 => (x"c4",x"92",x"c0",x"c0"),
   275 => (x"4a",x"92",x"b7",x"c0"),
   276 => (x"aa",x"b7",x"d2",x"c1"),
   277 => (x"87",x"c5",x"c0",x"05"),
   278 => (x"e6",x"c0",x"48",x"c1"),
   279 => (x"4a",x"66",x"d4",x"87"),
   280 => (x"27",x"49",x"66",x"d8"),
   281 => (x"00",x"00",x"04",x"ea"),
   282 => (x"c0",x"4a",x"70",x"0f"),
   283 => (x"c0",x"06",x"aa",x"b7"),
   284 => (x"48",x"73",x"87",x"cf"),
   285 => (x"7c",x"27",x"80",x"c7"),
   286 => (x"58",x"00",x"00",x"16"),
   287 => (x"c2",x"c0",x"48",x"c1"),
   288 => (x"26",x"48",x"c0",x"87"),
   289 => (x"4b",x"26",x"4c",x"26"),
   290 => (x"4f",x"26",x"4a",x"26"),
   291 => (x"49",x"66",x"c4",x"1e"),
   292 => (x"05",x"a9",x"b7",x"c2"),
   293 => (x"c1",x"87",x"c5",x"c0"),
   294 => (x"87",x"c2",x"c0",x"48"),
   295 => (x"4f",x"26",x"48",x"c0"),
   296 => (x"72",x"1e",x"73",x"1e"),
   297 => (x"87",x"d9",x"02",x"9a"),
   298 => (x"4b",x"c1",x"48",x"c0"),
   299 => (x"82",x"01",x"a9",x"72"),
   300 => (x"87",x"f8",x"83",x"73"),
   301 => (x"89",x"03",x"a9",x"72"),
   302 => (x"c1",x"07",x"80",x"73"),
   303 => (x"f3",x"05",x"2b",x"2a"),
   304 => (x"26",x"4b",x"26",x"87"),
   305 => (x"1e",x"75",x"1e",x"4f"),
   306 => (x"a1",x"71",x"4d",x"c0"),
   307 => (x"c1",x"b9",x"ff",x"04"),
   308 => (x"72",x"07",x"bd",x"81"),
   309 => (x"ba",x"ff",x"04",x"a2"),
   310 => (x"07",x"bd",x"82",x"c1"),
   311 => (x"9d",x"75",x"87",x"c2"),
   312 => (x"c1",x"b8",x"ff",x"05"),
   313 => (x"4d",x"25",x"07",x"80"),
   314 => (x"12",x"1e",x"4f",x"26"),
   315 => (x"c4",x"02",x"11",x"48"),
   316 => (x"f6",x"02",x"88",x"87"),
   317 => (x"1e",x"4f",x"26",x"87"),
   318 => (x"48",x"bf",x"c8",x"ff"),
   319 => (x"5e",x"0e",x"4f",x"26"),
   320 => (x"5d",x"5c",x"5b",x"5a"),
   321 => (x"c4",x"8e",x"d0",x"0e"),
   322 => (x"74",x"27",x"4c",x"66"),
   323 => (x"49",x"00",x"00",x"16"),
   324 => (x"00",x"3e",x"78",x"27"),
   325 => (x"70",x"27",x"79",x"00"),
   326 => (x"49",x"00",x"00",x"16"),
   327 => (x"00",x"3e",x"a8",x"27"),
   328 => (x"a8",x"27",x"79",x"00"),
   329 => (x"49",x"00",x"00",x"3e"),
   330 => (x"00",x"3e",x"78",x"27"),
   331 => (x"ac",x"27",x"79",x"00"),
   332 => (x"49",x"00",x"00",x"3e"),
   333 => (x"b0",x"27",x"79",x"c0"),
   334 => (x"49",x"00",x"00",x"3e"),
   335 => (x"b4",x"27",x"79",x"c2"),
   336 => (x"49",x"00",x"00",x"3e"),
   337 => (x"27",x"79",x"e8",x"c0"),
   338 => (x"00",x"00",x"3e",x"b8"),
   339 => (x"0f",x"d1",x"27",x"49"),
   340 => (x"72",x"48",x"00",x"00"),
   341 => (x"20",x"41",x"20",x"1e"),
   342 => (x"20",x"41",x"20",x"41"),
   343 => (x"20",x"41",x"20",x"41"),
   344 => (x"10",x"41",x"20",x"41"),
   345 => (x"10",x"51",x"10",x"51"),
   346 => (x"27",x"4a",x"26",x"51"),
   347 => (x"00",x"00",x"3e",x"d8"),
   348 => (x"0f",x"f0",x"27",x"49"),
   349 => (x"72",x"48",x"00",x"00"),
   350 => (x"20",x"41",x"20",x"1e"),
   351 => (x"20",x"41",x"20",x"41"),
   352 => (x"20",x"41",x"20",x"41"),
   353 => (x"10",x"41",x"20",x"41"),
   354 => (x"10",x"51",x"10",x"51"),
   355 => (x"27",x"4a",x"26",x"51"),
   356 => (x"00",x"00",x"1d",x"ac"),
   357 => (x"27",x"79",x"ca",x"49"),
   358 => (x"00",x"00",x"10",x"0f"),
   359 => (x"01",x"17",x"27",x"1e"),
   360 => (x"c4",x"0f",x"00",x"00"),
   361 => (x"10",x"11",x"27",x"86"),
   362 => (x"27",x"1e",x"00",x"00"),
   363 => (x"00",x"00",x"01",x"17"),
   364 => (x"27",x"86",x"c4",x"0f"),
   365 => (x"00",x"00",x"10",x"41"),
   366 => (x"01",x"17",x"27",x"1e"),
   367 => (x"c4",x"0f",x"00",x"00"),
   368 => (x"15",x"f4",x"27",x"86"),
   369 => (x"02",x"bf",x"00",x"00"),
   370 => (x"27",x"87",x"df",x"c0"),
   371 => (x"00",x"00",x"0e",x"58"),
   372 => (x"01",x"17",x"27",x"1e"),
   373 => (x"c4",x"0f",x"00",x"00"),
   374 => (x"0e",x"84",x"27",x"86"),
   375 => (x"27",x"1e",x"00",x"00"),
   376 => (x"00",x"00",x"01",x"17"),
   377 => (x"c0",x"86",x"c4",x"0f"),
   378 => (x"86",x"27",x"87",x"dc"),
   379 => (x"1e",x"00",x"00",x"0e"),
   380 => (x"00",x"01",x"17",x"27"),
   381 => (x"86",x"c4",x"0f",x"00"),
   382 => (x"00",x"0e",x"b5",x"27"),
   383 => (x"17",x"27",x"1e",x"00"),
   384 => (x"0f",x"00",x"00",x"01"),
   385 => (x"f8",x"27",x"86",x"c4"),
   386 => (x"bf",x"00",x"00",x"15"),
   387 => (x"10",x"43",x"27",x"1e"),
   388 => (x"27",x"1e",x"00",x"00"),
   389 => (x"00",x"00",x"01",x"17"),
   390 => (x"27",x"86",x"c8",x"0f"),
   391 => (x"00",x"00",x"04",x"f7"),
   392 => (x"3e",x"64",x"27",x"0f"),
   393 => (x"c1",x"58",x"00",x"00"),
   394 => (x"15",x"f8",x"27",x"4d"),
   395 => (x"49",x"bf",x"00",x"00"),
   396 => (x"06",x"a9",x"b7",x"c0"),
   397 => (x"27",x"87",x"f9",x"c6"),
   398 => (x"00",x"00",x"0e",x"42"),
   399 => (x"0e",x"01",x"27",x"0f"),
   400 => (x"76",x"0f",x"00",x"00"),
   401 => (x"c3",x"79",x"c2",x"49"),
   402 => (x"3e",x"f8",x"27",x"4c"),
   403 => (x"27",x"49",x"00",x"00"),
   404 => (x"00",x"00",x"0e",x"d6"),
   405 => (x"20",x"1e",x"72",x"48"),
   406 => (x"20",x"41",x"20",x"41"),
   407 => (x"20",x"41",x"20",x"41"),
   408 => (x"20",x"41",x"20",x"41"),
   409 => (x"10",x"51",x"10",x"41"),
   410 => (x"26",x"51",x"10",x"51"),
   411 => (x"49",x"a6",x"c8",x"4a"),
   412 => (x"f8",x"27",x"79",x"c1"),
   413 => (x"1e",x"00",x"00",x"3e"),
   414 => (x"00",x"3e",x"d8",x"27"),
   415 => (x"c3",x"27",x"1e",x"00"),
   416 => (x"0f",x"00",x"00",x"03"),
   417 => (x"4a",x"70",x"86",x"c8"),
   418 => (x"c0",x"05",x"9a",x"72"),
   419 => (x"4a",x"c1",x"87",x"c5"),
   420 => (x"c0",x"87",x"c2",x"c0"),
   421 => (x"16",x"7c",x"27",x"4a"),
   422 => (x"72",x"49",x"00",x"00"),
   423 => (x"74",x"49",x"6e",x"79"),
   424 => (x"c0",x"03",x"a9",x"b7"),
   425 => (x"4a",x"6e",x"87",x"ed"),
   426 => (x"48",x"72",x"92",x"c5"),
   427 => (x"a6",x"d0",x"88",x"74"),
   428 => (x"4a",x"a6",x"cc",x"58"),
   429 => (x"1e",x"74",x"1e",x"72"),
   430 => (x"27",x"1e",x"66",x"c8"),
   431 => (x"00",x"00",x"02",x"dc"),
   432 => (x"6e",x"86",x"cc",x"0f"),
   433 => (x"c4",x"80",x"c1",x"48"),
   434 => (x"49",x"6e",x"58",x"a6"),
   435 => (x"04",x"a9",x"b7",x"74"),
   436 => (x"cc",x"87",x"d3",x"ff"),
   437 => (x"66",x"c4",x"1e",x"66"),
   438 => (x"17",x"50",x"27",x"1e"),
   439 => (x"27",x"1e",x"00",x"00"),
   440 => (x"00",x"00",x"16",x"88"),
   441 => (x"02",x"f2",x"27",x"1e"),
   442 => (x"d0",x"0f",x"00",x"00"),
   443 => (x"16",x"70",x"27",x"86"),
   444 => (x"1e",x"bf",x"00",x"00"),
   445 => (x"00",x"0c",x"e2",x"27"),
   446 => (x"86",x"c4",x"0f",x"00"),
   447 => (x"c1",x"49",x"a6",x"c4"),
   448 => (x"81",x"27",x"51",x"c1"),
   449 => (x"97",x"00",x"00",x"16"),
   450 => (x"c0",x"c1",x"4a",x"bf"),
   451 => (x"92",x"c0",x"c0",x"c0"),
   452 => (x"92",x"b7",x"c0",x"c4"),
   453 => (x"b7",x"c1",x"c1",x"4a"),
   454 => (x"d8",x"c2",x"04",x"aa"),
   455 => (x"1e",x"c3",x"c1",x"87"),
   456 => (x"4a",x"66",x"c8",x"97"),
   457 => (x"c0",x"c0",x"c0",x"c1"),
   458 => (x"c0",x"c4",x"92",x"c0"),
   459 => (x"72",x"4a",x"92",x"b7"),
   460 => (x"03",x"7f",x"27",x"1e"),
   461 => (x"c8",x"0f",x"00",x"00"),
   462 => (x"c8",x"4a",x"70",x"86"),
   463 => (x"b7",x"72",x"49",x"66"),
   464 => (x"fd",x"c0",x"05",x"a9"),
   465 => (x"4a",x"a6",x"c8",x"87"),
   466 => (x"1e",x"c0",x"1e",x"72"),
   467 => (x"00",x"02",x"65",x"27"),
   468 => (x"86",x"c8",x"0f",x"00"),
   469 => (x"00",x"3e",x"f8",x"27"),
   470 => (x"b7",x"27",x"49",x"00"),
   471 => (x"48",x"00",x"00",x"0e"),
   472 => (x"41",x"20",x"1e",x"72"),
   473 => (x"41",x"20",x"41",x"20"),
   474 => (x"41",x"20",x"41",x"20"),
   475 => (x"41",x"20",x"41",x"20"),
   476 => (x"51",x"10",x"51",x"10"),
   477 => (x"4a",x"26",x"51",x"10"),
   478 => (x"78",x"27",x"4c",x"75"),
   479 => (x"49",x"00",x"00",x"16"),
   480 => (x"c4",x"97",x"79",x"75"),
   481 => (x"80",x"c1",x"48",x"66"),
   482 => (x"50",x"08",x"a6",x"c4"),
   483 => (x"4b",x"66",x"c4",x"97"),
   484 => (x"c0",x"c0",x"c0",x"c1"),
   485 => (x"c0",x"c4",x"93",x"c0"),
   486 => (x"27",x"4b",x"93",x"b7"),
   487 => (x"00",x"00",x"16",x"81"),
   488 => (x"c1",x"4a",x"bf",x"97"),
   489 => (x"c0",x"c0",x"c0",x"c0"),
   490 => (x"b7",x"c0",x"c4",x"92"),
   491 => (x"b7",x"72",x"4a",x"92"),
   492 => (x"e8",x"fd",x"06",x"ab"),
   493 => (x"74",x"94",x"6e",x"87"),
   494 => (x"d0",x"1e",x"72",x"49"),
   495 => (x"a0",x"27",x"4a",x"66"),
   496 => (x"0f",x"00",x"00",x"04"),
   497 => (x"48",x"70",x"4a",x"26"),
   498 => (x"74",x"58",x"a6",x"c4"),
   499 => (x"8a",x"66",x"cc",x"4a"),
   500 => (x"4c",x"72",x"92",x"c7"),
   501 => (x"4a",x"76",x"8c",x"6e"),
   502 => (x"7d",x"27",x"1e",x"72"),
   503 => (x"0f",x"00",x"00",x"0d"),
   504 => (x"85",x"c1",x"86",x"c4"),
   505 => (x"00",x"15",x"f8",x"27"),
   506 => (x"ad",x"b7",x"bf",x"00"),
   507 => (x"87",x"c7",x"f9",x"06"),
   508 => (x"00",x"04",x"f7",x"27"),
   509 => (x"68",x"27",x"0f",x"00"),
   510 => (x"58",x"00",x"00",x"3e"),
   511 => (x"00",x"10",x"70",x"27"),
   512 => (x"17",x"27",x"1e",x"00"),
   513 => (x"0f",x"00",x"00",x"01"),
   514 => (x"80",x"27",x"86",x"c4"),
   515 => (x"1e",x"00",x"00",x"10"),
   516 => (x"00",x"01",x"17",x"27"),
   517 => (x"86",x"c4",x"0f",x"00"),
   518 => (x"00",x"10",x"82",x"27"),
   519 => (x"17",x"27",x"1e",x"00"),
   520 => (x"0f",x"00",x"00",x"01"),
   521 => (x"b8",x"27",x"86",x"c4"),
   522 => (x"1e",x"00",x"00",x"10"),
   523 => (x"00",x"01",x"17",x"27"),
   524 => (x"86",x"c4",x"0f",x"00"),
   525 => (x"00",x"16",x"78",x"27"),
   526 => (x"27",x"1e",x"bf",x"00"),
   527 => (x"00",x"00",x"10",x"ba"),
   528 => (x"01",x"17",x"27",x"1e"),
   529 => (x"c8",x"0f",x"00",x"00"),
   530 => (x"27",x"1e",x"c5",x"86"),
   531 => (x"00",x"00",x"10",x"d3"),
   532 => (x"01",x"17",x"27",x"1e"),
   533 => (x"c8",x"0f",x"00",x"00"),
   534 => (x"16",x"7c",x"27",x"86"),
   535 => (x"1e",x"bf",x"00",x"00"),
   536 => (x"00",x"10",x"ec",x"27"),
   537 => (x"17",x"27",x"1e",x"00"),
   538 => (x"0f",x"00",x"00",x"01"),
   539 => (x"1e",x"c1",x"86",x"c8"),
   540 => (x"00",x"11",x"05",x"27"),
   541 => (x"17",x"27",x"1e",x"00"),
   542 => (x"0f",x"00",x"00",x"01"),
   543 => (x"80",x"27",x"86",x"c8"),
   544 => (x"97",x"00",x"00",x"16"),
   545 => (x"c0",x"c1",x"4a",x"bf"),
   546 => (x"92",x"c0",x"c0",x"c0"),
   547 => (x"92",x"b7",x"c0",x"c4"),
   548 => (x"27",x"1e",x"72",x"4a"),
   549 => (x"00",x"00",x"11",x"1e"),
   550 => (x"01",x"17",x"27",x"1e"),
   551 => (x"c8",x"0f",x"00",x"00"),
   552 => (x"1e",x"c1",x"c1",x"86"),
   553 => (x"00",x"11",x"37",x"27"),
   554 => (x"17",x"27",x"1e",x"00"),
   555 => (x"0f",x"00",x"00",x"01"),
   556 => (x"81",x"27",x"86",x"c8"),
   557 => (x"97",x"00",x"00",x"16"),
   558 => (x"c0",x"c1",x"4a",x"bf"),
   559 => (x"92",x"c0",x"c0",x"c0"),
   560 => (x"92",x"b7",x"c0",x"c4"),
   561 => (x"27",x"1e",x"72",x"4a"),
   562 => (x"00",x"00",x"11",x"50"),
   563 => (x"01",x"17",x"27",x"1e"),
   564 => (x"c8",x"0f",x"00",x"00"),
   565 => (x"1e",x"c2",x"c1",x"86"),
   566 => (x"00",x"11",x"69",x"27"),
   567 => (x"17",x"27",x"1e",x"00"),
   568 => (x"0f",x"00",x"00",x"01"),
   569 => (x"a8",x"27",x"86",x"c8"),
   570 => (x"bf",x"00",x"00",x"16"),
   571 => (x"11",x"82",x"27",x"1e"),
   572 => (x"27",x"1e",x"00",x"00"),
   573 => (x"00",x"00",x"01",x"17"),
   574 => (x"c7",x"86",x"c8",x"0f"),
   575 => (x"11",x"9b",x"27",x"1e"),
   576 => (x"27",x"1e",x"00",x"00"),
   577 => (x"00",x"00",x"01",x"17"),
   578 => (x"27",x"86",x"c8",x"0f"),
   579 => (x"00",x"00",x"1d",x"ac"),
   580 => (x"b4",x"27",x"1e",x"bf"),
   581 => (x"1e",x"00",x"00",x"11"),
   582 => (x"00",x"01",x"17",x"27"),
   583 => (x"86",x"c8",x"0f",x"00"),
   584 => (x"00",x"11",x"cd",x"27"),
   585 => (x"17",x"27",x"1e",x"00"),
   586 => (x"0f",x"00",x"00",x"01"),
   587 => (x"f7",x"27",x"86",x"c4"),
   588 => (x"1e",x"00",x"00",x"11"),
   589 => (x"00",x"01",x"17",x"27"),
   590 => (x"86",x"c4",x"0f",x"00"),
   591 => (x"00",x"16",x"70",x"27"),
   592 => (x"1e",x"bf",x"bf",x"00"),
   593 => (x"00",x"12",x"03",x"27"),
   594 => (x"17",x"27",x"1e",x"00"),
   595 => (x"0f",x"00",x"00",x"01"),
   596 => (x"1c",x"27",x"86",x"c8"),
   597 => (x"1e",x"00",x"00",x"12"),
   598 => (x"00",x"01",x"17",x"27"),
   599 => (x"86",x"c4",x"0f",x"00"),
   600 => (x"00",x"16",x"70",x"27"),
   601 => (x"c4",x"4a",x"bf",x"00"),
   602 => (x"27",x"1e",x"6a",x"82"),
   603 => (x"00",x"00",x"12",x"4d"),
   604 => (x"01",x"17",x"27",x"1e"),
   605 => (x"c8",x"0f",x"00",x"00"),
   606 => (x"27",x"1e",x"c0",x"86"),
   607 => (x"00",x"00",x"12",x"66"),
   608 => (x"01",x"17",x"27",x"1e"),
   609 => (x"c8",x"0f",x"00",x"00"),
   610 => (x"16",x"70",x"27",x"86"),
   611 => (x"4a",x"bf",x"00",x"00"),
   612 => (x"1e",x"6a",x"82",x"c8"),
   613 => (x"00",x"12",x"7f",x"27"),
   614 => (x"17",x"27",x"1e",x"00"),
   615 => (x"0f",x"00",x"00",x"01"),
   616 => (x"1e",x"c2",x"86",x"c8"),
   617 => (x"00",x"12",x"98",x"27"),
   618 => (x"17",x"27",x"1e",x"00"),
   619 => (x"0f",x"00",x"00",x"01"),
   620 => (x"70",x"27",x"86",x"c8"),
   621 => (x"bf",x"00",x"00",x"16"),
   622 => (x"6a",x"82",x"cc",x"4a"),
   623 => (x"12",x"b1",x"27",x"1e"),
   624 => (x"27",x"1e",x"00",x"00"),
   625 => (x"00",x"00",x"01",x"17"),
   626 => (x"d1",x"86",x"c8",x"0f"),
   627 => (x"12",x"ca",x"27",x"1e"),
   628 => (x"27",x"1e",x"00",x"00"),
   629 => (x"00",x"00",x"01",x"17"),
   630 => (x"27",x"86",x"c8",x"0f"),
   631 => (x"00",x"00",x"16",x"70"),
   632 => (x"82",x"d0",x"4a",x"bf"),
   633 => (x"e3",x"27",x"1e",x"72"),
   634 => (x"1e",x"00",x"00",x"12"),
   635 => (x"00",x"01",x"17",x"27"),
   636 => (x"86",x"c8",x"0f",x"00"),
   637 => (x"00",x"12",x"fc",x"27"),
   638 => (x"17",x"27",x"1e",x"00"),
   639 => (x"0f",x"00",x"00",x"01"),
   640 => (x"31",x"27",x"86",x"c4"),
   641 => (x"1e",x"00",x"00",x"13"),
   642 => (x"00",x"01",x"17",x"27"),
   643 => (x"86",x"c4",x"0f",x"00"),
   644 => (x"00",x"16",x"74",x"27"),
   645 => (x"1e",x"bf",x"bf",x"00"),
   646 => (x"00",x"13",x"42",x"27"),
   647 => (x"17",x"27",x"1e",x"00"),
   648 => (x"0f",x"00",x"00",x"01"),
   649 => (x"5b",x"27",x"86",x"c8"),
   650 => (x"1e",x"00",x"00",x"13"),
   651 => (x"00",x"01",x"17",x"27"),
   652 => (x"86",x"c4",x"0f",x"00"),
   653 => (x"00",x"16",x"74",x"27"),
   654 => (x"c4",x"4a",x"bf",x"00"),
   655 => (x"27",x"1e",x"6a",x"82"),
   656 => (x"00",x"00",x"13",x"9b"),
   657 => (x"01",x"17",x"27",x"1e"),
   658 => (x"c8",x"0f",x"00",x"00"),
   659 => (x"27",x"1e",x"c0",x"86"),
   660 => (x"00",x"00",x"13",x"b4"),
   661 => (x"01",x"17",x"27",x"1e"),
   662 => (x"c8",x"0f",x"00",x"00"),
   663 => (x"16",x"74",x"27",x"86"),
   664 => (x"4a",x"bf",x"00",x"00"),
   665 => (x"1e",x"6a",x"82",x"c8"),
   666 => (x"00",x"13",x"cd",x"27"),
   667 => (x"17",x"27",x"1e",x"00"),
   668 => (x"0f",x"00",x"00",x"01"),
   669 => (x"1e",x"c1",x"86",x"c8"),
   670 => (x"00",x"13",x"e6",x"27"),
   671 => (x"17",x"27",x"1e",x"00"),
   672 => (x"0f",x"00",x"00",x"01"),
   673 => (x"74",x"27",x"86",x"c8"),
   674 => (x"bf",x"00",x"00",x"16"),
   675 => (x"6a",x"82",x"cc",x"4a"),
   676 => (x"13",x"ff",x"27",x"1e"),
   677 => (x"27",x"1e",x"00",x"00"),
   678 => (x"00",x"00",x"01",x"17"),
   679 => (x"d2",x"86",x"c8",x"0f"),
   680 => (x"14",x"18",x"27",x"1e"),
   681 => (x"27",x"1e",x"00",x"00"),
   682 => (x"00",x"00",x"01",x"17"),
   683 => (x"27",x"86",x"c8",x"0f"),
   684 => (x"00",x"00",x"16",x"74"),
   685 => (x"82",x"d0",x"4a",x"bf"),
   686 => (x"31",x"27",x"1e",x"72"),
   687 => (x"1e",x"00",x"00",x"14"),
   688 => (x"00",x"01",x"17",x"27"),
   689 => (x"86",x"c8",x"0f",x"00"),
   690 => (x"00",x"14",x"4a",x"27"),
   691 => (x"17",x"27",x"1e",x"00"),
   692 => (x"0f",x"00",x"00",x"01"),
   693 => (x"1e",x"6e",x"86",x"c4"),
   694 => (x"00",x"14",x"7f",x"27"),
   695 => (x"17",x"27",x"1e",x"00"),
   696 => (x"0f",x"00",x"00",x"01"),
   697 => (x"1e",x"c5",x"86",x"c8"),
   698 => (x"00",x"14",x"98",x"27"),
   699 => (x"17",x"27",x"1e",x"00"),
   700 => (x"0f",x"00",x"00",x"01"),
   701 => (x"1e",x"74",x"86",x"c8"),
   702 => (x"00",x"14",x"b1",x"27"),
   703 => (x"17",x"27",x"1e",x"00"),
   704 => (x"0f",x"00",x"00",x"01"),
   705 => (x"1e",x"cd",x"86",x"c8"),
   706 => (x"00",x"14",x"ca",x"27"),
   707 => (x"17",x"27",x"1e",x"00"),
   708 => (x"0f",x"00",x"00",x"01"),
   709 => (x"66",x"cc",x"86",x"c8"),
   710 => (x"14",x"e3",x"27",x"1e"),
   711 => (x"27",x"1e",x"00",x"00"),
   712 => (x"00",x"00",x"01",x"17"),
   713 => (x"c7",x"86",x"c8",x"0f"),
   714 => (x"14",x"fc",x"27",x"1e"),
   715 => (x"27",x"1e",x"00",x"00"),
   716 => (x"00",x"00",x"01",x"17"),
   717 => (x"c8",x"86",x"c8",x"0f"),
   718 => (x"15",x"27",x"1e",x"66"),
   719 => (x"1e",x"00",x"00",x"15"),
   720 => (x"00",x"01",x"17",x"27"),
   721 => (x"86",x"c8",x"0f",x"00"),
   722 => (x"2e",x"27",x"1e",x"c1"),
   723 => (x"1e",x"00",x"00",x"15"),
   724 => (x"00",x"01",x"17",x"27"),
   725 => (x"86",x"c8",x"0f",x"00"),
   726 => (x"00",x"3e",x"d8",x"27"),
   727 => (x"47",x"27",x"1e",x"00"),
   728 => (x"1e",x"00",x"00",x"15"),
   729 => (x"00",x"01",x"17",x"27"),
   730 => (x"86",x"c8",x"0f",x"00"),
   731 => (x"00",x"15",x"60",x"27"),
   732 => (x"17",x"27",x"1e",x"00"),
   733 => (x"0f",x"00",x"00",x"01"),
   734 => (x"f8",x"27",x"86",x"c4"),
   735 => (x"1e",x"00",x"00",x"3e"),
   736 => (x"00",x"15",x"95",x"27"),
   737 => (x"17",x"27",x"1e",x"00"),
   738 => (x"0f",x"00",x"00",x"01"),
   739 => (x"ae",x"27",x"86",x"c8"),
   740 => (x"1e",x"00",x"00",x"15"),
   741 => (x"00",x"01",x"17",x"27"),
   742 => (x"86",x"c4",x"0f",x"00"),
   743 => (x"00",x"15",x"e3",x"27"),
   744 => (x"17",x"27",x"1e",x"00"),
   745 => (x"0f",x"00",x"00",x"01"),
   746 => (x"64",x"27",x"86",x"c4"),
   747 => (x"bf",x"00",x"00",x"3e"),
   748 => (x"3e",x"60",x"27",x"4a"),
   749 => (x"8a",x"bf",x"00",x"00"),
   750 => (x"00",x"3e",x"68",x"27"),
   751 => (x"79",x"72",x"49",x"00"),
   752 => (x"e5",x"27",x"1e",x"72"),
   753 => (x"1e",x"00",x"00",x"15"),
   754 => (x"00",x"01",x"17",x"27"),
   755 => (x"86",x"c8",x"0f",x"00"),
   756 => (x"00",x"3e",x"68",x"27"),
   757 => (x"c1",x"49",x"bf",x"00"),
   758 => (x"03",x"a9",x"b7",x"f8"),
   759 => (x"27",x"87",x"ea",x"c0"),
   760 => (x"00",x"00",x"0e",x"f5"),
   761 => (x"01",x"17",x"27",x"1e"),
   762 => (x"c4",x"0f",x"00",x"00"),
   763 => (x"0f",x"2b",x"27",x"86"),
   764 => (x"27",x"1e",x"00",x"00"),
   765 => (x"00",x"00",x"01",x"17"),
   766 => (x"27",x"86",x"c4",x"0f"),
   767 => (x"00",x"00",x"0f",x"4b"),
   768 => (x"01",x"17",x"27",x"1e"),
   769 => (x"c4",x"0f",x"00",x"00"),
   770 => (x"3e",x"68",x"27",x"86"),
   771 => (x"4a",x"bf",x"00",x"00"),
   772 => (x"e8",x"cf",x"4b",x"72"),
   773 => (x"72",x"49",x"73",x"93"),
   774 => (x"15",x"f8",x"27",x"1e"),
   775 => (x"4a",x"bf",x"00",x"00"),
   776 => (x"00",x"04",x"a0",x"27"),
   777 => (x"4a",x"26",x"0f",x"00"),
   778 => (x"70",x"27",x"48",x"70"),
   779 => (x"58",x"00",x"00",x"3e"),
   780 => (x"00",x"15",x"f8",x"27"),
   781 => (x"73",x"4b",x"bf",x"00"),
   782 => (x"94",x"e8",x"cf",x"4c"),
   783 => (x"1e",x"72",x"49",x"74"),
   784 => (x"a0",x"27",x"4a",x"72"),
   785 => (x"0f",x"00",x"00",x"04"),
   786 => (x"48",x"70",x"4a",x"26"),
   787 => (x"00",x"3e",x"74",x"27"),
   788 => (x"f9",x"c8",x"58",x"00"),
   789 => (x"72",x"49",x"73",x"93"),
   790 => (x"27",x"4a",x"72",x"1e"),
   791 => (x"00",x"00",x"04",x"a0"),
   792 => (x"70",x"4a",x"26",x"0f"),
   793 => (x"3e",x"78",x"27",x"48"),
   794 => (x"27",x"58",x"00",x"00"),
   795 => (x"00",x"00",x"0f",x"4d"),
   796 => (x"01",x"17",x"27",x"1e"),
   797 => (x"c4",x"0f",x"00",x"00"),
   798 => (x"3e",x"6c",x"27",x"86"),
   799 => (x"1e",x"bf",x"00",x"00"),
   800 => (x"00",x"0f",x"7a",x"27"),
   801 => (x"17",x"27",x"1e",x"00"),
   802 => (x"0f",x"00",x"00",x"01"),
   803 => (x"7f",x"27",x"86",x"c8"),
   804 => (x"1e",x"00",x"00",x"0f"),
   805 => (x"00",x"01",x"17",x"27"),
   806 => (x"86",x"c4",x"0f",x"00"),
   807 => (x"00",x"3e",x"70",x"27"),
   808 => (x"27",x"1e",x"bf",x"00"),
   809 => (x"00",x"00",x"0f",x"ac"),
   810 => (x"01",x"17",x"27",x"1e"),
   811 => (x"c8",x"0f",x"00",x"00"),
   812 => (x"3e",x"74",x"27",x"86"),
   813 => (x"1e",x"bf",x"00",x"00"),
   814 => (x"00",x"0f",x"b1",x"27"),
   815 => (x"17",x"27",x"1e",x"00"),
   816 => (x"0f",x"00",x"00",x"01"),
   817 => (x"cf",x"27",x"86",x"c8"),
   818 => (x"1e",x"00",x"00",x"0f"),
   819 => (x"00",x"01",x"17",x"27"),
   820 => (x"86",x"c4",x"0f",x"00"),
   821 => (x"86",x"d0",x"48",x"c0"),
   822 => (x"4c",x"26",x"4d",x"26"),
   823 => (x"4a",x"26",x"4b",x"26"),
   824 => (x"5e",x"0e",x"4f",x"26"),
   825 => (x"5d",x"5c",x"5b",x"5a"),
   826 => (x"bf",x"66",x"d4",x"0e"),
   827 => (x"27",x"4d",x"72",x"4a"),
   828 => (x"00",x"00",x"16",x"70"),
   829 => (x"1e",x"72",x"48",x"bf"),
   830 => (x"49",x"a2",x"f0",x"c0"),
   831 => (x"a9",x"72",x"42",x"20"),
   832 => (x"26",x"87",x"f9",x"05"),
   833 => (x"4c",x"66",x"d4",x"4a"),
   834 => (x"7c",x"c5",x"84",x"cc"),
   835 => (x"83",x"cc",x"4b",x"72"),
   836 => (x"66",x"d4",x"7b",x"6c"),
   837 => (x"1e",x"72",x"7a",x"bf"),
   838 => (x"00",x"0d",x"c9",x"27"),
   839 => (x"86",x"c4",x"0f",x"00"),
   840 => (x"9a",x"6a",x"82",x"c4"),
   841 => (x"87",x"f4",x"c0",x"05"),
   842 => (x"83",x"c8",x"4b",x"75"),
   843 => (x"82",x"cc",x"4a",x"75"),
   844 => (x"1e",x"73",x"7a",x"c6"),
   845 => (x"c8",x"4b",x"66",x"d8"),
   846 => (x"27",x"1e",x"6b",x"83"),
   847 => (x"00",x"00",x"02",x"65"),
   848 => (x"27",x"86",x"c8",x"0f"),
   849 => (x"00",x"00",x"16",x"70"),
   850 => (x"72",x"7d",x"bf",x"bf"),
   851 => (x"6a",x"1e",x"ca",x"1e"),
   852 => (x"02",x"dc",x"27",x"1e"),
   853 => (x"cc",x"0f",x"00",x"00"),
   854 => (x"87",x"d7",x"c0",x"86"),
   855 => (x"4a",x"bf",x"66",x"d4"),
   856 => (x"48",x"49",x"66",x"d4"),
   857 => (x"f0",x"c0",x"1e",x"72"),
   858 => (x"41",x"20",x"4a",x"a1"),
   859 => (x"f9",x"05",x"aa",x"71"),
   860 => (x"26",x"4a",x"26",x"87"),
   861 => (x"26",x"4c",x"26",x"4d"),
   862 => (x"26",x"4a",x"26",x"4b"),
   863 => (x"5a",x"5e",x"0e",x"4f"),
   864 => (x"0e",x"5d",x"5c",x"5b"),
   865 => (x"d8",x"4d",x"6e",x"1e"),
   866 => (x"4b",x"6c",x"4c",x"66"),
   867 => (x"80",x"27",x"83",x"ca"),
   868 => (x"97",x"00",x"00",x"16"),
   869 => (x"c0",x"c1",x"4a",x"bf"),
   870 => (x"92",x"c0",x"c0",x"c0"),
   871 => (x"92",x"b7",x"c0",x"c4"),
   872 => (x"b7",x"c1",x"c1",x"4a"),
   873 => (x"cf",x"c0",x"05",x"aa"),
   874 => (x"73",x"8b",x"c1",x"87"),
   875 => (x"16",x"78",x"27",x"48"),
   876 => (x"88",x"bf",x"00",x"00"),
   877 => (x"4d",x"c0",x"7c",x"70"),
   878 => (x"ff",x"05",x"9d",x"75"),
   879 => (x"26",x"26",x"87",x"d0"),
   880 => (x"26",x"4c",x"26",x"4d"),
   881 => (x"26",x"4a",x"26",x"4b"),
   882 => (x"1e",x"72",x"1e",x"4f"),
   883 => (x"00",x"16",x"70",x"27"),
   884 => (x"c0",x"02",x"bf",x"00"),
   885 => (x"66",x"c8",x"87",x"cb"),
   886 => (x"16",x"70",x"27",x"49"),
   887 => (x"bf",x"bf",x"00",x"00"),
   888 => (x"16",x"70",x"27",x"79"),
   889 => (x"4a",x"bf",x"00",x"00"),
   890 => (x"1e",x"72",x"82",x"cc"),
   891 => (x"00",x"16",x"78",x"27"),
   892 => (x"ca",x"1e",x"bf",x"00"),
   893 => (x"02",x"dc",x"27",x"1e"),
   894 => (x"cc",x"0f",x"00",x"00"),
   895 => (x"26",x"4a",x"26",x"86"),
   896 => (x"1e",x"72",x"1e",x"4f"),
   897 => (x"00",x"16",x"80",x"27"),
   898 => (x"4a",x"bf",x"97",x"00"),
   899 => (x"c0",x"c0",x"c0",x"c1"),
   900 => (x"c0",x"c4",x"92",x"c0"),
   901 => (x"c1",x"4a",x"92",x"b7"),
   902 => (x"02",x"aa",x"b7",x"c1"),
   903 => (x"c0",x"87",x"c5",x"c0"),
   904 => (x"87",x"c2",x"c0",x"4a"),
   905 => (x"7c",x"27",x"4a",x"c1"),
   906 => (x"bf",x"00",x"00",x"16"),
   907 => (x"27",x"b0",x"72",x"48"),
   908 => (x"00",x"00",x"16",x"80"),
   909 => (x"16",x"81",x"27",x"58"),
   910 => (x"c1",x"49",x"00",x"00"),
   911 => (x"4a",x"26",x"51",x"c2"),
   912 => (x"27",x"1e",x"4f",x"26"),
   913 => (x"00",x"00",x"16",x"80"),
   914 => (x"51",x"c1",x"c1",x"49"),
   915 => (x"00",x"16",x"7c",x"27"),
   916 => (x"79",x"c0",x"49",x"00"),
   917 => (x"00",x"00",x"4f",x"26"),
   918 => (x"67",x"6f",x"72",x"50"),
   919 => (x"20",x"6d",x"61",x"72"),
   920 => (x"70",x"6d",x"6f",x"63"),
   921 => (x"64",x"65",x"6c",x"69"),
   922 => (x"74",x"69",x"77",x"20"),
   923 => (x"72",x"27",x"20",x"68"),
   924 => (x"73",x"69",x"67",x"65"),
   925 => (x"27",x"72",x"65",x"74"),
   926 => (x"74",x"74",x"61",x"20"),
   927 => (x"75",x"62",x"69",x"72"),
   928 => (x"00",x"0a",x"65",x"74"),
   929 => (x"72",x"50",x"00",x"0a"),
   930 => (x"61",x"72",x"67",x"6f"),
   931 => (x"6f",x"63",x"20",x"6d"),
   932 => (x"6c",x"69",x"70",x"6d"),
   933 => (x"77",x"20",x"64",x"65"),
   934 => (x"6f",x"68",x"74",x"69"),
   935 => (x"27",x"20",x"74",x"75"),
   936 => (x"69",x"67",x"65",x"72"),
   937 => (x"72",x"65",x"74",x"73"),
   938 => (x"74",x"61",x"20",x"27"),
   939 => (x"62",x"69",x"72",x"74"),
   940 => (x"0a",x"65",x"74",x"75"),
   941 => (x"44",x"00",x"0a",x"00"),
   942 => (x"53",x"59",x"52",x"48"),
   943 => (x"45",x"4e",x"4f",x"54"),
   944 => (x"4f",x"52",x"50",x"20"),
   945 => (x"4d",x"41",x"52",x"47"),
   946 => (x"27",x"33",x"20",x"2c"),
   947 => (x"53",x"20",x"44",x"52"),
   948 => (x"4e",x"49",x"52",x"54"),
   949 => (x"48",x"44",x"00",x"47"),
   950 => (x"54",x"53",x"59",x"52"),
   951 => (x"20",x"45",x"4e",x"4f"),
   952 => (x"47",x"4f",x"52",x"50"),
   953 => (x"2c",x"4d",x"41",x"52"),
   954 => (x"4e",x"27",x"32",x"20"),
   955 => (x"54",x"53",x"20",x"44"),
   956 => (x"47",x"4e",x"49",x"52"),
   957 => (x"61",x"65",x"4d",x"00"),
   958 => (x"65",x"72",x"75",x"73"),
   959 => (x"69",x"74",x"20",x"64"),
   960 => (x"74",x"20",x"65",x"6d"),
   961 => (x"73",x"20",x"6f",x"6f"),
   962 => (x"6c",x"6c",x"61",x"6d"),
   963 => (x"20",x"6f",x"74",x"20"),
   964 => (x"61",x"74",x"62",x"6f"),
   965 => (x"6d",x"20",x"6e",x"69"),
   966 => (x"69",x"6e",x"61",x"65"),
   967 => (x"75",x"66",x"67",x"6e"),
   968 => (x"65",x"72",x"20",x"6c"),
   969 => (x"74",x"6c",x"75",x"73"),
   970 => (x"50",x"00",x"0a",x"73"),
   971 => (x"73",x"61",x"65",x"6c"),
   972 => (x"6e",x"69",x"20",x"65"),
   973 => (x"61",x"65",x"72",x"63"),
   974 => (x"6e",x"20",x"65",x"73"),
   975 => (x"65",x"62",x"6d",x"75"),
   976 => (x"66",x"6f",x"20",x"72"),
   977 => (x"6e",x"75",x"72",x"20"),
   978 => (x"0a",x"00",x"0a",x"73"),
   979 => (x"63",x"69",x"4d",x"00"),
   980 => (x"65",x"73",x"6f",x"72"),
   981 => (x"64",x"6e",x"6f",x"63"),
   982 => (x"6f",x"66",x"20",x"73"),
   983 => (x"6e",x"6f",x"20",x"72"),
   984 => (x"75",x"72",x"20",x"65"),
   985 => (x"68",x"74",x"20",x"6e"),
   986 => (x"67",x"75",x"6f",x"72"),
   987 => (x"68",x"44",x"20",x"68"),
   988 => (x"74",x"73",x"79",x"72"),
   989 => (x"3a",x"65",x"6e",x"6f"),
   990 => (x"64",x"25",x"00",x"20"),
   991 => (x"44",x"00",x"0a",x"20"),
   992 => (x"73",x"79",x"72",x"68"),
   993 => (x"65",x"6e",x"6f",x"74"),
   994 => (x"65",x"70",x"20",x"73"),
   995 => (x"65",x"53",x"20",x"72"),
   996 => (x"64",x"6e",x"6f",x"63"),
   997 => (x"20",x"20",x"20",x"3a"),
   998 => (x"20",x"20",x"20",x"20"),
   999 => (x"20",x"20",x"20",x"20"),
  1000 => (x"20",x"20",x"20",x"20"),
  1001 => (x"20",x"20",x"20",x"20"),
  1002 => (x"00",x"20",x"20",x"20"),
  1003 => (x"0a",x"20",x"64",x"25"),
  1004 => (x"58",x"41",x"56",x"00"),
  1005 => (x"50",x"49",x"4d",x"20"),
  1006 => (x"61",x"72",x"20",x"53"),
  1007 => (x"67",x"6e",x"69",x"74"),
  1008 => (x"31",x"20",x"2a",x"20"),
  1009 => (x"20",x"30",x"30",x"30"),
  1010 => (x"64",x"25",x"20",x"3d"),
  1011 => (x"0a",x"00",x"0a",x"20"),
  1012 => (x"52",x"48",x"44",x"00"),
  1013 => (x"4f",x"54",x"53",x"59"),
  1014 => (x"50",x"20",x"45",x"4e"),
  1015 => (x"52",x"47",x"4f",x"52"),
  1016 => (x"20",x"2c",x"4d",x"41"),
  1017 => (x"45",x"4d",x"4f",x"53"),
  1018 => (x"52",x"54",x"53",x"20"),
  1019 => (x"00",x"47",x"4e",x"49"),
  1020 => (x"59",x"52",x"48",x"44"),
  1021 => (x"4e",x"4f",x"54",x"53"),
  1022 => (x"52",x"50",x"20",x"45"),
  1023 => (x"41",x"52",x"47",x"4f"),
  1024 => (x"31",x"20",x"2c",x"4d"),
  1025 => (x"20",x"54",x"53",x"27"),
  1026 => (x"49",x"52",x"54",x"53"),
  1027 => (x"0a",x"00",x"47",x"4e"),
  1028 => (x"72",x"68",x"44",x"00"),
  1029 => (x"6f",x"74",x"73",x"79"),
  1030 => (x"42",x"20",x"65",x"6e"),
  1031 => (x"68",x"63",x"6e",x"65"),
  1032 => (x"6b",x"72",x"61",x"6d"),
  1033 => (x"65",x"56",x"20",x"2c"),
  1034 => (x"6f",x"69",x"73",x"72"),
  1035 => (x"2e",x"32",x"20",x"6e"),
  1036 => (x"4c",x"28",x"20",x"31"),
  1037 => (x"75",x"67",x"6e",x"61"),
  1038 => (x"3a",x"65",x"67",x"61"),
  1039 => (x"0a",x"29",x"43",x"20"),
  1040 => (x"45",x"00",x"0a",x"00"),
  1041 => (x"75",x"63",x"65",x"78"),
  1042 => (x"6e",x"6f",x"69",x"74"),
  1043 => (x"61",x"74",x"73",x"20"),
  1044 => (x"2c",x"73",x"74",x"72"),
  1045 => (x"20",x"64",x"25",x"20"),
  1046 => (x"73",x"6e",x"75",x"72"),
  1047 => (x"72",x"68",x"74",x"20"),
  1048 => (x"68",x"67",x"75",x"6f"),
  1049 => (x"72",x"68",x"44",x"20"),
  1050 => (x"6f",x"74",x"73",x"79"),
  1051 => (x"00",x"0a",x"65",x"6e"),
  1052 => (x"63",x"65",x"78",x"45"),
  1053 => (x"6f",x"69",x"74",x"75"),
  1054 => (x"6e",x"65",x"20",x"6e"),
  1055 => (x"00",x"0a",x"73",x"64"),
  1056 => (x"69",x"46",x"00",x"0a"),
  1057 => (x"20",x"6c",x"61",x"6e"),
  1058 => (x"75",x"6c",x"61",x"76"),
  1059 => (x"6f",x"20",x"73",x"65"),
  1060 => (x"68",x"74",x"20",x"66"),
  1061 => (x"61",x"76",x"20",x"65"),
  1062 => (x"62",x"61",x"69",x"72"),
  1063 => (x"20",x"73",x"65",x"6c"),
  1064 => (x"64",x"65",x"73",x"75"),
  1065 => (x"20",x"6e",x"69",x"20"),
  1066 => (x"20",x"65",x"68",x"74"),
  1067 => (x"63",x"6e",x"65",x"62"),
  1068 => (x"72",x"61",x"6d",x"68"),
  1069 => (x"00",x"0a",x"3a",x"6b"),
  1070 => (x"6e",x"49",x"00",x"0a"),
  1071 => (x"6c",x"47",x"5f",x"74"),
  1072 => (x"20",x"3a",x"62",x"6f"),
  1073 => (x"20",x"20",x"20",x"20"),
  1074 => (x"20",x"20",x"20",x"20"),
  1075 => (x"25",x"20",x"20",x"20"),
  1076 => (x"20",x"00",x"0a",x"64"),
  1077 => (x"20",x"20",x"20",x"20"),
  1078 => (x"73",x"20",x"20",x"20"),
  1079 => (x"6c",x"75",x"6f",x"68"),
  1080 => (x"65",x"62",x"20",x"64"),
  1081 => (x"20",x"20",x"20",x"3a"),
  1082 => (x"00",x"0a",x"64",x"25"),
  1083 => (x"6c",x"6f",x"6f",x"42"),
  1084 => (x"6f",x"6c",x"47",x"5f"),
  1085 => (x"20",x"20",x"3a",x"62"),
  1086 => (x"20",x"20",x"20",x"20"),
  1087 => (x"20",x"20",x"20",x"20"),
  1088 => (x"0a",x"64",x"25",x"20"),
  1089 => (x"20",x"20",x"20",x"00"),
  1090 => (x"20",x"20",x"20",x"20"),
  1091 => (x"6f",x"68",x"73",x"20"),
  1092 => (x"20",x"64",x"6c",x"75"),
  1093 => (x"20",x"3a",x"65",x"62"),
  1094 => (x"64",x"25",x"20",x"20"),
  1095 => (x"68",x"43",x"00",x"0a"),
  1096 => (x"47",x"5f",x"31",x"5f"),
  1097 => (x"3a",x"62",x"6f",x"6c"),
  1098 => (x"20",x"20",x"20",x"20"),
  1099 => (x"20",x"20",x"20",x"20"),
  1100 => (x"25",x"20",x"20",x"20"),
  1101 => (x"20",x"00",x"0a",x"63"),
  1102 => (x"20",x"20",x"20",x"20"),
  1103 => (x"73",x"20",x"20",x"20"),
  1104 => (x"6c",x"75",x"6f",x"68"),
  1105 => (x"65",x"62",x"20",x"64"),
  1106 => (x"20",x"20",x"20",x"3a"),
  1107 => (x"00",x"0a",x"63",x"25"),
  1108 => (x"32",x"5f",x"68",x"43"),
  1109 => (x"6f",x"6c",x"47",x"5f"),
  1110 => (x"20",x"20",x"3a",x"62"),
  1111 => (x"20",x"20",x"20",x"20"),
  1112 => (x"20",x"20",x"20",x"20"),
  1113 => (x"0a",x"63",x"25",x"20"),
  1114 => (x"20",x"20",x"20",x"00"),
  1115 => (x"20",x"20",x"20",x"20"),
  1116 => (x"6f",x"68",x"73",x"20"),
  1117 => (x"20",x"64",x"6c",x"75"),
  1118 => (x"20",x"3a",x"65",x"62"),
  1119 => (x"63",x"25",x"20",x"20"),
  1120 => (x"72",x"41",x"00",x"0a"),
  1121 => (x"5f",x"31",x"5f",x"72"),
  1122 => (x"62",x"6f",x"6c",x"47"),
  1123 => (x"3a",x"5d",x"38",x"5b"),
  1124 => (x"20",x"20",x"20",x"20"),
  1125 => (x"25",x"20",x"20",x"20"),
  1126 => (x"20",x"00",x"0a",x"64"),
  1127 => (x"20",x"20",x"20",x"20"),
  1128 => (x"73",x"20",x"20",x"20"),
  1129 => (x"6c",x"75",x"6f",x"68"),
  1130 => (x"65",x"62",x"20",x"64"),
  1131 => (x"20",x"20",x"20",x"3a"),
  1132 => (x"00",x"0a",x"64",x"25"),
  1133 => (x"5f",x"72",x"72",x"41"),
  1134 => (x"6c",x"47",x"5f",x"32"),
  1135 => (x"38",x"5b",x"62",x"6f"),
  1136 => (x"5d",x"37",x"5b",x"5d"),
  1137 => (x"20",x"20",x"20",x"3a"),
  1138 => (x"0a",x"64",x"25",x"20"),
  1139 => (x"20",x"20",x"20",x"00"),
  1140 => (x"20",x"20",x"20",x"20"),
  1141 => (x"6f",x"68",x"73",x"20"),
  1142 => (x"20",x"64",x"6c",x"75"),
  1143 => (x"20",x"3a",x"65",x"62"),
  1144 => (x"75",x"4e",x"20",x"20"),
  1145 => (x"72",x"65",x"62",x"6d"),
  1146 => (x"5f",x"66",x"4f",x"5f"),
  1147 => (x"73",x"6e",x"75",x"52"),
  1148 => (x"31",x"20",x"2b",x"20"),
  1149 => (x"50",x"00",x"0a",x"30"),
  1150 => (x"47",x"5f",x"72",x"74"),
  1151 => (x"2d",x"62",x"6f",x"6c"),
  1152 => (x"20",x"00",x"0a",x"3e"),
  1153 => (x"72",x"74",x"50",x"20"),
  1154 => (x"6d",x"6f",x"43",x"5f"),
  1155 => (x"20",x"20",x"3a",x"70"),
  1156 => (x"20",x"20",x"20",x"20"),
  1157 => (x"20",x"20",x"20",x"20"),
  1158 => (x"00",x"0a",x"64",x"25"),
  1159 => (x"20",x"20",x"20",x"20"),
  1160 => (x"20",x"20",x"20",x"20"),
  1161 => (x"75",x"6f",x"68",x"73"),
  1162 => (x"62",x"20",x"64",x"6c"),
  1163 => (x"20",x"20",x"3a",x"65"),
  1164 => (x"6d",x"69",x"28",x"20"),
  1165 => (x"6d",x"65",x"6c",x"70"),
  1166 => (x"61",x"74",x"6e",x"65"),
  1167 => (x"6e",x"6f",x"69",x"74"),
  1168 => (x"70",x"65",x"64",x"2d"),
  1169 => (x"65",x"64",x"6e",x"65"),
  1170 => (x"0a",x"29",x"74",x"6e"),
  1171 => (x"44",x"20",x"20",x"00"),
  1172 => (x"72",x"63",x"73",x"69"),
  1173 => (x"20",x"20",x"20",x"3a"),
  1174 => (x"20",x"20",x"20",x"20"),
  1175 => (x"20",x"20",x"20",x"20"),
  1176 => (x"64",x"25",x"20",x"20"),
  1177 => (x"20",x"20",x"00",x"0a"),
  1178 => (x"20",x"20",x"20",x"20"),
  1179 => (x"68",x"73",x"20",x"20"),
  1180 => (x"64",x"6c",x"75",x"6f"),
  1181 => (x"3a",x"65",x"62",x"20"),
  1182 => (x"25",x"20",x"20",x"20"),
  1183 => (x"20",x"00",x"0a",x"64"),
  1184 => (x"75",x"6e",x"45",x"20"),
  1185 => (x"6f",x"43",x"5f",x"6d"),
  1186 => (x"20",x"3a",x"70",x"6d"),
  1187 => (x"20",x"20",x"20",x"20"),
  1188 => (x"20",x"20",x"20",x"20"),
  1189 => (x"00",x"0a",x"64",x"25"),
  1190 => (x"20",x"20",x"20",x"20"),
  1191 => (x"20",x"20",x"20",x"20"),
  1192 => (x"75",x"6f",x"68",x"73"),
  1193 => (x"62",x"20",x"64",x"6c"),
  1194 => (x"20",x"20",x"3a",x"65"),
  1195 => (x"0a",x"64",x"25",x"20"),
  1196 => (x"49",x"20",x"20",x"00"),
  1197 => (x"43",x"5f",x"74",x"6e"),
  1198 => (x"3a",x"70",x"6d",x"6f"),
  1199 => (x"20",x"20",x"20",x"20"),
  1200 => (x"20",x"20",x"20",x"20"),
  1201 => (x"64",x"25",x"20",x"20"),
  1202 => (x"20",x"20",x"00",x"0a"),
  1203 => (x"20",x"20",x"20",x"20"),
  1204 => (x"68",x"73",x"20",x"20"),
  1205 => (x"64",x"6c",x"75",x"6f"),
  1206 => (x"3a",x"65",x"62",x"20"),
  1207 => (x"25",x"20",x"20",x"20"),
  1208 => (x"20",x"00",x"0a",x"64"),
  1209 => (x"72",x"74",x"53",x"20"),
  1210 => (x"6d",x"6f",x"43",x"5f"),
  1211 => (x"20",x"20",x"3a",x"70"),
  1212 => (x"20",x"20",x"20",x"20"),
  1213 => (x"20",x"20",x"20",x"20"),
  1214 => (x"00",x"0a",x"73",x"25"),
  1215 => (x"20",x"20",x"20",x"20"),
  1216 => (x"20",x"20",x"20",x"20"),
  1217 => (x"75",x"6f",x"68",x"73"),
  1218 => (x"62",x"20",x"64",x"6c"),
  1219 => (x"20",x"20",x"3a",x"65"),
  1220 => (x"52",x"48",x"44",x"20"),
  1221 => (x"4f",x"54",x"53",x"59"),
  1222 => (x"50",x"20",x"45",x"4e"),
  1223 => (x"52",x"47",x"4f",x"52"),
  1224 => (x"20",x"2c",x"4d",x"41"),
  1225 => (x"45",x"4d",x"4f",x"53"),
  1226 => (x"52",x"54",x"53",x"20"),
  1227 => (x"0a",x"47",x"4e",x"49"),
  1228 => (x"78",x"65",x"4e",x"00"),
  1229 => (x"74",x"50",x"5f",x"74"),
  1230 => (x"6c",x"47",x"5f",x"72"),
  1231 => (x"3e",x"2d",x"62",x"6f"),
  1232 => (x"20",x"20",x"00",x"0a"),
  1233 => (x"5f",x"72",x"74",x"50"),
  1234 => (x"70",x"6d",x"6f",x"43"),
  1235 => (x"20",x"20",x"20",x"3a"),
  1236 => (x"20",x"20",x"20",x"20"),
  1237 => (x"25",x"20",x"20",x"20"),
  1238 => (x"20",x"00",x"0a",x"64"),
  1239 => (x"20",x"20",x"20",x"20"),
  1240 => (x"73",x"20",x"20",x"20"),
  1241 => (x"6c",x"75",x"6f",x"68"),
  1242 => (x"65",x"62",x"20",x"64"),
  1243 => (x"20",x"20",x"20",x"3a"),
  1244 => (x"70",x"6d",x"69",x"28"),
  1245 => (x"65",x"6d",x"65",x"6c"),
  1246 => (x"74",x"61",x"74",x"6e"),
  1247 => (x"2d",x"6e",x"6f",x"69"),
  1248 => (x"65",x"70",x"65",x"64"),
  1249 => (x"6e",x"65",x"64",x"6e"),
  1250 => (x"20",x"2c",x"29",x"74"),
  1251 => (x"65",x"6d",x"61",x"73"),
  1252 => (x"20",x"73",x"61",x"20"),
  1253 => (x"76",x"6f",x"62",x"61"),
  1254 => (x"20",x"00",x"0a",x"65"),
  1255 => (x"73",x"69",x"44",x"20"),
  1256 => (x"20",x"3a",x"72",x"63"),
  1257 => (x"20",x"20",x"20",x"20"),
  1258 => (x"20",x"20",x"20",x"20"),
  1259 => (x"20",x"20",x"20",x"20"),
  1260 => (x"00",x"0a",x"64",x"25"),
  1261 => (x"20",x"20",x"20",x"20"),
  1262 => (x"20",x"20",x"20",x"20"),
  1263 => (x"75",x"6f",x"68",x"73"),
  1264 => (x"62",x"20",x"64",x"6c"),
  1265 => (x"20",x"20",x"3a",x"65"),
  1266 => (x"0a",x"64",x"25",x"20"),
  1267 => (x"45",x"20",x"20",x"00"),
  1268 => (x"5f",x"6d",x"75",x"6e"),
  1269 => (x"70",x"6d",x"6f",x"43"),
  1270 => (x"20",x"20",x"20",x"3a"),
  1271 => (x"20",x"20",x"20",x"20"),
  1272 => (x"64",x"25",x"20",x"20"),
  1273 => (x"20",x"20",x"00",x"0a"),
  1274 => (x"20",x"20",x"20",x"20"),
  1275 => (x"68",x"73",x"20",x"20"),
  1276 => (x"64",x"6c",x"75",x"6f"),
  1277 => (x"3a",x"65",x"62",x"20"),
  1278 => (x"25",x"20",x"20",x"20"),
  1279 => (x"20",x"00",x"0a",x"64"),
  1280 => (x"74",x"6e",x"49",x"20"),
  1281 => (x"6d",x"6f",x"43",x"5f"),
  1282 => (x"20",x"20",x"3a",x"70"),
  1283 => (x"20",x"20",x"20",x"20"),
  1284 => (x"20",x"20",x"20",x"20"),
  1285 => (x"00",x"0a",x"64",x"25"),
  1286 => (x"20",x"20",x"20",x"20"),
  1287 => (x"20",x"20",x"20",x"20"),
  1288 => (x"75",x"6f",x"68",x"73"),
  1289 => (x"62",x"20",x"64",x"6c"),
  1290 => (x"20",x"20",x"3a",x"65"),
  1291 => (x"0a",x"64",x"25",x"20"),
  1292 => (x"53",x"20",x"20",x"00"),
  1293 => (x"43",x"5f",x"72",x"74"),
  1294 => (x"3a",x"70",x"6d",x"6f"),
  1295 => (x"20",x"20",x"20",x"20"),
  1296 => (x"20",x"20",x"20",x"20"),
  1297 => (x"73",x"25",x"20",x"20"),
  1298 => (x"20",x"20",x"00",x"0a"),
  1299 => (x"20",x"20",x"20",x"20"),
  1300 => (x"68",x"73",x"20",x"20"),
  1301 => (x"64",x"6c",x"75",x"6f"),
  1302 => (x"3a",x"65",x"62",x"20"),
  1303 => (x"44",x"20",x"20",x"20"),
  1304 => (x"53",x"59",x"52",x"48"),
  1305 => (x"45",x"4e",x"4f",x"54"),
  1306 => (x"4f",x"52",x"50",x"20"),
  1307 => (x"4d",x"41",x"52",x"47"),
  1308 => (x"4f",x"53",x"20",x"2c"),
  1309 => (x"53",x"20",x"45",x"4d"),
  1310 => (x"4e",x"49",x"52",x"54"),
  1311 => (x"49",x"00",x"0a",x"47"),
  1312 => (x"31",x"5f",x"74",x"6e"),
  1313 => (x"63",x"6f",x"4c",x"5f"),
  1314 => (x"20",x"20",x"20",x"3a"),
  1315 => (x"20",x"20",x"20",x"20"),
  1316 => (x"20",x"20",x"20",x"20"),
  1317 => (x"00",x"0a",x"64",x"25"),
  1318 => (x"20",x"20",x"20",x"20"),
  1319 => (x"20",x"20",x"20",x"20"),
  1320 => (x"75",x"6f",x"68",x"73"),
  1321 => (x"62",x"20",x"64",x"6c"),
  1322 => (x"20",x"20",x"3a",x"65"),
  1323 => (x"0a",x"64",x"25",x"20"),
  1324 => (x"74",x"6e",x"49",x"00"),
  1325 => (x"4c",x"5f",x"32",x"5f"),
  1326 => (x"20",x"3a",x"63",x"6f"),
  1327 => (x"20",x"20",x"20",x"20"),
  1328 => (x"20",x"20",x"20",x"20"),
  1329 => (x"64",x"25",x"20",x"20"),
  1330 => (x"20",x"20",x"00",x"0a"),
  1331 => (x"20",x"20",x"20",x"20"),
  1332 => (x"68",x"73",x"20",x"20"),
  1333 => (x"64",x"6c",x"75",x"6f"),
  1334 => (x"3a",x"65",x"62",x"20"),
  1335 => (x"25",x"20",x"20",x"20"),
  1336 => (x"49",x"00",x"0a",x"64"),
  1337 => (x"33",x"5f",x"74",x"6e"),
  1338 => (x"63",x"6f",x"4c",x"5f"),
  1339 => (x"20",x"20",x"20",x"3a"),
  1340 => (x"20",x"20",x"20",x"20"),
  1341 => (x"20",x"20",x"20",x"20"),
  1342 => (x"00",x"0a",x"64",x"25"),
  1343 => (x"20",x"20",x"20",x"20"),
  1344 => (x"20",x"20",x"20",x"20"),
  1345 => (x"75",x"6f",x"68",x"73"),
  1346 => (x"62",x"20",x"64",x"6c"),
  1347 => (x"20",x"20",x"3a",x"65"),
  1348 => (x"0a",x"64",x"25",x"20"),
  1349 => (x"75",x"6e",x"45",x"00"),
  1350 => (x"6f",x"4c",x"5f",x"6d"),
  1351 => (x"20",x"20",x"3a",x"63"),
  1352 => (x"20",x"20",x"20",x"20"),
  1353 => (x"20",x"20",x"20",x"20"),
  1354 => (x"64",x"25",x"20",x"20"),
  1355 => (x"20",x"20",x"00",x"0a"),
  1356 => (x"20",x"20",x"20",x"20"),
  1357 => (x"68",x"73",x"20",x"20"),
  1358 => (x"64",x"6c",x"75",x"6f"),
  1359 => (x"3a",x"65",x"62",x"20"),
  1360 => (x"25",x"20",x"20",x"20"),
  1361 => (x"53",x"00",x"0a",x"64"),
  1362 => (x"31",x"5f",x"72",x"74"),
  1363 => (x"63",x"6f",x"4c",x"5f"),
  1364 => (x"20",x"20",x"20",x"3a"),
  1365 => (x"20",x"20",x"20",x"20"),
  1366 => (x"20",x"20",x"20",x"20"),
  1367 => (x"00",x"0a",x"73",x"25"),
  1368 => (x"20",x"20",x"20",x"20"),
  1369 => (x"20",x"20",x"20",x"20"),
  1370 => (x"75",x"6f",x"68",x"73"),
  1371 => (x"62",x"20",x"64",x"6c"),
  1372 => (x"20",x"20",x"3a",x"65"),
  1373 => (x"52",x"48",x"44",x"20"),
  1374 => (x"4f",x"54",x"53",x"59"),
  1375 => (x"50",x"20",x"45",x"4e"),
  1376 => (x"52",x"47",x"4f",x"52"),
  1377 => (x"20",x"2c",x"4d",x"41"),
  1378 => (x"54",x"53",x"27",x"31"),
  1379 => (x"52",x"54",x"53",x"20"),
  1380 => (x"0a",x"47",x"4e",x"49"),
  1381 => (x"72",x"74",x"53",x"00"),
  1382 => (x"4c",x"5f",x"32",x"5f"),
  1383 => (x"20",x"3a",x"63",x"6f"),
  1384 => (x"20",x"20",x"20",x"20"),
  1385 => (x"20",x"20",x"20",x"20"),
  1386 => (x"73",x"25",x"20",x"20"),
  1387 => (x"20",x"20",x"00",x"0a"),
  1388 => (x"20",x"20",x"20",x"20"),
  1389 => (x"68",x"73",x"20",x"20"),
  1390 => (x"64",x"6c",x"75",x"6f"),
  1391 => (x"3a",x"65",x"62",x"20"),
  1392 => (x"44",x"20",x"20",x"20"),
  1393 => (x"53",x"59",x"52",x"48"),
  1394 => (x"45",x"4e",x"4f",x"54"),
  1395 => (x"4f",x"52",x"50",x"20"),
  1396 => (x"4d",x"41",x"52",x"47"),
  1397 => (x"27",x"32",x"20",x"2c"),
  1398 => (x"53",x"20",x"44",x"4e"),
  1399 => (x"4e",x"49",x"52",x"54"),
  1400 => (x"0a",x"00",x"0a",x"47"),
  1401 => (x"65",x"73",x"55",x"00"),
  1402 => (x"69",x"74",x"20",x"72"),
  1403 => (x"20",x"3a",x"65",x"6d"),
  1404 => (x"00",x"0a",x"64",x"25"),
  1405 => (x"00",x"00",x"00",x"00"),
  1406 => (x"00",x"00",x"61",x"a8"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
