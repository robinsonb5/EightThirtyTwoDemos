
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"3b",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"38"),
    10 => (x"20",x"00",x"27",x"4f"),
    11 => (x"27",x"4e",x"00",x"00"),
    12 => (x"00",x"00",x"13",x"64"),
    13 => (x"87",x"fd",x"00",x"0f"),
    14 => (x"4f",x"87",x"fd",x"00"),
    15 => (x"ff",x"86",x"fc",x"1e"),
    16 => (x"48",x"69",x"49",x"c0"),
    17 => (x"c4",x"98",x"c0",x"c4"),
    18 => (x"02",x"6e",x"58",x"a6"),
    19 => (x"66",x"c8",x"87",x"f4"),
    20 => (x"8e",x"fc",x"48",x"79"),
    21 => (x"5e",x"0e",x"4f",x"26"),
    22 => (x"0e",x"5d",x"5c",x"5b"),
    23 => (x"c0",x"4b",x"66",x"d0"),
    24 => (x"c3",x"49",x"13",x"4c"),
    25 => (x"99",x"71",x"99",x"ff"),
    26 => (x"71",x"87",x"db",x"02"),
    27 => (x"4a",x"c0",x"ff",x"4d"),
    28 => (x"c0",x"c4",x"49",x"6a"),
    29 => (x"87",x"f8",x"02",x"99"),
    30 => (x"84",x"c1",x"7a",x"75"),
    31 => (x"ff",x"c3",x"49",x"13"),
    32 => (x"05",x"99",x"71",x"99"),
    33 => (x"48",x"74",x"87",x"e5"),
    34 => (x"4c",x"26",x"4d",x"26"),
    35 => (x"4f",x"26",x"4b",x"26"),
    36 => (x"5c",x"5b",x"5e",x"0e"),
    37 => (x"86",x"f0",x"0e",x"5d"),
    38 => (x"a6",x"c4",x"4b",x"c0"),
    39 => (x"c0",x"78",x"c0",x"48"),
    40 => (x"c0",x"4c",x"a6",x"e4"),
    41 => (x"48",x"49",x"66",x"e0"),
    42 => (x"e4",x"c0",x"80",x"c1"),
    43 => (x"4a",x"11",x"58",x"a6"),
    44 => (x"ba",x"82",x"c0",x"fe"),
    45 => (x"c4",x"02",x"9a",x"72"),
    46 => (x"66",x"c4",x"87",x"d2"),
    47 => (x"87",x"e1",x"c3",x"02"),
    48 => (x"c0",x"48",x"a6",x"c4"),
    49 => (x"c0",x"49",x"72",x"78"),
    50 => (x"c2",x"02",x"aa",x"f0"),
    51 => (x"e3",x"c1",x"87",x"f1"),
    52 => (x"f2",x"c2",x"02",x"a9"),
    53 => (x"a9",x"e4",x"c1",x"87"),
    54 => (x"87",x"e1",x"c0",x"02"),
    55 => (x"02",x"a9",x"ec",x"c1"),
    56 => (x"c1",x"87",x"dc",x"c2"),
    57 => (x"d4",x"02",x"a9",x"f0"),
    58 => (x"a9",x"f3",x"c1",x"87"),
    59 => (x"87",x"fa",x"c1",x"02"),
    60 => (x"02",x"a9",x"f5",x"c1"),
    61 => (x"f8",x"c1",x"87",x"c7"),
    62 => (x"db",x"c2",x"05",x"a9"),
    63 => (x"74",x"84",x"c4",x"87"),
    64 => (x"76",x"89",x"c4",x"49"),
    65 => (x"6e",x"78",x"69",x"48"),
    66 => (x"87",x"d1",x"c1",x"02"),
    67 => (x"78",x"c0",x"80",x"c8"),
    68 => (x"c0",x"48",x"a6",x"cc"),
    69 => (x"dc",x"4a",x"6e",x"78"),
    70 => (x"9a",x"cf",x"2a",x"b7"),
    71 => (x"30",x"c4",x"48",x"6e"),
    72 => (x"72",x"58",x"a6",x"c4"),
    73 => (x"87",x"c5",x"02",x"9a"),
    74 => (x"c1",x"48",x"a6",x"c8"),
    75 => (x"06",x"aa",x"c9",x"78"),
    76 => (x"f7",x"c0",x"87",x"c5"),
    77 => (x"c0",x"87",x"c3",x"82"),
    78 => (x"66",x"c8",x"82",x"f0"),
    79 => (x"72",x"87",x"c9",x"02"),
    80 => (x"87",x"f8",x"fb",x"1e"),
    81 => (x"83",x"c1",x"86",x"c4"),
    82 => (x"c1",x"48",x"66",x"cc"),
    83 => (x"58",x"a6",x"d0",x"80"),
    84 => (x"c8",x"48",x"66",x"cc"),
    85 => (x"fe",x"04",x"a8",x"b7"),
    86 => (x"d8",x"c1",x"87",x"fb"),
    87 => (x"1e",x"f0",x"c0",x"87"),
    88 => (x"c4",x"87",x"d9",x"fb"),
    89 => (x"c1",x"83",x"c1",x"86"),
    90 => (x"84",x"c4",x"87",x"cb"),
    91 => (x"89",x"c4",x"49",x"74"),
    92 => (x"e1",x"fb",x"1e",x"69"),
    93 => (x"70",x"86",x"c4",x"87"),
    94 => (x"4b",x"a3",x"71",x"49"),
    95 => (x"c4",x"87",x"f6",x"c0"),
    96 => (x"78",x"c1",x"48",x"a6"),
    97 => (x"c4",x"87",x"ee",x"c0"),
    98 => (x"c4",x"49",x"74",x"84"),
    99 => (x"fa",x"1e",x"69",x"89"),
   100 => (x"86",x"c4",x"87",x"ea"),
   101 => (x"87",x"dd",x"83",x"c1"),
   102 => (x"df",x"fa",x"1e",x"72"),
   103 => (x"d4",x"86",x"c4",x"87"),
   104 => (x"aa",x"e5",x"c0",x"87"),
   105 => (x"c4",x"87",x"c7",x"05"),
   106 => (x"78",x"c1",x"48",x"a6"),
   107 => (x"1e",x"72",x"87",x"c7"),
   108 => (x"c4",x"87",x"c9",x"fa"),
   109 => (x"66",x"e0",x"c0",x"86"),
   110 => (x"80",x"c1",x"48",x"49"),
   111 => (x"58",x"a6",x"e4",x"c0"),
   112 => (x"c0",x"fe",x"4a",x"11"),
   113 => (x"9a",x"72",x"ba",x"82"),
   114 => (x"87",x"ee",x"fb",x"05"),
   115 => (x"8e",x"f0",x"48",x"73"),
   116 => (x"4c",x"26",x"4d",x"26"),
   117 => (x"4f",x"26",x"4b",x"26"),
   118 => (x"e8",x"0e",x"5e",x"0e"),
   119 => (x"4a",x"d4",x"ff",x"86"),
   120 => (x"6a",x"7a",x"ff",x"c3"),
   121 => (x"7a",x"ff",x"c3",x"49"),
   122 => (x"30",x"c8",x"48",x"6a"),
   123 => (x"c8",x"58",x"a6",x"c4"),
   124 => (x"b1",x"6e",x"59",x"a6"),
   125 => (x"6a",x"7a",x"ff",x"c3"),
   126 => (x"cc",x"30",x"d0",x"48"),
   127 => (x"a6",x"d0",x"58",x"a6"),
   128 => (x"b1",x"66",x"c8",x"59"),
   129 => (x"6a",x"7a",x"ff",x"c3"),
   130 => (x"d4",x"30",x"d8",x"48"),
   131 => (x"a6",x"d8",x"58",x"a6"),
   132 => (x"b1",x"66",x"d0",x"59"),
   133 => (x"8e",x"e8",x"48",x"71"),
   134 => (x"5e",x"0e",x"4f",x"26"),
   135 => (x"ff",x"86",x"f4",x"0e"),
   136 => (x"ff",x"c3",x"4a",x"d4"),
   137 => (x"c3",x"49",x"6a",x"7a"),
   138 => (x"48",x"71",x"7a",x"ff"),
   139 => (x"a6",x"c4",x"30",x"c8"),
   140 => (x"6e",x"49",x"6a",x"58"),
   141 => (x"7a",x"ff",x"c3",x"b1"),
   142 => (x"30",x"c8",x"48",x"71"),
   143 => (x"6a",x"58",x"a6",x"c8"),
   144 => (x"b1",x"66",x"c4",x"49"),
   145 => (x"71",x"7a",x"ff",x"c3"),
   146 => (x"cc",x"30",x"c8",x"48"),
   147 => (x"49",x"6a",x"58",x"a6"),
   148 => (x"71",x"b1",x"66",x"c8"),
   149 => (x"26",x"8e",x"f4",x"48"),
   150 => (x"5b",x"5e",x"0e",x"4f"),
   151 => (x"c3",x"0e",x"5d",x"5c"),
   152 => (x"d4",x"ff",x"4d",x"ff"),
   153 => (x"48",x"66",x"d0",x"4c"),
   154 => (x"70",x"98",x"ff",x"c3"),
   155 => (x"c0",x"d2",x"c1",x"7c"),
   156 => (x"87",x"c8",x"05",x"bf"),
   157 => (x"c9",x"48",x"66",x"d4"),
   158 => (x"58",x"a6",x"d8",x"30"),
   159 => (x"d8",x"49",x"66",x"d4"),
   160 => (x"c3",x"48",x"71",x"29"),
   161 => (x"7c",x"70",x"98",x"ff"),
   162 => (x"d0",x"49",x"66",x"d4"),
   163 => (x"c3",x"48",x"71",x"29"),
   164 => (x"7c",x"70",x"98",x"ff"),
   165 => (x"c8",x"49",x"66",x"d4"),
   166 => (x"c3",x"48",x"71",x"29"),
   167 => (x"7c",x"70",x"98",x"ff"),
   168 => (x"c3",x"48",x"66",x"d4"),
   169 => (x"7c",x"70",x"98",x"ff"),
   170 => (x"d0",x"49",x"66",x"d0"),
   171 => (x"c3",x"48",x"71",x"29"),
   172 => (x"7c",x"70",x"98",x"ff"),
   173 => (x"f0",x"c9",x"4b",x"6c"),
   174 => (x"ab",x"75",x"4a",x"ff"),
   175 => (x"75",x"87",x"ce",x"05"),
   176 => (x"c1",x"4b",x"6c",x"7c"),
   177 => (x"87",x"c5",x"02",x"8a"),
   178 => (x"f2",x"02",x"ab",x"75"),
   179 => (x"26",x"48",x"73",x"87"),
   180 => (x"26",x"4c",x"26",x"4d"),
   181 => (x"1e",x"4f",x"26",x"4b"),
   182 => (x"d4",x"ff",x"49",x"c0"),
   183 => (x"78",x"ff",x"c3",x"48"),
   184 => (x"c8",x"c3",x"81",x"c1"),
   185 => (x"f1",x"04",x"a9",x"b7"),
   186 => (x"0e",x"4f",x"26",x"87"),
   187 => (x"5d",x"5c",x"5b",x"5e"),
   188 => (x"f0",x"ff",x"c0",x"0e"),
   189 => (x"c1",x"4d",x"f7",x"c1"),
   190 => (x"c0",x"c0",x"c0",x"c0"),
   191 => (x"d6",x"ff",x"4b",x"c0"),
   192 => (x"df",x"f8",x"c4",x"87"),
   193 => (x"75",x"1e",x"c0",x"4c"),
   194 => (x"87",x"cd",x"fd",x"1e"),
   195 => (x"a8",x"c1",x"86",x"c8"),
   196 => (x"87",x"e5",x"c0",x"05"),
   197 => (x"c3",x"48",x"d4",x"ff"),
   198 => (x"1e",x"73",x"78",x"ff"),
   199 => (x"c1",x"f0",x"e1",x"c0"),
   200 => (x"f4",x"fc",x"1e",x"e9"),
   201 => (x"70",x"86",x"c8",x"87"),
   202 => (x"87",x"ca",x"05",x"98"),
   203 => (x"c3",x"48",x"d4",x"ff"),
   204 => (x"48",x"c1",x"78",x"ff"),
   205 => (x"de",x"fe",x"87",x"cb"),
   206 => (x"05",x"8c",x"c1",x"87"),
   207 => (x"c0",x"87",x"c6",x"ff"),
   208 => (x"26",x"4d",x"26",x"48"),
   209 => (x"26",x"4b",x"26",x"4c"),
   210 => (x"5b",x"5e",x"0e",x"4f"),
   211 => (x"ff",x"c0",x"0e",x"5c"),
   212 => (x"4c",x"c1",x"c1",x"f0"),
   213 => (x"c3",x"48",x"d4",x"ff"),
   214 => (x"e5",x"c0",x"78",x"ff"),
   215 => (x"f5",x"f3",x"1e",x"e0"),
   216 => (x"d3",x"86",x"c4",x"87"),
   217 => (x"74",x"1e",x"c0",x"4b"),
   218 => (x"87",x"ed",x"fb",x"1e"),
   219 => (x"98",x"70",x"86",x"c8"),
   220 => (x"ff",x"87",x"ca",x"05"),
   221 => (x"ff",x"c3",x"48",x"d4"),
   222 => (x"cb",x"48",x"c1",x"78"),
   223 => (x"87",x"d7",x"fd",x"87"),
   224 => (x"ff",x"05",x"8b",x"c1"),
   225 => (x"48",x"c0",x"87",x"df"),
   226 => (x"4b",x"26",x"4c",x"26"),
   227 => (x"5e",x"0e",x"4f",x"26"),
   228 => (x"0e",x"5d",x"5c",x"5b"),
   229 => (x"fc",x"4c",x"d4",x"ff"),
   230 => (x"ea",x"c6",x"87",x"fd"),
   231 => (x"f0",x"e1",x"c0",x"1e"),
   232 => (x"fa",x"1e",x"c8",x"c1"),
   233 => (x"86",x"c8",x"87",x"f3"),
   234 => (x"1e",x"73",x"4b",x"70"),
   235 => (x"f3",x"1e",x"da",x"d2"),
   236 => (x"86",x"c8",x"87",x"de"),
   237 => (x"c8",x"02",x"ab",x"c1"),
   238 => (x"87",x"cd",x"fe",x"87"),
   239 => (x"cf",x"c2",x"48",x"c0"),
   240 => (x"87",x"d6",x"f9",x"87"),
   241 => (x"ff",x"cf",x"49",x"70"),
   242 => (x"ea",x"c6",x"99",x"ff"),
   243 => (x"87",x"c8",x"02",x"a9"),
   244 => (x"c0",x"87",x"f6",x"fd"),
   245 => (x"87",x"f8",x"c1",x"48"),
   246 => (x"c0",x"7c",x"ff",x"c3"),
   247 => (x"ca",x"fc",x"4d",x"f1"),
   248 => (x"02",x"98",x"70",x"87"),
   249 => (x"c0",x"87",x"d0",x"c1"),
   250 => (x"f0",x"ff",x"c0",x"1e"),
   251 => (x"f9",x"1e",x"fa",x"c1"),
   252 => (x"86",x"c8",x"87",x"e7"),
   253 => (x"9b",x"73",x"4b",x"70"),
   254 => (x"87",x"f1",x"c0",x"05"),
   255 => (x"d8",x"d1",x"1e",x"73"),
   256 => (x"87",x"cc",x"f2",x"1e"),
   257 => (x"ff",x"c3",x"86",x"c8"),
   258 => (x"73",x"4b",x"6c",x"7c"),
   259 => (x"1e",x"e4",x"d1",x"1e"),
   260 => (x"c8",x"87",x"fd",x"f1"),
   261 => (x"7c",x"ff",x"c3",x"86"),
   262 => (x"73",x"7c",x"7c",x"7c"),
   263 => (x"99",x"c0",x"c1",x"49"),
   264 => (x"c1",x"87",x"c5",x"02"),
   265 => (x"87",x"e8",x"c0",x"48"),
   266 => (x"e3",x"c0",x"48",x"c0"),
   267 => (x"d1",x"1e",x"73",x"87"),
   268 => (x"db",x"f1",x"1e",x"f2"),
   269 => (x"c2",x"86",x"c8",x"87"),
   270 => (x"87",x"cc",x"05",x"ad"),
   271 => (x"f1",x"1e",x"fe",x"d1"),
   272 => (x"86",x"c4",x"87",x"ce"),
   273 => (x"87",x"c8",x"48",x"c0"),
   274 => (x"fe",x"05",x"8d",x"c1"),
   275 => (x"48",x"c0",x"87",x"d0"),
   276 => (x"4c",x"26",x"4d",x"26"),
   277 => (x"4f",x"26",x"4b",x"26"),
   278 => (x"35",x"44",x"4d",x"43"),
   279 => (x"64",x"25",x"20",x"38"),
   280 => (x"00",x"20",x"20",x"0a"),
   281 => (x"35",x"44",x"4d",x"43"),
   282 => (x"20",x"32",x"5f",x"38"),
   283 => (x"20",x"0a",x"64",x"25"),
   284 => (x"4d",x"43",x"00",x"20"),
   285 => (x"20",x"38",x"35",x"44"),
   286 => (x"20",x"0a",x"64",x"25"),
   287 => (x"44",x"53",x"00",x"20"),
   288 => (x"49",x"20",x"43",x"48"),
   289 => (x"69",x"74",x"69",x"6e"),
   290 => (x"7a",x"69",x"6c",x"61"),
   291 => (x"6f",x"69",x"74",x"61"),
   292 => (x"72",x"65",x"20",x"6e"),
   293 => (x"21",x"72",x"6f",x"72"),
   294 => (x"6d",x"63",x"00",x"0a"),
   295 => (x"4d",x"43",x"5f",x"64"),
   296 => (x"72",x"20",x"38",x"44"),
   297 => (x"6f",x"70",x"73",x"65"),
   298 => (x"3a",x"65",x"73",x"6e"),
   299 => (x"0a",x"64",x"25",x"20"),
   300 => (x"5b",x"5e",x"0e",x"00"),
   301 => (x"fc",x"0e",x"5d",x"5c"),
   302 => (x"4c",x"d0",x"ff",x"86"),
   303 => (x"4b",x"c0",x"c0",x"c8"),
   304 => (x"48",x"c0",x"d2",x"c1"),
   305 => (x"da",x"d6",x"78",x"c1"),
   306 => (x"87",x"ca",x"ee",x"1e"),
   307 => (x"4d",x"c7",x"86",x"c4"),
   308 => (x"98",x"73",x"48",x"6c"),
   309 => (x"6e",x"58",x"a6",x"c4"),
   310 => (x"6c",x"87",x"cc",x"02"),
   311 => (x"c4",x"98",x"73",x"48"),
   312 => (x"05",x"6e",x"58",x"a6"),
   313 => (x"c0",x"87",x"f4",x"ff"),
   314 => (x"87",x"eb",x"f7",x"7c"),
   315 => (x"98",x"73",x"48",x"6c"),
   316 => (x"6e",x"58",x"a6",x"c4"),
   317 => (x"6c",x"87",x"cc",x"02"),
   318 => (x"c4",x"98",x"73",x"48"),
   319 => (x"05",x"6e",x"58",x"a6"),
   320 => (x"c1",x"87",x"f4",x"ff"),
   321 => (x"c0",x"1e",x"c0",x"7c"),
   322 => (x"c0",x"c1",x"d0",x"e5"),
   323 => (x"87",x"c9",x"f5",x"1e"),
   324 => (x"a8",x"c1",x"86",x"c8"),
   325 => (x"87",x"c2",x"c0",x"05"),
   326 => (x"ad",x"c2",x"4d",x"c1"),
   327 => (x"87",x"cd",x"c0",x"05"),
   328 => (x"ec",x"1e",x"d5",x"d6"),
   329 => (x"86",x"c4",x"87",x"f0"),
   330 => (x"de",x"c1",x"48",x"c0"),
   331 => (x"05",x"8d",x"c1",x"87"),
   332 => (x"f9",x"87",x"dd",x"fe"),
   333 => (x"d2",x"c1",x"87",x"d8"),
   334 => (x"d2",x"c1",x"58",x"c4"),
   335 => (x"c0",x"05",x"bf",x"c0"),
   336 => (x"1e",x"c1",x"87",x"cd"),
   337 => (x"c1",x"f0",x"ff",x"c0"),
   338 => (x"cc",x"f4",x"1e",x"d0"),
   339 => (x"ff",x"86",x"c8",x"87"),
   340 => (x"ff",x"c3",x"48",x"d4"),
   341 => (x"87",x"ca",x"ca",x"78"),
   342 => (x"58",x"c8",x"d2",x"c1"),
   343 => (x"bf",x"c4",x"d2",x"c1"),
   344 => (x"1e",x"de",x"d6",x"1e"),
   345 => (x"c8",x"87",x"e9",x"ec"),
   346 => (x"73",x"48",x"6c",x"86"),
   347 => (x"58",x"a6",x"c4",x"98"),
   348 => (x"cc",x"c0",x"02",x"6e"),
   349 => (x"73",x"48",x"6c",x"87"),
   350 => (x"58",x"a6",x"c4",x"98"),
   351 => (x"f4",x"ff",x"05",x"6e"),
   352 => (x"ff",x"7c",x"c0",x"87"),
   353 => (x"ff",x"c3",x"48",x"d4"),
   354 => (x"fc",x"48",x"c1",x"78"),
   355 => (x"26",x"4d",x"26",x"8e"),
   356 => (x"26",x"4b",x"26",x"4c"),
   357 => (x"52",x"45",x"49",x"4f"),
   358 => (x"50",x"53",x"00",x"52"),
   359 => (x"44",x"53",x"00",x"49"),
   360 => (x"72",x"61",x"63",x"20"),
   361 => (x"69",x"73",x"20",x"64"),
   362 => (x"69",x"20",x"65",x"7a"),
   363 => (x"64",x"25",x"20",x"73"),
   364 => (x"5e",x"0e",x"00",x"0a"),
   365 => (x"0e",x"5d",x"5c",x"5b"),
   366 => (x"c0",x"c8",x"86",x"fc"),
   367 => (x"ff",x"c3",x"4d",x"c0"),
   368 => (x"4b",x"d4",x"ff",x"4c"),
   369 => (x"d0",x"ff",x"7b",x"74"),
   370 => (x"98",x"75",x"48",x"bf"),
   371 => (x"6e",x"58",x"a6",x"c4"),
   372 => (x"87",x"ce",x"c0",x"02"),
   373 => (x"48",x"bf",x"d0",x"ff"),
   374 => (x"a6",x"c4",x"98",x"75"),
   375 => (x"ff",x"05",x"6e",x"58"),
   376 => (x"d0",x"ff",x"87",x"f2"),
   377 => (x"78",x"c1",x"c4",x"48"),
   378 => (x"66",x"d4",x"7b",x"74"),
   379 => (x"f0",x"ff",x"c0",x"1e"),
   380 => (x"f1",x"1e",x"d8",x"c1"),
   381 => (x"86",x"c8",x"87",x"e3"),
   382 => (x"c0",x"02",x"98",x"70"),
   383 => (x"da",x"da",x"87",x"cd"),
   384 => (x"87",x"d2",x"e9",x"1e"),
   385 => (x"48",x"c1",x"86",x"c4"),
   386 => (x"74",x"87",x"c5",x"c2"),
   387 => (x"7b",x"fe",x"c3",x"7b"),
   388 => (x"78",x"c0",x"48",x"76"),
   389 => (x"25",x"4d",x"66",x"d8"),
   390 => (x"d8",x"4a",x"71",x"49"),
   391 => (x"48",x"72",x"2a",x"b7"),
   392 => (x"7b",x"70",x"98",x"74"),
   393 => (x"b7",x"d0",x"4a",x"71"),
   394 => (x"74",x"48",x"72",x"2a"),
   395 => (x"71",x"7b",x"70",x"98"),
   396 => (x"2a",x"b7",x"c8",x"4a"),
   397 => (x"98",x"74",x"48",x"72"),
   398 => (x"48",x"71",x"7b",x"70"),
   399 => (x"7b",x"70",x"98",x"74"),
   400 => (x"80",x"c1",x"48",x"6e"),
   401 => (x"6e",x"58",x"a6",x"c4"),
   402 => (x"b7",x"c0",x"c2",x"48"),
   403 => (x"c6",x"ff",x"04",x"a8"),
   404 => (x"c0",x"c0",x"c8",x"87"),
   405 => (x"74",x"7b",x"74",x"4d"),
   406 => (x"d8",x"7b",x"74",x"7b"),
   407 => (x"74",x"49",x"e0",x"da"),
   408 => (x"c0",x"05",x"6b",x"7b"),
   409 => (x"89",x"c1",x"87",x"c6"),
   410 => (x"87",x"f3",x"ff",x"05"),
   411 => (x"d0",x"ff",x"7b",x"74"),
   412 => (x"98",x"75",x"48",x"bf"),
   413 => (x"6e",x"58",x"a6",x"c4"),
   414 => (x"87",x"ce",x"c0",x"02"),
   415 => (x"48",x"bf",x"d0",x"ff"),
   416 => (x"a6",x"c4",x"98",x"75"),
   417 => (x"ff",x"05",x"6e",x"58"),
   418 => (x"d0",x"ff",x"87",x"f2"),
   419 => (x"48",x"78",x"c0",x"48"),
   420 => (x"4d",x"26",x"8e",x"fc"),
   421 => (x"4b",x"26",x"4c",x"26"),
   422 => (x"72",x"57",x"4f",x"26"),
   423 => (x"20",x"65",x"74",x"69"),
   424 => (x"6c",x"69",x"61",x"66"),
   425 => (x"00",x"0a",x"64",x"65"),
   426 => (x"5c",x"5b",x"5e",x"0e"),
   427 => (x"d4",x"ff",x"0e",x"5d"),
   428 => (x"4c",x"66",x"d4",x"4d"),
   429 => (x"c0",x"4b",x"66",x"d0"),
   430 => (x"cd",x"ee",x"c5",x"4a"),
   431 => (x"ff",x"c3",x"49",x"df"),
   432 => (x"c3",x"48",x"6d",x"7d"),
   433 => (x"c1",x"05",x"a8",x"fe"),
   434 => (x"d1",x"c1",x"87",x"d4"),
   435 => (x"78",x"c0",x"48",x"fc"),
   436 => (x"04",x"ac",x"b7",x"c4"),
   437 => (x"eb",x"87",x"dc",x"c0"),
   438 => (x"49",x"70",x"87",x"fe"),
   439 => (x"83",x"c4",x"7b",x"71"),
   440 => (x"bf",x"fc",x"d1",x"c1"),
   441 => (x"c1",x"80",x"71",x"48"),
   442 => (x"c4",x"58",x"c0",x"d2"),
   443 => (x"03",x"ac",x"b7",x"8c"),
   444 => (x"c0",x"87",x"e4",x"ff"),
   445 => (x"c0",x"06",x"ac",x"b7"),
   446 => (x"ff",x"c3",x"87",x"e1"),
   447 => (x"71",x"49",x"6d",x"7d"),
   448 => (x"ff",x"c3",x"7b",x"97"),
   449 => (x"c1",x"83",x"c1",x"98"),
   450 => (x"48",x"bf",x"fc",x"d1"),
   451 => (x"d2",x"c1",x"80",x"71"),
   452 => (x"8c",x"c1",x"58",x"c0"),
   453 => (x"01",x"ac",x"b7",x"c0"),
   454 => (x"c1",x"87",x"df",x"ff"),
   455 => (x"89",x"c1",x"4a",x"49"),
   456 => (x"87",x"da",x"fe",x"05"),
   457 => (x"72",x"7d",x"ff",x"c3"),
   458 => (x"26",x"4d",x"26",x"48"),
   459 => (x"26",x"4b",x"26",x"4c"),
   460 => (x"5b",x"5e",x"0e",x"4f"),
   461 => (x"fc",x"0e",x"5d",x"5c"),
   462 => (x"4c",x"d0",x"ff",x"86"),
   463 => (x"4b",x"c0",x"c0",x"c8"),
   464 => (x"d4",x"ff",x"4d",x"c0"),
   465 => (x"78",x"ff",x"c3",x"48"),
   466 => (x"98",x"73",x"48",x"6c"),
   467 => (x"6e",x"58",x"a6",x"c4"),
   468 => (x"87",x"cc",x"c0",x"02"),
   469 => (x"98",x"73",x"48",x"6c"),
   470 => (x"6e",x"58",x"a6",x"c4"),
   471 => (x"87",x"f4",x"ff",x"05"),
   472 => (x"ff",x"7c",x"c1",x"c4"),
   473 => (x"ff",x"c3",x"48",x"d4"),
   474 => (x"1e",x"66",x"d4",x"78"),
   475 => (x"c1",x"f0",x"ff",x"c0"),
   476 => (x"e4",x"eb",x"1e",x"d1"),
   477 => (x"70",x"86",x"c8",x"87"),
   478 => (x"02",x"99",x"71",x"49"),
   479 => (x"71",x"87",x"d0",x"c0"),
   480 => (x"1e",x"66",x"d8",x"1e"),
   481 => (x"e4",x"1e",x"c2",x"df"),
   482 => (x"86",x"cc",x"87",x"c6"),
   483 => (x"c8",x"87",x"e7",x"c0"),
   484 => (x"66",x"dc",x"1e",x"c0"),
   485 => (x"87",x"d0",x"fc",x"1e"),
   486 => (x"4d",x"70",x"86",x"c8"),
   487 => (x"98",x"73",x"48",x"6c"),
   488 => (x"6e",x"58",x"a6",x"c4"),
   489 => (x"87",x"cc",x"c0",x"02"),
   490 => (x"98",x"73",x"48",x"6c"),
   491 => (x"6e",x"58",x"a6",x"c4"),
   492 => (x"87",x"f4",x"ff",x"05"),
   493 => (x"48",x"75",x"7c",x"c0"),
   494 => (x"4d",x"26",x"8e",x"fc"),
   495 => (x"4b",x"26",x"4c",x"26"),
   496 => (x"65",x"52",x"4f",x"26"),
   497 => (x"63",x"20",x"64",x"61"),
   498 => (x"61",x"6d",x"6d",x"6f"),
   499 => (x"66",x"20",x"64",x"6e"),
   500 => (x"65",x"6c",x"69",x"61"),
   501 => (x"74",x"61",x"20",x"64"),
   502 => (x"20",x"64",x"25",x"20"),
   503 => (x"29",x"64",x"25",x"28"),
   504 => (x"5e",x"0e",x"00",x"0a"),
   505 => (x"0e",x"5d",x"5c",x"5b"),
   506 => (x"1e",x"c0",x"86",x"fc"),
   507 => (x"c1",x"f0",x"ff",x"c0"),
   508 => (x"e4",x"e9",x"1e",x"c9"),
   509 => (x"d2",x"86",x"c8",x"87"),
   510 => (x"ce",x"d2",x"c1",x"1e"),
   511 => (x"87",x"e8",x"fa",x"1e"),
   512 => (x"4d",x"c0",x"86",x"c8"),
   513 => (x"b7",x"d2",x"85",x"c1"),
   514 => (x"f7",x"ff",x"04",x"ad"),
   515 => (x"ce",x"d2",x"c1",x"87"),
   516 => (x"c3",x"49",x"bf",x"97"),
   517 => (x"c0",x"c1",x"99",x"c0"),
   518 => (x"e8",x"c0",x"05",x"a9"),
   519 => (x"d5",x"d2",x"c1",x"87"),
   520 => (x"d0",x"49",x"bf",x"97"),
   521 => (x"d6",x"d2",x"c1",x"31"),
   522 => (x"c8",x"4a",x"bf",x"97"),
   523 => (x"c1",x"b1",x"72",x"32"),
   524 => (x"bf",x"97",x"d7",x"d2"),
   525 => (x"cf",x"b1",x"72",x"4a"),
   526 => (x"99",x"ff",x"ff",x"ff"),
   527 => (x"85",x"c1",x"4d",x"71"),
   528 => (x"eb",x"c2",x"35",x"ca"),
   529 => (x"d7",x"d2",x"c1",x"87"),
   530 => (x"c1",x"4b",x"bf",x"97"),
   531 => (x"c1",x"9b",x"c6",x"33"),
   532 => (x"bf",x"97",x"d8",x"d2"),
   533 => (x"29",x"b7",x"c7",x"49"),
   534 => (x"d2",x"c1",x"b3",x"71"),
   535 => (x"49",x"bf",x"97",x"d3"),
   536 => (x"98",x"cf",x"48",x"71"),
   537 => (x"c1",x"58",x"a6",x"c4"),
   538 => (x"bf",x"97",x"d4",x"d2"),
   539 => (x"ca",x"9c",x"c3",x"4c"),
   540 => (x"d5",x"d2",x"c1",x"34"),
   541 => (x"c2",x"49",x"bf",x"97"),
   542 => (x"c1",x"b4",x"71",x"31"),
   543 => (x"bf",x"97",x"d6",x"d2"),
   544 => (x"99",x"c0",x"c3",x"49"),
   545 => (x"71",x"29",x"b7",x"c6"),
   546 => (x"c4",x"1e",x"74",x"b4"),
   547 => (x"1e",x"73",x"1e",x"66"),
   548 => (x"1e",x"fc",x"e3",x"c0"),
   549 => (x"87",x"f8",x"df",x"ff"),
   550 => (x"83",x"c2",x"86",x"d0"),
   551 => (x"30",x"73",x"48",x"c1"),
   552 => (x"1e",x"73",x"4b",x"70"),
   553 => (x"1e",x"e9",x"e4",x"c0"),
   554 => (x"87",x"e4",x"df",x"ff"),
   555 => (x"48",x"c1",x"86",x"c8"),
   556 => (x"a6",x"c4",x"30",x"6e"),
   557 => (x"c1",x"49",x"74",x"58"),
   558 => (x"73",x"4d",x"71",x"81"),
   559 => (x"1e",x"6e",x"95",x"b7"),
   560 => (x"e4",x"c0",x"1e",x"75"),
   561 => (x"df",x"ff",x"1e",x"f2"),
   562 => (x"86",x"cc",x"87",x"c6"),
   563 => (x"c0",x"c8",x"48",x"6e"),
   564 => (x"c0",x"06",x"a8",x"b7"),
   565 => (x"4b",x"6e",x"87",x"ce"),
   566 => (x"2b",x"b7",x"35",x"c1"),
   567 => (x"ab",x"b7",x"c0",x"c8"),
   568 => (x"87",x"f4",x"ff",x"01"),
   569 => (x"e5",x"c0",x"1e",x"75"),
   570 => (x"de",x"ff",x"1e",x"c8"),
   571 => (x"86",x"c8",x"87",x"e2"),
   572 => (x"8e",x"fc",x"48",x"75"),
   573 => (x"4c",x"26",x"4d",x"26"),
   574 => (x"4f",x"26",x"4b",x"26"),
   575 => (x"69",x"73",x"5f",x"63"),
   576 => (x"6d",x"5f",x"65",x"7a"),
   577 => (x"3a",x"74",x"6c",x"75"),
   578 => (x"2c",x"64",x"25",x"20"),
   579 => (x"61",x"65",x"72",x"20"),
   580 => (x"6c",x"62",x"5f",x"64"),
   581 => (x"6e",x"65",x"6c",x"5f"),
   582 => (x"64",x"25",x"20",x"3a"),
   583 => (x"73",x"63",x"20",x"2c"),
   584 => (x"3a",x"65",x"7a",x"69"),
   585 => (x"0a",x"64",x"25",x"20"),
   586 => (x"6c",x"75",x"4d",x"00"),
   587 => (x"64",x"25",x"20",x"74"),
   588 => (x"64",x"25",x"00",x"0a"),
   589 => (x"6f",x"6c",x"62",x"20"),
   590 => (x"20",x"73",x"6b",x"63"),
   591 => (x"73",x"20",x"66",x"6f"),
   592 => (x"20",x"65",x"7a",x"69"),
   593 => (x"00",x"0a",x"64",x"25"),
   594 => (x"62",x"20",x"64",x"25"),
   595 => (x"6b",x"63",x"6f",x"6c"),
   596 => (x"66",x"6f",x"20",x"73"),
   597 => (x"32",x"31",x"35",x"20"),
   598 => (x"74",x"79",x"62",x"20"),
   599 => (x"00",x"0a",x"73",x"65"),
   600 => (x"00",x"44",x"4d",x"43"),
   601 => (x"c0",x"1e",x"73",x"1e"),
   602 => (x"48",x"66",x"d0",x"4b"),
   603 => (x"06",x"a8",x"b7",x"c0"),
   604 => (x"c8",x"87",x"f6",x"c0"),
   605 => (x"4a",x"bf",x"97",x"66"),
   606 => (x"ba",x"82",x"c0",x"fe"),
   607 => (x"c1",x"48",x"66",x"c8"),
   608 => (x"58",x"a6",x"cc",x"80"),
   609 => (x"bf",x"97",x"66",x"cc"),
   610 => (x"81",x"c0",x"fe",x"49"),
   611 => (x"48",x"66",x"cc",x"b9"),
   612 => (x"a6",x"d0",x"80",x"c1"),
   613 => (x"aa",x"b7",x"71",x"58"),
   614 => (x"c1",x"87",x"c4",x"02"),
   615 => (x"c1",x"87",x"cc",x"48"),
   616 => (x"b7",x"66",x"d0",x"83"),
   617 => (x"ca",x"ff",x"04",x"ab"),
   618 => (x"c4",x"48",x"c0",x"87"),
   619 => (x"26",x"4d",x"26",x"87"),
   620 => (x"26",x"4b",x"26",x"4c"),
   621 => (x"5b",x"5e",x"0e",x"4f"),
   622 => (x"c1",x"0e",x"5d",x"5c"),
   623 => (x"c0",x"48",x"e8",x"da"),
   624 => (x"d9",x"f6",x"c0",x"78"),
   625 => (x"cd",x"da",x"ff",x"1e"),
   626 => (x"c1",x"86",x"c4",x"87"),
   627 => (x"c0",x"1e",x"e0",x"d2"),
   628 => (x"87",x"dd",x"f5",x"1e"),
   629 => (x"98",x"70",x"86",x"c8"),
   630 => (x"c0",x"87",x"cf",x"05"),
   631 => (x"ff",x"1e",x"c5",x"f3"),
   632 => (x"c4",x"87",x"f3",x"d9"),
   633 => (x"cb",x"48",x"c0",x"86"),
   634 => (x"f6",x"c0",x"87",x"d8"),
   635 => (x"d9",x"ff",x"1e",x"e6"),
   636 => (x"86",x"c4",x"87",x"e4"),
   637 => (x"db",x"c1",x"4b",x"c0"),
   638 => (x"78",x"c1",x"48",x"d4"),
   639 => (x"f6",x"c0",x"1e",x"c8"),
   640 => (x"d3",x"c1",x"1e",x"fd"),
   641 => (x"db",x"fd",x"1e",x"d6"),
   642 => (x"70",x"86",x"cc",x"87"),
   643 => (x"87",x"c6",x"05",x"98"),
   644 => (x"48",x"d4",x"db",x"c1"),
   645 => (x"1e",x"c8",x"78",x"c0"),
   646 => (x"1e",x"c6",x"f7",x"c0"),
   647 => (x"1e",x"f2",x"d3",x"c1"),
   648 => (x"cc",x"87",x"c1",x"fd"),
   649 => (x"05",x"98",x"70",x"86"),
   650 => (x"db",x"c1",x"87",x"c6"),
   651 => (x"78",x"c0",x"48",x"d4"),
   652 => (x"bf",x"d4",x"db",x"c1"),
   653 => (x"cf",x"f7",x"c0",x"1e"),
   654 => (x"d3",x"d9",x"ff",x"1e"),
   655 => (x"c1",x"86",x"c8",x"87"),
   656 => (x"02",x"bf",x"d4",x"db"),
   657 => (x"c1",x"87",x"d5",x"c2"),
   658 => (x"c1",x"4d",x"e0",x"d2"),
   659 => (x"c1",x"4c",x"de",x"d9"),
   660 => (x"bf",x"9f",x"de",x"da"),
   661 => (x"c1",x"1e",x"71",x"49"),
   662 => (x"c1",x"49",x"de",x"da"),
   663 => (x"71",x"89",x"e0",x"d2"),
   664 => (x"c8",x"1e",x"d0",x"1e"),
   665 => (x"f3",x"c0",x"1e",x"c0"),
   666 => (x"d8",x"ff",x"1e",x"f7"),
   667 => (x"86",x"d4",x"87",x"e2"),
   668 => (x"69",x"49",x"a4",x"c8"),
   669 => (x"de",x"da",x"c1",x"4b"),
   670 => (x"c5",x"49",x"bf",x"9f"),
   671 => (x"05",x"a9",x"ea",x"d6"),
   672 => (x"c8",x"87",x"cf",x"c0"),
   673 => (x"1e",x"69",x"49",x"a4"),
   674 => (x"c4",x"87",x"ff",x"d8"),
   675 => (x"c0",x"4b",x"70",x"86"),
   676 => (x"fe",x"c7",x"87",x"de"),
   677 => (x"69",x"9f",x"49",x"a5"),
   678 => (x"d5",x"e9",x"ca",x"49"),
   679 => (x"cf",x"c0",x"02",x"a9"),
   680 => (x"d9",x"f3",x"c0",x"87"),
   681 => (x"ed",x"d6",x"ff",x"1e"),
   682 => (x"c0",x"86",x"c4",x"87"),
   683 => (x"87",x"d2",x"c8",x"48"),
   684 => (x"f4",x"c0",x"1e",x"73"),
   685 => (x"d7",x"ff",x"1e",x"f4"),
   686 => (x"86",x"c8",x"87",x"d6"),
   687 => (x"1e",x"e0",x"d2",x"c1"),
   688 => (x"ec",x"f1",x"1e",x"73"),
   689 => (x"70",x"86",x"c8",x"87"),
   690 => (x"c5",x"c0",x"05",x"98"),
   691 => (x"c7",x"48",x"c0",x"87"),
   692 => (x"f5",x"c0",x"87",x"f0"),
   693 => (x"d5",x"ff",x"1e",x"cc"),
   694 => (x"86",x"c4",x"87",x"fc"),
   695 => (x"1e",x"e2",x"f7",x"c0"),
   696 => (x"87",x"ec",x"d6",x"ff"),
   697 => (x"1e",x"c8",x"86",x"c4"),
   698 => (x"1e",x"fa",x"f7",x"c0"),
   699 => (x"1e",x"f2",x"d3",x"c1"),
   700 => (x"cc",x"87",x"f1",x"f9"),
   701 => (x"05",x"98",x"70",x"86"),
   702 => (x"c1",x"87",x"c9",x"c0"),
   703 => (x"c1",x"48",x"e8",x"da"),
   704 => (x"87",x"e4",x"c0",x"78"),
   705 => (x"f8",x"c0",x"1e",x"c8"),
   706 => (x"d3",x"c1",x"1e",x"c3"),
   707 => (x"d3",x"f9",x"1e",x"d6"),
   708 => (x"70",x"86",x"cc",x"87"),
   709 => (x"cf",x"c0",x"02",x"98"),
   710 => (x"f3",x"f5",x"c0",x"87"),
   711 => (x"ef",x"d5",x"ff",x"1e"),
   712 => (x"c0",x"86",x"c4",x"87"),
   713 => (x"87",x"da",x"c6",x"48"),
   714 => (x"97",x"de",x"da",x"c1"),
   715 => (x"d5",x"c1",x"49",x"bf"),
   716 => (x"cd",x"c0",x"05",x"a9"),
   717 => (x"df",x"da",x"c1",x"87"),
   718 => (x"c2",x"49",x"bf",x"97"),
   719 => (x"c0",x"02",x"a9",x"ea"),
   720 => (x"48",x"c0",x"87",x"c5"),
   721 => (x"c1",x"87",x"fb",x"c5"),
   722 => (x"bf",x"97",x"e0",x"d2"),
   723 => (x"a9",x"e9",x"c3",x"49"),
   724 => (x"87",x"d2",x"c0",x"02"),
   725 => (x"97",x"e0",x"d2",x"c1"),
   726 => (x"eb",x"c3",x"49",x"bf"),
   727 => (x"c5",x"c0",x"02",x"a9"),
   728 => (x"c5",x"48",x"c0",x"87"),
   729 => (x"d2",x"c1",x"87",x"dc"),
   730 => (x"49",x"bf",x"97",x"eb"),
   731 => (x"c0",x"05",x"99",x"71"),
   732 => (x"d2",x"c1",x"87",x"cc"),
   733 => (x"49",x"bf",x"97",x"ec"),
   734 => (x"c0",x"02",x"a9",x"c2"),
   735 => (x"48",x"c0",x"87",x"c5"),
   736 => (x"c1",x"87",x"ff",x"c4"),
   737 => (x"bf",x"97",x"ed",x"d2"),
   738 => (x"e4",x"da",x"c1",x"48"),
   739 => (x"e0",x"da",x"c1",x"58"),
   740 => (x"4a",x"71",x"49",x"bf"),
   741 => (x"da",x"c1",x"8a",x"c1"),
   742 => (x"1e",x"72",x"5a",x"e8"),
   743 => (x"f8",x"c0",x"1e",x"71"),
   744 => (x"d3",x"ff",x"1e",x"cc"),
   745 => (x"86",x"cc",x"87",x"ea"),
   746 => (x"97",x"ee",x"d2",x"c1"),
   747 => (x"81",x"73",x"49",x"bf"),
   748 => (x"97",x"ef",x"d2",x"c1"),
   749 => (x"32",x"c8",x"4a",x"bf"),
   750 => (x"48",x"f4",x"da",x"c1"),
   751 => (x"c1",x"78",x"a1",x"72"),
   752 => (x"bf",x"97",x"f0",x"d2"),
   753 => (x"cc",x"db",x"c1",x"48"),
   754 => (x"e8",x"da",x"c1",x"58"),
   755 => (x"df",x"c2",x"02",x"bf"),
   756 => (x"c0",x"1e",x"c8",x"87"),
   757 => (x"c1",x"1e",x"d0",x"f6"),
   758 => (x"f6",x"1e",x"f2",x"d3"),
   759 => (x"86",x"cc",x"87",x"c6"),
   760 => (x"c0",x"02",x"98",x"70"),
   761 => (x"48",x"c0",x"87",x"c5"),
   762 => (x"c1",x"87",x"d7",x"c3"),
   763 => (x"4a",x"bf",x"e0",x"da"),
   764 => (x"30",x"c4",x"48",x"72"),
   765 => (x"58",x"d0",x"db",x"c1"),
   766 => (x"5a",x"c8",x"db",x"c1"),
   767 => (x"97",x"c5",x"d3",x"c1"),
   768 => (x"31",x"c8",x"49",x"bf"),
   769 => (x"97",x"c4",x"d3",x"c1"),
   770 => (x"a1",x"73",x"4b",x"bf"),
   771 => (x"c6",x"d3",x"c1",x"49"),
   772 => (x"d0",x"4b",x"bf",x"97"),
   773 => (x"49",x"a1",x"73",x"33"),
   774 => (x"97",x"c7",x"d3",x"c1"),
   775 => (x"33",x"d8",x"4b",x"bf"),
   776 => (x"c1",x"49",x"a1",x"73"),
   777 => (x"c1",x"59",x"d4",x"db"),
   778 => (x"91",x"bf",x"c8",x"db"),
   779 => (x"bf",x"f4",x"da",x"c1"),
   780 => (x"fc",x"da",x"c1",x"81"),
   781 => (x"cd",x"d3",x"c1",x"59"),
   782 => (x"c8",x"4b",x"bf",x"97"),
   783 => (x"cc",x"d3",x"c1",x"33"),
   784 => (x"74",x"4c",x"bf",x"97"),
   785 => (x"d3",x"c1",x"4b",x"a3"),
   786 => (x"4c",x"bf",x"97",x"ce"),
   787 => (x"a3",x"74",x"34",x"d0"),
   788 => (x"cf",x"d3",x"c1",x"4b"),
   789 => (x"cf",x"4c",x"bf",x"97"),
   790 => (x"74",x"34",x"d8",x"9c"),
   791 => (x"db",x"c1",x"4b",x"a3"),
   792 => (x"8b",x"c2",x"5b",x"c0"),
   793 => (x"db",x"c1",x"92",x"73"),
   794 => (x"a1",x"72",x"48",x"c0"),
   795 => (x"87",x"d0",x"c1",x"78"),
   796 => (x"97",x"f2",x"d2",x"c1"),
   797 => (x"31",x"c8",x"49",x"bf"),
   798 => (x"97",x"f1",x"d2",x"c1"),
   799 => (x"a1",x"72",x"4a",x"bf"),
   800 => (x"d0",x"db",x"c1",x"49"),
   801 => (x"c7",x"31",x"c5",x"59"),
   802 => (x"29",x"c9",x"81",x"ff"),
   803 => (x"59",x"c8",x"db",x"c1"),
   804 => (x"97",x"f7",x"d2",x"c1"),
   805 => (x"32",x"c8",x"4a",x"bf"),
   806 => (x"97",x"f6",x"d2",x"c1"),
   807 => (x"a2",x"73",x"4b",x"bf"),
   808 => (x"d4",x"db",x"c1",x"4a"),
   809 => (x"c8",x"db",x"c1",x"5a"),
   810 => (x"da",x"c1",x"92",x"bf"),
   811 => (x"c1",x"82",x"bf",x"f4"),
   812 => (x"c1",x"5a",x"c4",x"db"),
   813 => (x"c0",x"48",x"fc",x"da"),
   814 => (x"f8",x"da",x"c1",x"78"),
   815 => (x"78",x"a1",x"72",x"48"),
   816 => (x"e8",x"f3",x"48",x"c1"),
   817 => (x"61",x"65",x"52",x"87"),
   818 => (x"66",x"6f",x"20",x"64"),
   819 => (x"52",x"42",x"4d",x"20"),
   820 => (x"69",x"61",x"66",x"20"),
   821 => (x"0a",x"64",x"65",x"6c"),
   822 => (x"20",x"6f",x"4e",x"00"),
   823 => (x"74",x"72",x"61",x"70"),
   824 => (x"6f",x"69",x"74",x"69"),
   825 => (x"69",x"73",x"20",x"6e"),
   826 => (x"74",x"61",x"6e",x"67"),
   827 => (x"20",x"65",x"72",x"75"),
   828 => (x"6e",x"75",x"6f",x"66"),
   829 => (x"4d",x"00",x"0a",x"64"),
   830 => (x"69",x"73",x"52",x"42"),
   831 => (x"20",x"3a",x"65",x"7a"),
   832 => (x"20",x"2c",x"64",x"25"),
   833 => (x"74",x"72",x"61",x"70"),
   834 => (x"6f",x"69",x"74",x"69"),
   835 => (x"7a",x"69",x"73",x"6e"),
   836 => (x"25",x"20",x"3a",x"65"),
   837 => (x"6f",x"20",x"2c",x"64"),
   838 => (x"65",x"73",x"66",x"66"),
   839 => (x"66",x"6f",x"20",x"74"),
   840 => (x"67",x"69",x"73",x"20"),
   841 => (x"64",x"25",x"20",x"3a"),
   842 => (x"69",x"73",x"20",x"2c"),
   843 => (x"78",x"30",x"20",x"67"),
   844 => (x"00",x"0a",x"78",x"25"),
   845 => (x"64",x"61",x"65",x"52"),
   846 => (x"20",x"67",x"6e",x"69"),
   847 => (x"74",x"6f",x"6f",x"62"),
   848 => (x"63",x"65",x"73",x"20"),
   849 => (x"20",x"72",x"6f",x"74"),
   850 => (x"00",x"0a",x"64",x"25"),
   851 => (x"64",x"61",x"65",x"52"),
   852 => (x"6f",x"6f",x"62",x"20"),
   853 => (x"65",x"73",x"20",x"74"),
   854 => (x"72",x"6f",x"74",x"63"),
   855 => (x"6f",x"72",x"66",x"20"),
   856 => (x"69",x"66",x"20",x"6d"),
   857 => (x"20",x"74",x"73",x"72"),
   858 => (x"74",x"72",x"61",x"70"),
   859 => (x"6f",x"69",x"74",x"69"),
   860 => (x"55",x"00",x"0a",x"6e"),
   861 => (x"70",x"75",x"73",x"6e"),
   862 => (x"74",x"72",x"6f",x"70"),
   863 => (x"70",x"20",x"64",x"65"),
   864 => (x"69",x"74",x"72",x"61"),
   865 => (x"6e",x"6f",x"69",x"74"),
   866 => (x"70",x"79",x"74",x"20"),
   867 => (x"00",x"0d",x"21",x"65"),
   868 => (x"33",x"54",x"41",x"46"),
   869 => (x"20",x"20",x"20",x"32"),
   870 => (x"61",x"65",x"52",x"00"),
   871 => (x"67",x"6e",x"69",x"64"),
   872 => (x"52",x"42",x"4d",x"20"),
   873 => (x"42",x"4d",x"00",x"0a"),
   874 => (x"75",x"73",x"20",x"52"),
   875 => (x"73",x"65",x"63",x"63"),
   876 => (x"6c",x"75",x"66",x"73"),
   877 => (x"72",x"20",x"79",x"6c"),
   878 => (x"0a",x"64",x"61",x"65"),
   879 => (x"54",x"41",x"46",x"00"),
   880 => (x"20",x"20",x"36",x"31"),
   881 => (x"41",x"46",x"00",x"20"),
   882 => (x"20",x"32",x"33",x"54"),
   883 => (x"50",x"00",x"20",x"20"),
   884 => (x"69",x"74",x"72",x"61"),
   885 => (x"6e",x"6f",x"69",x"74"),
   886 => (x"6e",x"75",x"6f",x"63"),
   887 => (x"64",x"25",x"20",x"74"),
   888 => (x"75",x"48",x"00",x"0a"),
   889 => (x"6e",x"69",x"74",x"6e"),
   890 => (x"6f",x"66",x"20",x"67"),
   891 => (x"69",x"66",x"20",x"72"),
   892 => (x"79",x"73",x"65",x"6c"),
   893 => (x"6d",x"65",x"74",x"73"),
   894 => (x"41",x"46",x"00",x"0a"),
   895 => (x"20",x"32",x"33",x"54"),
   896 => (x"46",x"00",x"20",x"20"),
   897 => (x"36",x"31",x"54",x"41"),
   898 => (x"00",x"20",x"20",x"20"),
   899 => (x"73",x"75",x"6c",x"43"),
   900 => (x"20",x"72",x"65",x"74"),
   901 => (x"65",x"7a",x"69",x"73"),
   902 => (x"64",x"25",x"20",x"3a"),
   903 => (x"6c",x"43",x"20",x"2c"),
   904 => (x"65",x"74",x"73",x"75"),
   905 => (x"61",x"6d",x"20",x"72"),
   906 => (x"20",x"2c",x"6b",x"73"),
   907 => (x"00",x"0a",x"64",x"25"),
   908 => (x"5c",x"5b",x"5e",x"0e"),
   909 => (x"e8",x"da",x"c1",x"0e"),
   910 => (x"87",x"ce",x"02",x"bf"),
   911 => (x"c7",x"4a",x"66",x"cc"),
   912 => (x"66",x"cc",x"2a",x"b7"),
   913 => (x"9b",x"ff",x"c1",x"4b"),
   914 => (x"66",x"cc",x"87",x"cc"),
   915 => (x"2a",x"b7",x"c8",x"4a"),
   916 => (x"c3",x"4b",x"66",x"cc"),
   917 => (x"d2",x"c1",x"9b",x"ff"),
   918 => (x"da",x"c1",x"1e",x"e0"),
   919 => (x"72",x"49",x"bf",x"f4"),
   920 => (x"e3",x"1e",x"71",x"81"),
   921 => (x"86",x"c8",x"87",x"cb"),
   922 => (x"c5",x"05",x"98",x"70"),
   923 => (x"c0",x"48",x"c0",x"87"),
   924 => (x"da",x"c1",x"87",x"e6"),
   925 => (x"d2",x"02",x"bf",x"e8"),
   926 => (x"c4",x"49",x"73",x"87"),
   927 => (x"e0",x"d2",x"c1",x"91"),
   928 => (x"cf",x"4c",x"69",x"81"),
   929 => (x"ff",x"ff",x"ff",x"ff"),
   930 => (x"73",x"87",x"cb",x"9c"),
   931 => (x"c1",x"91",x"c2",x"49"),
   932 => (x"9f",x"81",x"e0",x"d2"),
   933 => (x"48",x"74",x"4c",x"69"),
   934 => (x"0e",x"87",x"d4",x"ec"),
   935 => (x"5d",x"5c",x"5b",x"5e"),
   936 => (x"c0",x"86",x"f4",x"0e"),
   937 => (x"c1",x"48",x"76",x"4b"),
   938 => (x"78",x"bf",x"fc",x"da"),
   939 => (x"db",x"c1",x"80",x"c4"),
   940 => (x"c1",x"78",x"bf",x"c0"),
   941 => (x"02",x"bf",x"e8",x"da"),
   942 => (x"da",x"c1",x"87",x"c9"),
   943 => (x"c4",x"49",x"bf",x"e0"),
   944 => (x"c1",x"87",x"c7",x"31"),
   945 => (x"49",x"bf",x"c4",x"db"),
   946 => (x"a6",x"cc",x"31",x"c4"),
   947 => (x"c8",x"4d",x"c0",x"59"),
   948 => (x"a8",x"c0",x"48",x"66"),
   949 => (x"87",x"e9",x"c2",x"06"),
   950 => (x"99",x"cf",x"49",x"75"),
   951 => (x"c1",x"87",x"da",x"05"),
   952 => (x"c8",x"1e",x"e0",x"d2"),
   953 => (x"c1",x"48",x"49",x"66"),
   954 => (x"58",x"a6",x"cc",x"80"),
   955 => (x"c0",x"e1",x"1e",x"71"),
   956 => (x"c1",x"86",x"c8",x"87"),
   957 => (x"c3",x"4b",x"e0",x"d2"),
   958 => (x"83",x"e0",x"c0",x"87"),
   959 => (x"71",x"49",x"6b",x"97"),
   960 => (x"f3",x"c1",x"02",x"99"),
   961 => (x"49",x"6b",x"97",x"87"),
   962 => (x"02",x"a9",x"e5",x"c3"),
   963 => (x"cb",x"87",x"e9",x"c1"),
   964 => (x"69",x"97",x"49",x"a3"),
   965 => (x"05",x"99",x"d8",x"49"),
   966 => (x"73",x"87",x"dd",x"c1"),
   967 => (x"f5",x"c4",x"ff",x"1e"),
   968 => (x"cb",x"86",x"c4",x"87"),
   969 => (x"66",x"e4",x"c0",x"1e"),
   970 => (x"e8",x"1e",x"73",x"1e"),
   971 => (x"86",x"cc",x"87",x"f6"),
   972 => (x"c1",x"05",x"98",x"70"),
   973 => (x"a3",x"dc",x"87",x"c2"),
   974 => (x"49",x"66",x"dc",x"4a"),
   975 => (x"79",x"6a",x"81",x"c4"),
   976 => (x"dc",x"4a",x"a3",x"da"),
   977 => (x"81",x"c8",x"49",x"66"),
   978 => (x"70",x"48",x"6a",x"9f"),
   979 => (x"c1",x"4c",x"71",x"79"),
   980 => (x"02",x"bf",x"e8",x"da"),
   981 => (x"a3",x"d4",x"87",x"d0"),
   982 => (x"49",x"69",x"9f",x"49"),
   983 => (x"ff",x"c0",x"4a",x"71"),
   984 => (x"32",x"d0",x"9a",x"ff"),
   985 => (x"4a",x"c0",x"87",x"c2"),
   986 => (x"80",x"6c",x"48",x"72"),
   987 => (x"66",x"dc",x"7c",x"70"),
   988 => (x"c1",x"78",x"c0",x"48"),
   989 => (x"87",x"ff",x"c0",x"48"),
   990 => (x"66",x"c8",x"85",x"c1"),
   991 => (x"d7",x"fd",x"04",x"ad"),
   992 => (x"e8",x"da",x"c1",x"87"),
   993 => (x"ec",x"c0",x"02",x"bf"),
   994 => (x"fa",x"1e",x"6e",x"87"),
   995 => (x"86",x"c4",x"87",x"e2"),
   996 => (x"6e",x"58",x"a6",x"c4"),
   997 => (x"ff",x"ff",x"cf",x"49"),
   998 => (x"a9",x"99",x"f8",x"ff"),
   999 => (x"6e",x"87",x"d6",x"02"),
  1000 => (x"c1",x"89",x"c2",x"49"),
  1001 => (x"91",x"bf",x"e0",x"da"),
  1002 => (x"bf",x"f8",x"da",x"c1"),
  1003 => (x"c8",x"80",x"71",x"48"),
  1004 => (x"d8",x"fc",x"58",x"a6"),
  1005 => (x"f4",x"48",x"c0",x"87"),
  1006 => (x"87",x"f1",x"e7",x"8e"),
  1007 => (x"c8",x"1e",x"73",x"1e"),
  1008 => (x"c1",x"49",x"bf",x"66"),
  1009 => (x"09",x"66",x"c8",x"81"),
  1010 => (x"da",x"c1",x"09",x"79"),
  1011 => (x"05",x"99",x"bf",x"e4"),
  1012 => (x"66",x"c8",x"87",x"d0"),
  1013 => (x"6b",x"83",x"c8",x"4b"),
  1014 => (x"87",x"d4",x"f9",x"1e"),
  1015 => (x"49",x"70",x"86",x"c4"),
  1016 => (x"48",x"c1",x"7b",x"71"),
  1017 => (x"1e",x"87",x"ca",x"e7"),
  1018 => (x"bf",x"f8",x"da",x"c1"),
  1019 => (x"4a",x"66",x"c4",x"49"),
  1020 => (x"4a",x"6a",x"82",x"c8"),
  1021 => (x"da",x"c1",x"8a",x"c2"),
  1022 => (x"72",x"92",x"bf",x"e0"),
  1023 => (x"da",x"c1",x"49",x"a1"),
  1024 => (x"c4",x"4a",x"bf",x"e4"),
  1025 => (x"72",x"9a",x"bf",x"66"),
  1026 => (x"66",x"c8",x"49",x"a1"),
  1027 => (x"ff",x"1e",x"71",x"1e"),
  1028 => (x"c8",x"87",x"de",x"dc"),
  1029 => (x"05",x"98",x"70",x"86"),
  1030 => (x"48",x"c0",x"87",x"c4"),
  1031 => (x"48",x"c1",x"87",x"c2"),
  1032 => (x"0e",x"87",x"d0",x"e6"),
  1033 => (x"0e",x"5c",x"5b",x"5e"),
  1034 => (x"c1",x"1e",x"66",x"cc"),
  1035 => (x"f9",x"1e",x"d8",x"db"),
  1036 => (x"86",x"c8",x"87",x"e9"),
  1037 => (x"c1",x"02",x"98",x"70"),
  1038 => (x"db",x"c1",x"87",x"d2"),
  1039 => (x"c7",x"49",x"bf",x"dc"),
  1040 => (x"29",x"c9",x"81",x"ff"),
  1041 => (x"4b",x"c0",x"4c",x"71"),
  1042 => (x"1e",x"e2",x"c2",x"c1"),
  1043 => (x"87",x"c6",x"c0",x"ff"),
  1044 => (x"b7",x"c0",x"86",x"c4"),
  1045 => (x"c4",x"c1",x"06",x"ac"),
  1046 => (x"1e",x"66",x"d0",x"87"),
  1047 => (x"1e",x"d8",x"db",x"c1"),
  1048 => (x"c8",x"87",x"c4",x"fe"),
  1049 => (x"05",x"98",x"70",x"86"),
  1050 => (x"48",x"c0",x"87",x"c5"),
  1051 => (x"c1",x"87",x"f0",x"c0"),
  1052 => (x"fd",x"1e",x"d8",x"db"),
  1053 => (x"86",x"c4",x"87",x"c6"),
  1054 => (x"c8",x"48",x"66",x"d0"),
  1055 => (x"a6",x"d4",x"80",x"c0"),
  1056 => (x"74",x"83",x"c1",x"58"),
  1057 => (x"ff",x"04",x"ab",x"b7"),
  1058 => (x"87",x"d1",x"87",x"cf"),
  1059 => (x"c1",x"1e",x"66",x"cc"),
  1060 => (x"fe",x"1e",x"fb",x"c2"),
  1061 => (x"c8",x"87",x"f9",x"ff"),
  1062 => (x"c2",x"48",x"c0",x"86"),
  1063 => (x"e4",x"48",x"c1",x"87"),
  1064 => (x"70",x"4f",x"87",x"cd"),
  1065 => (x"64",x"65",x"6e",x"65"),
  1066 => (x"6c",x"69",x"66",x"20"),
  1067 => (x"6c",x"20",x"2c",x"65"),
  1068 => (x"69",x"64",x"61",x"6f"),
  1069 => (x"2e",x"2e",x"67",x"6e"),
  1070 => (x"43",x"00",x"0a",x"2e"),
  1071 => (x"74",x"27",x"6e",x"61"),
  1072 => (x"65",x"70",x"6f",x"20"),
  1073 => (x"73",x"25",x"20",x"6e"),
  1074 => (x"c4",x"1e",x"00",x"0a"),
  1075 => (x"29",x"d8",x"49",x"66"),
  1076 => (x"c4",x"99",x"ff",x"c3"),
  1077 => (x"2a",x"c8",x"4a",x"66"),
  1078 => (x"9a",x"c0",x"fc",x"cf"),
  1079 => (x"66",x"c4",x"b1",x"72"),
  1080 => (x"c0",x"32",x"c8",x"4a"),
  1081 => (x"c0",x"c0",x"f0",x"ff"),
  1082 => (x"c4",x"b1",x"72",x"9a"),
  1083 => (x"32",x"d8",x"4a",x"66"),
  1084 => (x"c0",x"c0",x"c0",x"ff"),
  1085 => (x"b1",x"72",x"9a",x"c0"),
  1086 => (x"87",x"c6",x"48",x"71"),
  1087 => (x"4c",x"26",x"4d",x"26"),
  1088 => (x"4f",x"26",x"4b",x"26"),
  1089 => (x"d0",x"1e",x"73",x"1e"),
  1090 => (x"c0",x"c0",x"c0",x"c0"),
  1091 => (x"fe",x"0f",x"73",x"4b"),
  1092 => (x"26",x"87",x"c4",x"87"),
  1093 => (x"26",x"4c",x"26",x"4d"),
  1094 => (x"1e",x"4f",x"26",x"4b"),
  1095 => (x"c3",x"49",x"66",x"c8"),
  1096 => (x"f7",x"c0",x"99",x"df"),
  1097 => (x"a9",x"b7",x"c0",x"89"),
  1098 => (x"c0",x"87",x"c3",x"03"),
  1099 => (x"66",x"c4",x"81",x"e7"),
  1100 => (x"c8",x"30",x"c4",x"48"),
  1101 => (x"66",x"c4",x"58",x"a6"),
  1102 => (x"c8",x"b0",x"71",x"48"),
  1103 => (x"66",x"c4",x"58",x"a6"),
  1104 => (x"87",x"d5",x"ff",x"48"),
  1105 => (x"5c",x"5b",x"5e",x"0e"),
  1106 => (x"c0",x"c0",x"d0",x"0e"),
  1107 => (x"c1",x"4c",x"c0",x"c0"),
  1108 => (x"48",x"bf",x"e4",x"db"),
  1109 => (x"db",x"c1",x"80",x"c1"),
  1110 => (x"cc",x"97",x"58",x"e8"),
  1111 => (x"c0",x"fe",x"49",x"66"),
  1112 => (x"d3",x"c1",x"b9",x"81"),
  1113 => (x"87",x"db",x"05",x"a9"),
  1114 => (x"48",x"e4",x"db",x"c1"),
  1115 => (x"db",x"c1",x"78",x"c0"),
  1116 => (x"78",x"c0",x"48",x"e8"),
  1117 => (x"48",x"f0",x"db",x"c1"),
  1118 => (x"db",x"c1",x"78",x"c0"),
  1119 => (x"78",x"c0",x"48",x"f4"),
  1120 => (x"c1",x"87",x"fb",x"c6"),
  1121 => (x"48",x"bf",x"e4",x"db"),
  1122 => (x"c0",x"05",x"a8",x"c1"),
  1123 => (x"cc",x"97",x"87",x"f8"),
  1124 => (x"c0",x"fe",x"49",x"66"),
  1125 => (x"1e",x"71",x"b9",x"81"),
  1126 => (x"bf",x"f4",x"db",x"c1"),
  1127 => (x"87",x"fb",x"fd",x"1e"),
  1128 => (x"db",x"c1",x"86",x"c8"),
  1129 => (x"db",x"c1",x"58",x"f8"),
  1130 => (x"c3",x"4a",x"bf",x"f4"),
  1131 => (x"c6",x"06",x"aa",x"b7"),
  1132 => (x"72",x"48",x"ca",x"87"),
  1133 => (x"72",x"4a",x"70",x"88"),
  1134 => (x"71",x"81",x"c1",x"49"),
  1135 => (x"c1",x"30",x"c1",x"48"),
  1136 => (x"c5",x"58",x"f0",x"db"),
  1137 => (x"db",x"c1",x"87",x"f8"),
  1138 => (x"c9",x"48",x"bf",x"f4"),
  1139 => (x"c5",x"01",x"a8",x"b7"),
  1140 => (x"db",x"c1",x"87",x"ec"),
  1141 => (x"c0",x"48",x"bf",x"f4"),
  1142 => (x"c5",x"06",x"a8",x"b7"),
  1143 => (x"db",x"c1",x"87",x"e0"),
  1144 => (x"c3",x"48",x"bf",x"e4"),
  1145 => (x"db",x"01",x"a8",x"b7"),
  1146 => (x"66",x"cc",x"97",x"87"),
  1147 => (x"81",x"c0",x"fe",x"49"),
  1148 => (x"c1",x"1e",x"71",x"b9"),
  1149 => (x"1e",x"bf",x"f0",x"db"),
  1150 => (x"c8",x"87",x"e0",x"fc"),
  1151 => (x"f4",x"db",x"c1",x"86"),
  1152 => (x"87",x"fa",x"c4",x"58"),
  1153 => (x"bf",x"ec",x"db",x"c1"),
  1154 => (x"c1",x"81",x"c3",x"49"),
  1155 => (x"b7",x"bf",x"e4",x"db"),
  1156 => (x"e1",x"c0",x"04",x"a9"),
  1157 => (x"66",x"cc",x"97",x"87"),
  1158 => (x"81",x"c0",x"fe",x"49"),
  1159 => (x"c1",x"1e",x"71",x"b9"),
  1160 => (x"1e",x"bf",x"e8",x"db"),
  1161 => (x"c8",x"87",x"f4",x"fb"),
  1162 => (x"ec",x"db",x"c1",x"86"),
  1163 => (x"f8",x"db",x"c1",x"58"),
  1164 => (x"c4",x"78",x"c1",x"48"),
  1165 => (x"db",x"c1",x"87",x"c8"),
  1166 => (x"c0",x"48",x"bf",x"f4"),
  1167 => (x"c2",x"06",x"a8",x"b7"),
  1168 => (x"db",x"c1",x"87",x"db"),
  1169 => (x"c3",x"48",x"bf",x"f4"),
  1170 => (x"c2",x"01",x"a8",x"b7"),
  1171 => (x"db",x"c1",x"87",x"cf"),
  1172 => (x"c1",x"49",x"bf",x"f0"),
  1173 => (x"db",x"c1",x"81",x"31"),
  1174 => (x"a9",x"b7",x"bf",x"e4"),
  1175 => (x"87",x"df",x"c1",x"04"),
  1176 => (x"49",x"66",x"cc",x"97"),
  1177 => (x"b9",x"81",x"c0",x"fe"),
  1178 => (x"db",x"c1",x"1e",x"71"),
  1179 => (x"fa",x"1e",x"bf",x"fc"),
  1180 => (x"86",x"c8",x"87",x"e9"),
  1181 => (x"58",x"c0",x"dc",x"c1"),
  1182 => (x"bf",x"f8",x"db",x"c1"),
  1183 => (x"c1",x"89",x"c1",x"49"),
  1184 => (x"c0",x"59",x"fc",x"db"),
  1185 => (x"c2",x"03",x"a9",x"b7"),
  1186 => (x"db",x"c1",x"87",x"f4"),
  1187 => (x"c1",x"49",x"bf",x"e8"),
  1188 => (x"bf",x"97",x"fc",x"db"),
  1189 => (x"98",x"ff",x"c3",x"51"),
  1190 => (x"bf",x"e8",x"db",x"c1"),
  1191 => (x"c1",x"81",x"c1",x"49"),
  1192 => (x"c1",x"59",x"ec",x"db"),
  1193 => (x"b7",x"bf",x"c0",x"dc"),
  1194 => (x"c9",x"c0",x"06",x"a9"),
  1195 => (x"c0",x"dc",x"c1",x"87"),
  1196 => (x"e8",x"db",x"c1",x"48"),
  1197 => (x"db",x"c1",x"78",x"bf"),
  1198 => (x"78",x"c1",x"48",x"f8"),
  1199 => (x"c1",x"87",x"ff",x"c1"),
  1200 => (x"05",x"bf",x"f8",x"db"),
  1201 => (x"c1",x"87",x"f7",x"c1"),
  1202 => (x"49",x"bf",x"fc",x"db"),
  1203 => (x"dc",x"c1",x"31",x"c4"),
  1204 => (x"db",x"c1",x"59",x"c0"),
  1205 => (x"97",x"09",x"bf",x"e8"),
  1206 => (x"e1",x"c1",x"09",x"79"),
  1207 => (x"f4",x"db",x"c1",x"87"),
  1208 => (x"b7",x"c7",x"48",x"bf"),
  1209 => (x"d5",x"c1",x"04",x"a8"),
  1210 => (x"fe",x"4b",x"c0",x"87"),
  1211 => (x"78",x"c1",x"48",x"f4"),
  1212 => (x"bf",x"c0",x"dc",x"c1"),
  1213 => (x"c1",x"1e",x"74",x"1e"),
  1214 => (x"fe",x"1e",x"c1",x"cd"),
  1215 => (x"cc",x"87",x"d1",x"f6"),
  1216 => (x"ec",x"db",x"c1",x"86"),
  1217 => (x"e8",x"db",x"c1",x"5c"),
  1218 => (x"dc",x"c1",x"48",x"bf"),
  1219 => (x"a8",x"b7",x"bf",x"c0"),
  1220 => (x"87",x"db",x"c0",x"03"),
  1221 => (x"bf",x"e8",x"db",x"c1"),
  1222 => (x"db",x"c1",x"83",x"bf"),
  1223 => (x"c4",x"49",x"bf",x"e8"),
  1224 => (x"ec",x"db",x"c1",x"81"),
  1225 => (x"c0",x"dc",x"c1",x"59"),
  1226 => (x"04",x"a9",x"b7",x"bf"),
  1227 => (x"73",x"87",x"e5",x"ff"),
  1228 => (x"e0",x"cd",x"c1",x"1e"),
  1229 => (x"d7",x"f5",x"fe",x"1e"),
  1230 => (x"f7",x"86",x"c8",x"87"),
  1231 => (x"d4",x"f7",x"87",x"c6"),
  1232 => (x"65",x"68",x"43",x"87"),
  1233 => (x"75",x"73",x"6b",x"63"),
  1234 => (x"6e",x"69",x"6d",x"6d"),
  1235 => (x"72",x"66",x"20",x"67"),
  1236 => (x"25",x"20",x"6d",x"6f"),
  1237 => (x"6f",x"74",x"20",x"64"),
  1238 => (x"2e",x"64",x"25",x"20"),
  1239 => (x"00",x"20",x"2e",x"2e"),
  1240 => (x"00",x"0a",x"64",x"25"),
  1241 => (x"5c",x"5b",x"5e",x"0e"),
  1242 => (x"d0",x"c1",x"0e",x"5d"),
  1243 => (x"f3",x"fe",x"1e",x"fb"),
  1244 => (x"86",x"c4",x"87",x"e4"),
  1245 => (x"87",x"f9",x"c4",x"ff"),
  1246 => (x"cd",x"02",x"98",x"70"),
  1247 => (x"f4",x"d8",x"ff",x"87"),
  1248 => (x"02",x"98",x"70",x"87"),
  1249 => (x"49",x"c1",x"87",x"c4"),
  1250 => (x"49",x"c0",x"87",x"c2"),
  1251 => (x"d1",x"c1",x"4d",x"71"),
  1252 => (x"f3",x"fe",x"1e",x"d1"),
  1253 => (x"86",x"c4",x"87",x"c0"),
  1254 => (x"48",x"c0",x"dc",x"c1"),
  1255 => (x"ee",x"c0",x"78",x"c0"),
  1256 => (x"d7",x"f2",x"fe",x"1e"),
  1257 => (x"c3",x"86",x"c4",x"87"),
  1258 => (x"4a",x"ff",x"c8",x"f4"),
  1259 => (x"4c",x"bf",x"c0",x"ff"),
  1260 => (x"c0",x"c8",x"49",x"74"),
  1261 => (x"ca",x"c1",x"02",x"99"),
  1262 => (x"c3",x"4b",x"74",x"87"),
  1263 => (x"ab",x"db",x"9b",x"ff"),
  1264 => (x"87",x"f3",x"c0",x"05"),
  1265 => (x"c0",x"02",x"9d",x"75"),
  1266 => (x"c0",x"d0",x"87",x"e3"),
  1267 => (x"1e",x"c0",x"c0",x"c0"),
  1268 => (x"1e",x"df",x"d0",x"c1"),
  1269 => (x"c8",x"87",x"cc",x"f1"),
  1270 => (x"02",x"98",x"70",x"86"),
  1271 => (x"d0",x"c1",x"87",x"cf"),
  1272 => (x"f1",x"fe",x"1e",x"d3"),
  1273 => (x"86",x"c4",x"87",x"f0"),
  1274 => (x"ca",x"87",x"d9",x"f4"),
  1275 => (x"eb",x"d0",x"c1",x"87"),
  1276 => (x"e1",x"f1",x"fe",x"1e"),
  1277 => (x"73",x"86",x"c4",x"87"),
  1278 => (x"87",x"c8",x"f5",x"1e"),
  1279 => (x"f4",x"c3",x"86",x"c4"),
  1280 => (x"72",x"4a",x"c0",x"c9"),
  1281 => (x"71",x"8a",x"c1",x"49"),
  1282 => (x"df",x"fe",x"05",x"99"),
  1283 => (x"87",x"ce",x"fe",x"87"),
  1284 => (x"42",x"87",x"c0",x"f4"),
  1285 => (x"69",x"74",x"6f",x"6f"),
  1286 => (x"2e",x"2e",x"67",x"6e"),
  1287 => (x"42",x"00",x"0a",x"2e"),
  1288 => (x"38",x"54",x"4f",x"4f"),
  1289 => (x"42",x"20",x"32",x"33"),
  1290 => (x"53",x"00",x"4e",x"49"),
  1291 => (x"6f",x"62",x"20",x"44"),
  1292 => (x"66",x"20",x"74",x"6f"),
  1293 => (x"65",x"6c",x"69",x"61"),
  1294 => (x"49",x"00",x"0a",x"64"),
  1295 => (x"69",x"74",x"69",x"6e"),
  1296 => (x"7a",x"69",x"6c",x"61"),
  1297 => (x"20",x"67",x"6e",x"69"),
  1298 => (x"63",x"20",x"44",x"53"),
  1299 => (x"0a",x"64",x"72",x"61"),
  1300 => (x"32",x"53",x"52",x"00"),
  1301 => (x"62",x"20",x"32",x"33"),
  1302 => (x"20",x"74",x"6f",x"6f"),
  1303 => (x"72",x"70",x"20",x"2d"),
  1304 => (x"20",x"73",x"73",x"65"),
  1305 => (x"20",x"43",x"53",x"45"),
  1306 => (x"62",x"20",x"6f",x"74"),
  1307 => (x"20",x"74",x"6f",x"6f"),
  1308 => (x"6d",x"6f",x"72",x"66"),
  1309 => (x"2e",x"44",x"53",x"20"),
  1310 => (x"2e",x"44",x"53",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
