
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"46",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"38"),
    10 => (x"41",x"b0",x"27",x"4f"),
    11 => (x"27",x"4e",x"00",x"00"),
    12 => (x"00",x"00",x"06",x"41"),
    13 => (x"87",x"fd",x"00",x"0f"),
    14 => (x"4e",x"c0",x"f0",x"c1"),
    15 => (x"00",x"00",x"45",x"27"),
    16 => (x"fd",x"00",x"0f",x"00"),
    17 => (x"1e",x"4f",x"4f",x"87"),
    18 => (x"c0",x"ff",x"86",x"fc"),
    19 => (x"c4",x"48",x"69",x"49"),
    20 => (x"a6",x"c4",x"98",x"c0"),
    21 => (x"ff",x"02",x"6e",x"58"),
    22 => (x"66",x"c8",x"87",x"f3"),
    23 => (x"8e",x"fc",x"48",x"79"),
    24 => (x"5e",x"0e",x"4f",x"26"),
    25 => (x"cc",x"0e",x"5c",x"5b"),
    26 => (x"4c",x"c0",x"4b",x"66"),
    27 => (x"9a",x"72",x"4a",x"13"),
    28 => (x"87",x"d9",x"c0",x"02"),
    29 => (x"ff",x"c3",x"49",x"72"),
    30 => (x"27",x"1e",x"71",x"99"),
    31 => (x"00",x"00",x"00",x"47"),
    32 => (x"c1",x"86",x"c4",x"0f"),
    33 => (x"72",x"4a",x"13",x"84"),
    34 => (x"e7",x"ff",x"05",x"9a"),
    35 => (x"26",x"48",x"74",x"87"),
    36 => (x"26",x"4b",x"26",x"4c"),
    37 => (x"5b",x"5e",x"0e",x"4f"),
    38 => (x"d0",x"0e",x"5d",x"5c"),
    39 => (x"f8",x"27",x"4a",x"66"),
    40 => (x"4b",x"00",x"00",x"16"),
    41 => (x"00",x"0f",x"40",x"27"),
    42 => (x"4c",x"c0",x"4d",x"00"),
    43 => (x"c0",x"05",x"9a",x"72"),
    44 => (x"f0",x"c0",x"87",x"c6"),
    45 => (x"87",x"f0",x"c0",x"53"),
    46 => (x"c0",x"02",x"9a",x"72"),
    47 => (x"1e",x"72",x"87",x"ea"),
    48 => (x"66",x"d8",x"49",x"72"),
    49 => (x"05",x"c5",x"27",x"4a"),
    50 => (x"26",x"0f",x"00",x"00"),
    51 => (x"11",x"81",x"75",x"4a"),
    52 => (x"72",x"1e",x"71",x"53"),
    53 => (x"4a",x"66",x"d8",x"49"),
    54 => (x"00",x"05",x"c5",x"27"),
    55 => (x"4a",x"70",x"0f",x"00"),
    56 => (x"9a",x"72",x"49",x"26"),
    57 => (x"87",x"d6",x"ff",x"05"),
    58 => (x"00",x"16",x"f8",x"27"),
    59 => (x"c0",x"02",x"ab",x"00"),
    60 => (x"66",x"d8",x"87",x"e5"),
    61 => (x"1e",x"66",x"dc",x"4d"),
    62 => (x"6b",x"97",x"8b",x"c1"),
    63 => (x"81",x"c0",x"fe",x"49"),
    64 => (x"b9",x"04",x"b1",x"03"),
    65 => (x"75",x"1e",x"71",x"07"),
    66 => (x"c1",x"86",x"c8",x"0f"),
    67 => (x"16",x"f8",x"27",x"84"),
    68 => (x"05",x"ab",x"00",x"00"),
    69 => (x"74",x"87",x"de",x"ff"),
    70 => (x"26",x"4d",x"26",x"48"),
    71 => (x"26",x"4b",x"26",x"4c"),
    72 => (x"5b",x"5e",x"0e",x"4f"),
    73 => (x"d0",x"0e",x"5d",x"5c"),
    74 => (x"4d",x"ff",x"4c",x"66"),
    75 => (x"c0",x"fe",x"4b",x"14"),
    76 => (x"04",x"b3",x"03",x"83"),
    77 => (x"9b",x"73",x"07",x"bb"),
    78 => (x"87",x"e2",x"c0",x"02"),
    79 => (x"66",x"d8",x"85",x"c1"),
    80 => (x"dc",x"1e",x"73",x"1e"),
    81 => (x"86",x"c8",x"0f",x"66"),
    82 => (x"c0",x"05",x"a8",x"73"),
    83 => (x"4b",x"14",x"87",x"d0"),
    84 => (x"03",x"83",x"c0",x"fe"),
    85 => (x"07",x"bb",x"04",x"b3"),
    86 => (x"ff",x"05",x"9b",x"73"),
    87 => (x"48",x"75",x"87",x"de"),
    88 => (x"4c",x"26",x"4d",x"26"),
    89 => (x"4f",x"26",x"4b",x"26"),
    90 => (x"5c",x"5b",x"5e",x"0e"),
    91 => (x"86",x"f4",x"0e",x"5d"),
    92 => (x"4b",x"66",x"e4",x"c0"),
    93 => (x"a6",x"c4",x"4c",x"c0"),
    94 => (x"dc",x"78",x"c0",x"48"),
    95 => (x"4d",x"bf",x"97",x"66"),
    96 => (x"03",x"85",x"c0",x"fe"),
    97 => (x"07",x"bd",x"04",x"b5"),
    98 => (x"c1",x"48",x"66",x"dc"),
    99 => (x"a6",x"e0",x"c0",x"80"),
   100 => (x"02",x"9d",x"75",x"58"),
   101 => (x"c4",x"87",x"c7",x"c5"),
   102 => (x"cc",x"c4",x"02",x"66"),
   103 => (x"48",x"a6",x"c8",x"87"),
   104 => (x"a6",x"c4",x"78",x"c0"),
   105 => (x"75",x"78",x"c0",x"48"),
   106 => (x"ad",x"f0",x"c0",x"49"),
   107 => (x"87",x"e7",x"c1",x"02"),
   108 => (x"02",x"a9",x"e3",x"c1"),
   109 => (x"c1",x"87",x"e8",x"c1"),
   110 => (x"c0",x"02",x"a9",x"e4"),
   111 => (x"ec",x"c1",x"87",x"e6"),
   112 => (x"d2",x"c1",x"02",x"a9"),
   113 => (x"a9",x"f0",x"c1",x"87"),
   114 => (x"87",x"e0",x"c0",x"02"),
   115 => (x"02",x"a9",x"f3",x"c1"),
   116 => (x"c1",x"87",x"e1",x"c0"),
   117 => (x"c0",x"02",x"a9",x"f5"),
   118 => (x"f8",x"c1",x"87",x"ca"),
   119 => (x"cb",x"c0",x"02",x"a9"),
   120 => (x"87",x"da",x"c1",x"87"),
   121 => (x"ca",x"48",x"a6",x"c8"),
   122 => (x"87",x"e9",x"c1",x"78"),
   123 => (x"d0",x"48",x"a6",x"c8"),
   124 => (x"87",x"e1",x"c1",x"78"),
   125 => (x"1e",x"66",x"e8",x"c0"),
   126 => (x"e8",x"c0",x"1e",x"73"),
   127 => (x"80",x"c4",x"48",x"66"),
   128 => (x"58",x"a6",x"ec",x"c0"),
   129 => (x"49",x"66",x"e8",x"c0"),
   130 => (x"1e",x"69",x"89",x"c4"),
   131 => (x"cc",x"87",x"d2",x"fc"),
   132 => (x"84",x"49",x"70",x"86"),
   133 => (x"c4",x"87",x"fe",x"c0"),
   134 => (x"78",x"c1",x"48",x"a6"),
   135 => (x"c0",x"87",x"f6",x"c0"),
   136 => (x"c0",x"1e",x"66",x"e8"),
   137 => (x"c4",x"48",x"66",x"e4"),
   138 => (x"a6",x"e8",x"c0",x"80"),
   139 => (x"66",x"e4",x"c0",x"58"),
   140 => (x"69",x"89",x"c4",x"49"),
   141 => (x"c8",x"0f",x"73",x"1e"),
   142 => (x"c0",x"84",x"c1",x"86"),
   143 => (x"e8",x"c0",x"87",x"d7"),
   144 => (x"e5",x"c0",x"1e",x"66"),
   145 => (x"c8",x"0f",x"73",x"1e"),
   146 => (x"66",x"e8",x"c0",x"86"),
   147 => (x"73",x"1e",x"75",x"1e"),
   148 => (x"c1",x"86",x"c8",x"0f"),
   149 => (x"02",x"66",x"c8",x"84"),
   150 => (x"c0",x"87",x"e7",x"c1"),
   151 => (x"c4",x"48",x"66",x"e0"),
   152 => (x"a6",x"e4",x"c0",x"80"),
   153 => (x"66",x"e0",x"c0",x"58"),
   154 => (x"76",x"89",x"c4",x"49"),
   155 => (x"c1",x"78",x"69",x"48"),
   156 => (x"c0",x"05",x"ad",x"e4"),
   157 => (x"48",x"6e",x"87",x"dc"),
   158 => (x"03",x"a8",x"b7",x"c0"),
   159 => (x"c0",x"87",x"d3",x"c0"),
   160 => (x"47",x"27",x"1e",x"ed"),
   161 => (x"0f",x"00",x"00",x"00"),
   162 => (x"48",x"6e",x"86",x"c4"),
   163 => (x"c4",x"88",x"08",x"c0"),
   164 => (x"e8",x"c0",x"58",x"a6"),
   165 => (x"1e",x"73",x"1e",x"66"),
   166 => (x"cc",x"1e",x"66",x"d0"),
   167 => (x"f4",x"f7",x"1e",x"66"),
   168 => (x"70",x"86",x"d0",x"87"),
   169 => (x"d9",x"c0",x"84",x"49"),
   170 => (x"ad",x"e5",x"c0",x"87"),
   171 => (x"87",x"c8",x"c0",x"05"),
   172 => (x"c1",x"48",x"a6",x"c4"),
   173 => (x"87",x"ca",x"c0",x"78"),
   174 => (x"1e",x"66",x"e8",x"c0"),
   175 => (x"0f",x"73",x"1e",x"75"),
   176 => (x"66",x"dc",x"86",x"c8"),
   177 => (x"fe",x"4d",x"bf",x"97"),
   178 => (x"b5",x"03",x"85",x"c0"),
   179 => (x"dc",x"07",x"bd",x"04"),
   180 => (x"80",x"c1",x"48",x"66"),
   181 => (x"58",x"a6",x"e0",x"c0"),
   182 => (x"fa",x"05",x"9d",x"75"),
   183 => (x"48",x"74",x"87",x"f9"),
   184 => (x"4d",x"26",x"8e",x"f4"),
   185 => (x"4b",x"26",x"4c",x"26"),
   186 => (x"c0",x"1e",x"4f",x"26"),
   187 => (x"00",x"47",x"27",x"1e"),
   188 => (x"d0",x"1e",x"00",x"00"),
   189 => (x"66",x"d0",x"1e",x"66"),
   190 => (x"01",x"68",x"27",x"1e"),
   191 => (x"d0",x"0f",x"00",x"00"),
   192 => (x"1e",x"4f",x"26",x"86"),
   193 => (x"47",x"27",x"1e",x"c0"),
   194 => (x"1e",x"00",x"00",x"00"),
   195 => (x"d0",x"1e",x"a6",x"d0"),
   196 => (x"68",x"27",x"1e",x"66"),
   197 => (x"0f",x"00",x"00",x"01"),
   198 => (x"4f",x"26",x"86",x"d0"),
   199 => (x"4a",x"66",x"c8",x"1e"),
   200 => (x"69",x"81",x"c4",x"49"),
   201 => (x"87",x"da",x"c0",x"02"),
   202 => (x"81",x"c4",x"49",x"72"),
   203 => (x"88",x"c1",x"48",x"69"),
   204 => (x"49",x"6a",x"79",x"70"),
   205 => (x"80",x"c1",x"48",x"71"),
   206 => (x"c4",x"97",x"7a",x"70"),
   207 => (x"c0",x"48",x"51",x"66"),
   208 => (x"48",x"c0",x"87",x"c2"),
   209 => (x"f8",x"1e",x"4f",x"26"),
   210 => (x"cc",x"48",x"76",x"86"),
   211 => (x"a6",x"c4",x"78",x"66"),
   212 => (x"76",x"78",x"ff",x"48"),
   213 => (x"03",x"1c",x"27",x"1e"),
   214 => (x"dc",x"1e",x"00",x"00"),
   215 => (x"66",x"dc",x"1e",x"a6"),
   216 => (x"01",x"68",x"27",x"1e"),
   217 => (x"d0",x"0f",x"00",x"00"),
   218 => (x"26",x"8e",x"f8",x"86"),
   219 => (x"86",x"f8",x"1e",x"4f"),
   220 => (x"66",x"cc",x"48",x"76"),
   221 => (x"48",x"a6",x"c4",x"78"),
   222 => (x"76",x"78",x"66",x"d0"),
   223 => (x"03",x"1c",x"27",x"1e"),
   224 => (x"c0",x"1e",x"00",x"00"),
   225 => (x"c0",x"1e",x"a6",x"e0"),
   226 => (x"27",x"1e",x"66",x"e0"),
   227 => (x"00",x"00",x"01",x"68"),
   228 => (x"f8",x"86",x"d0",x"0f"),
   229 => (x"1e",x"4f",x"26",x"8e"),
   230 => (x"48",x"76",x"86",x"f8"),
   231 => (x"c4",x"78",x"66",x"cc"),
   232 => (x"78",x"ff",x"48",x"a6"),
   233 => (x"1c",x"27",x"1e",x"76"),
   234 => (x"1e",x"00",x"00",x"03"),
   235 => (x"dc",x"1e",x"66",x"dc"),
   236 => (x"68",x"27",x"1e",x"66"),
   237 => (x"0f",x"00",x"00",x"01"),
   238 => (x"8e",x"f8",x"86",x"d0"),
   239 => (x"73",x"1e",x"4f",x"26"),
   240 => (x"4b",x"66",x"cc",x"1e"),
   241 => (x"1e",x"7b",x"66",x"c8"),
   242 => (x"00",x"05",x"b2",x"27"),
   243 => (x"86",x"c4",x"0f",x"00"),
   244 => (x"c0",x"05",x"98",x"70"),
   245 => (x"7b",x"c3",x"87",x"c2"),
   246 => (x"48",x"49",x"66",x"c8"),
   247 => (x"c0",x"02",x"a8",x"c0"),
   248 => (x"a9",x"c1",x"87",x"db"),
   249 => (x"87",x"da",x"c0",x"02"),
   250 => (x"c0",x"02",x"a9",x"c2"),
   251 => (x"a9",x"c3",x"87",x"ed"),
   252 => (x"87",x"ee",x"c0",x"02"),
   253 => (x"c0",x"02",x"a9",x"c4"),
   254 => (x"e5",x"c0",x"87",x"e6"),
   255 => (x"c0",x"7b",x"c0",x"87"),
   256 => (x"10",x"27",x"87",x"e0"),
   257 => (x"bf",x"00",x"00",x"17"),
   258 => (x"b7",x"e4",x"c1",x"48"),
   259 => (x"c5",x"c0",x"06",x"a8"),
   260 => (x"c0",x"7b",x"c0",x"87"),
   261 => (x"7b",x"c3",x"87",x"cc"),
   262 => (x"c1",x"87",x"c7",x"c0"),
   263 => (x"87",x"c2",x"c0",x"7b"),
   264 => (x"4b",x"26",x"7b",x"c2"),
   265 => (x"c4",x"1e",x"4f",x"26"),
   266 => (x"81",x"c2",x"49",x"66"),
   267 => (x"71",x"48",x"66",x"c8"),
   268 => (x"08",x"66",x"cc",x"80"),
   269 => (x"4f",x"26",x"08",x"78"),
   270 => (x"5c",x"5b",x"5e",x"0e"),
   271 => (x"66",x"d8",x"0e",x"5d"),
   272 => (x"74",x"84",x"c5",x"4c"),
   273 => (x"d0",x"93",x"c4",x"4b"),
   274 => (x"66",x"dc",x"83",x"66"),
   275 => (x"c1",x"49",x"74",x"7b"),
   276 => (x"c4",x"4a",x"71",x"81"),
   277 => (x"82",x"66",x"d0",x"92"),
   278 => (x"4a",x"74",x"7a",x"6b"),
   279 => (x"92",x"c4",x"82",x"de"),
   280 => (x"74",x"82",x"66",x"d0"),
   281 => (x"b7",x"71",x"4d",x"7a"),
   282 => (x"dd",x"c0",x"01",x"ac"),
   283 => (x"c3",x"4a",x"74",x"87"),
   284 => (x"66",x"d4",x"92",x"c8"),
   285 => (x"c4",x"49",x"75",x"82"),
   286 => (x"74",x"81",x"72",x"91"),
   287 => (x"74",x"85",x"c1",x"79"),
   288 => (x"71",x"81",x"c1",x"49"),
   289 => (x"ff",x"06",x"ad",x"b7"),
   290 => (x"4a",x"74",x"87",x"e3"),
   291 => (x"d4",x"92",x"c8",x"c3"),
   292 => (x"49",x"74",x"82",x"66"),
   293 => (x"91",x"c4",x"89",x"c1"),
   294 => (x"48",x"69",x"81",x"72"),
   295 => (x"79",x"70",x"80",x"c1"),
   296 => (x"91",x"c4",x"49",x"74"),
   297 => (x"71",x"4a",x"66",x"d0"),
   298 => (x"d4",x"4b",x"74",x"82"),
   299 => (x"93",x"c8",x"c3",x"83"),
   300 => (x"73",x"83",x"66",x"d4"),
   301 => (x"27",x"79",x"6a",x"81"),
   302 => (x"00",x"00",x"17",x"10"),
   303 => (x"26",x"78",x"c5",x"48"),
   304 => (x"26",x"4c",x"26",x"4d"),
   305 => (x"0e",x"4f",x"26",x"4b"),
   306 => (x"97",x"0e",x"5b",x"5e"),
   307 => (x"73",x"4b",x"66",x"c8"),
   308 => (x"82",x"c0",x"fe",x"4a"),
   309 => (x"ba",x"04",x"b2",x"03"),
   310 => (x"66",x"cc",x"97",x"07"),
   311 => (x"81",x"c0",x"fe",x"49"),
   312 => (x"b9",x"04",x"b1",x"03"),
   313 => (x"aa",x"b7",x"71",x"07"),
   314 => (x"87",x"c5",x"c0",x"02"),
   315 => (x"c9",x"c0",x"48",x"c0"),
   316 => (x"17",x"1c",x"27",x"87"),
   317 => (x"5b",x"97",x"00",x"00"),
   318 => (x"4b",x"26",x"48",x"c1"),
   319 => (x"5e",x"0e",x"4f",x"26"),
   320 => (x"fc",x"0e",x"5c",x"5b"),
   321 => (x"4c",x"6e",x"97",x"86"),
   322 => (x"66",x"d4",x"4b",x"c2"),
   323 => (x"73",x"81",x"c1",x"49"),
   324 => (x"49",x"69",x"97",x"81"),
   325 => (x"03",x"81",x"c0",x"fe"),
   326 => (x"07",x"b9",x"04",x"b1"),
   327 => (x"66",x"d4",x"1e",x"71"),
   328 => (x"97",x"81",x"73",x"49"),
   329 => (x"c0",x"fe",x"49",x"69"),
   330 => (x"04",x"b1",x"03",x"81"),
   331 => (x"1e",x"71",x"07",x"b9"),
   332 => (x"00",x"04",x"c7",x"27"),
   333 => (x"86",x"c8",x"0f",x"00"),
   334 => (x"c0",x"05",x"98",x"70"),
   335 => (x"c1",x"c1",x"87",x"c5"),
   336 => (x"c2",x"83",x"c1",x"4c"),
   337 => (x"ff",x"06",x"ab",x"b7"),
   338 => (x"49",x"74",x"87",x"c0"),
   339 => (x"03",x"81",x"c0",x"fe"),
   340 => (x"07",x"b9",x"04",x"b1"),
   341 => (x"a9",x"b7",x"d7",x"c1"),
   342 => (x"87",x"d4",x"c0",x"04"),
   343 => (x"c0",x"fe",x"49",x"74"),
   344 => (x"04",x"b1",x"03",x"81"),
   345 => (x"da",x"c1",x"07",x"b9"),
   346 => (x"c0",x"03",x"a9",x"b7"),
   347 => (x"4b",x"c7",x"87",x"c2"),
   348 => (x"c0",x"fe",x"49",x"74"),
   349 => (x"04",x"b1",x"03",x"81"),
   350 => (x"d2",x"c1",x"07",x"b9"),
   351 => (x"c5",x"c0",x"05",x"a9"),
   352 => (x"c0",x"48",x"c1",x"87"),
   353 => (x"66",x"d0",x"87",x"e4"),
   354 => (x"49",x"66",x"d4",x"4a"),
   355 => (x"00",x"06",x"29",x"27"),
   356 => (x"b7",x"c0",x"0f",x"00"),
   357 => (x"cf",x"c0",x"06",x"a8"),
   358 => (x"c7",x"48",x"73",x"87"),
   359 => (x"17",x"14",x"27",x"80"),
   360 => (x"c1",x"58",x"00",x"00"),
   361 => (x"87",x"c2",x"c0",x"48"),
   362 => (x"8e",x"fc",x"48",x"c0"),
   363 => (x"4b",x"26",x"4c",x"26"),
   364 => (x"c4",x"1e",x"4f",x"26"),
   365 => (x"a8",x"c2",x"48",x"66"),
   366 => (x"87",x"c5",x"c0",x"05"),
   367 => (x"c2",x"c0",x"48",x"c1"),
   368 => (x"26",x"48",x"c0",x"87"),
   369 => (x"1e",x"73",x"1e",x"4f"),
   370 => (x"e7",x"02",x"9a",x"72"),
   371 => (x"c1",x"48",x"c0",x"87"),
   372 => (x"06",x"a9",x"72",x"4b"),
   373 => (x"82",x"72",x"87",x"d1"),
   374 => (x"73",x"87",x"c9",x"06"),
   375 => (x"01",x"a9",x"72",x"83"),
   376 => (x"87",x"c3",x"87",x"f4"),
   377 => (x"72",x"3a",x"b2",x"c1"),
   378 => (x"73",x"89",x"03",x"a9"),
   379 => (x"2a",x"c1",x"07",x"80"),
   380 => (x"87",x"f3",x"05",x"2b"),
   381 => (x"4f",x"26",x"4b",x"26"),
   382 => (x"c4",x"1e",x"75",x"1e"),
   383 => (x"a1",x"b7",x"71",x"4d"),
   384 => (x"c1",x"b9",x"ff",x"04"),
   385 => (x"07",x"bd",x"c3",x"81"),
   386 => (x"04",x"a2",x"b7",x"72"),
   387 => (x"82",x"c1",x"ba",x"ff"),
   388 => (x"fe",x"07",x"bd",x"c1"),
   389 => (x"2d",x"c1",x"87",x"ef"),
   390 => (x"c1",x"b8",x"ff",x"04"),
   391 => (x"04",x"2d",x"07",x"80"),
   392 => (x"81",x"c1",x"b9",x"ff"),
   393 => (x"26",x"4d",x"26",x"07"),
   394 => (x"1e",x"72",x"1e",x"4f"),
   395 => (x"02",x"11",x"48",x"12"),
   396 => (x"02",x"88",x"87",x"c4"),
   397 => (x"4a",x"26",x"87",x"f6"),
   398 => (x"ff",x"1e",x"4f",x"26"),
   399 => (x"26",x"48",x"bf",x"c8"),
   400 => (x"5b",x"5e",x"0e",x"4f"),
   401 => (x"f0",x"0e",x"5d",x"5c"),
   402 => (x"4b",x"66",x"c4",x"86"),
   403 => (x"00",x"17",x"0c",x"27"),
   404 => (x"10",x"27",x"48",x"00"),
   405 => (x"78",x"00",x"00",x"3f"),
   406 => (x"00",x"17",x"08",x"27"),
   407 => (x"40",x"27",x"48",x"00"),
   408 => (x"78",x"00",x"00",x"3f"),
   409 => (x"00",x"3f",x"40",x"27"),
   410 => (x"10",x"27",x"48",x"00"),
   411 => (x"78",x"00",x"00",x"3f"),
   412 => (x"00",x"3f",x"44",x"27"),
   413 => (x"78",x"c0",x"48",x"00"),
   414 => (x"00",x"3f",x"48",x"27"),
   415 => (x"78",x"c2",x"48",x"00"),
   416 => (x"00",x"3f",x"4c",x"27"),
   417 => (x"e8",x"c0",x"48",x"00"),
   418 => (x"3f",x"50",x"27",x"78"),
   419 => (x"27",x"4a",x"00",x"00"),
   420 => (x"00",x"00",x"10",x"ca"),
   421 => (x"20",x"42",x"20",x"48"),
   422 => (x"20",x"42",x"20",x"42"),
   423 => (x"20",x"42",x"20",x"42"),
   424 => (x"10",x"42",x"20",x"42"),
   425 => (x"10",x"52",x"10",x"52"),
   426 => (x"3f",x"70",x"27",x"52"),
   427 => (x"27",x"4a",x"00",x"00"),
   428 => (x"00",x"00",x"10",x"e9"),
   429 => (x"20",x"42",x"20",x"48"),
   430 => (x"20",x"42",x"20",x"42"),
   431 => (x"20",x"42",x"20",x"42"),
   432 => (x"10",x"42",x"20",x"42"),
   433 => (x"10",x"52",x"10",x"52"),
   434 => (x"1e",x"44",x"27",x"52"),
   435 => (x"ca",x"48",x"00",x"00"),
   436 => (x"11",x"08",x"27",x"78"),
   437 => (x"27",x"1e",x"00",x"00"),
   438 => (x"00",x"00",x"03",x"03"),
   439 => (x"27",x"86",x"c4",x"0f"),
   440 => (x"00",x"00",x"11",x"0a"),
   441 => (x"03",x"03",x"27",x"1e"),
   442 => (x"c4",x"0f",x"00",x"00"),
   443 => (x"11",x"3a",x"27",x"86"),
   444 => (x"27",x"1e",x"00",x"00"),
   445 => (x"00",x"00",x"03",x"03"),
   446 => (x"27",x"86",x"c4",x"0f"),
   447 => (x"00",x"00",x"16",x"f0"),
   448 => (x"df",x"c0",x"02",x"bf"),
   449 => (x"0f",x"51",x"27",x"87"),
   450 => (x"27",x"1e",x"00",x"00"),
   451 => (x"00",x"00",x"03",x"03"),
   452 => (x"27",x"86",x"c4",x"0f"),
   453 => (x"00",x"00",x"0f",x"7d"),
   454 => (x"03",x"03",x"27",x"1e"),
   455 => (x"c4",x"0f",x"00",x"00"),
   456 => (x"87",x"dc",x"c0",x"86"),
   457 => (x"00",x"0f",x"7f",x"27"),
   458 => (x"03",x"27",x"1e",x"00"),
   459 => (x"0f",x"00",x"00",x"03"),
   460 => (x"ae",x"27",x"86",x"c4"),
   461 => (x"1e",x"00",x"00",x"0f"),
   462 => (x"00",x"03",x"03",x"27"),
   463 => (x"86",x"c4",x"0f",x"00"),
   464 => (x"00",x"16",x"f4",x"27"),
   465 => (x"27",x"1e",x"bf",x"00"),
   466 => (x"00",x"00",x"11",x"3c"),
   467 => (x"03",x"03",x"27",x"1e"),
   468 => (x"c8",x"0f",x"00",x"00"),
   469 => (x"06",x"3a",x"27",x"86"),
   470 => (x"27",x"0f",x"00",x"00"),
   471 => (x"00",x"00",x"3e",x"fc"),
   472 => (x"27",x"4c",x"c1",x"58"),
   473 => (x"00",x"00",x"16",x"f4"),
   474 => (x"b7",x"c0",x"48",x"bf"),
   475 => (x"c3",x"c6",x"06",x"a8"),
   476 => (x"0f",x"2c",x"27",x"87"),
   477 => (x"27",x"0f",x"00",x"00"),
   478 => (x"00",x"00",x"0e",x"f3"),
   479 => (x"c2",x"48",x"76",x"0f"),
   480 => (x"27",x"4b",x"c3",x"78"),
   481 => (x"00",x"00",x"3f",x"90"),
   482 => (x"0f",x"cf",x"27",x"4a"),
   483 => (x"20",x"48",x"00",x"00"),
   484 => (x"20",x"42",x"20",x"42"),
   485 => (x"20",x"42",x"20",x"42"),
   486 => (x"20",x"42",x"20",x"42"),
   487 => (x"10",x"52",x"10",x"42"),
   488 => (x"c8",x"52",x"10",x"52"),
   489 => (x"78",x"c1",x"48",x"a6"),
   490 => (x"00",x"3f",x"90",x"27"),
   491 => (x"70",x"27",x"1e",x"00"),
   492 => (x"1e",x"00",x"00",x"3f"),
   493 => (x"00",x"04",x"fe",x"27"),
   494 => (x"86",x"c8",x"0f",x"00"),
   495 => (x"c0",x"05",x"98",x"70"),
   496 => (x"49",x"c1",x"87",x"c5"),
   497 => (x"c0",x"87",x"c2",x"c0"),
   498 => (x"17",x"18",x"27",x"49"),
   499 => (x"6e",x"59",x"00",x"00"),
   500 => (x"c0",x"06",x"ab",x"b7"),
   501 => (x"49",x"6e",x"87",x"e9"),
   502 => (x"48",x"71",x"91",x"c5"),
   503 => (x"a6",x"d0",x"88",x"73"),
   504 => (x"1e",x"a6",x"cc",x"58"),
   505 => (x"66",x"c8",x"1e",x"73"),
   506 => (x"04",x"26",x"27",x"1e"),
   507 => (x"cc",x"0f",x"00",x"00"),
   508 => (x"c1",x"48",x"6e",x"86"),
   509 => (x"58",x"a6",x"c4",x"80"),
   510 => (x"01",x"ab",x"b7",x"6e"),
   511 => (x"cc",x"87",x"d7",x"ff"),
   512 => (x"66",x"c4",x"1e",x"66"),
   513 => (x"17",x"e8",x"27",x"1e"),
   514 => (x"27",x"1e",x"00",x"00"),
   515 => (x"00",x"00",x"17",x"20"),
   516 => (x"04",x"38",x"27",x"1e"),
   517 => (x"d0",x"0f",x"00",x"00"),
   518 => (x"17",x"08",x"27",x"86"),
   519 => (x"1e",x"bf",x"00",x"00"),
   520 => (x"00",x"0d",x"e0",x"27"),
   521 => (x"86",x"c4",x"0f",x"00"),
   522 => (x"27",x"4d",x"c1",x"c1"),
   523 => (x"00",x"00",x"17",x"19"),
   524 => (x"fe",x"49",x"bf",x"97"),
   525 => (x"b1",x"03",x"81",x"c0"),
   526 => (x"c1",x"07",x"b9",x"04"),
   527 => (x"04",x"a9",x"b7",x"c1"),
   528 => (x"c1",x"87",x"f6",x"c1"),
   529 => (x"49",x"75",x"1e",x"c3"),
   530 => (x"03",x"81",x"c0",x"fe"),
   531 => (x"07",x"b9",x"04",x"b1"),
   532 => (x"c7",x"27",x"1e",x"71"),
   533 => (x"0f",x"00",x"00",x"04"),
   534 => (x"66",x"c8",x"86",x"c8"),
   535 => (x"f5",x"c0",x"05",x"a8"),
   536 => (x"1e",x"a6",x"c8",x"87"),
   537 => (x"be",x"27",x"1e",x"c0"),
   538 => (x"0f",x"00",x"00",x"03"),
   539 => (x"90",x"27",x"86",x"c8"),
   540 => (x"4a",x"00",x"00",x"3f"),
   541 => (x"00",x"0f",x"b0",x"27"),
   542 => (x"42",x"20",x"48",x"00"),
   543 => (x"42",x"20",x"42",x"20"),
   544 => (x"42",x"20",x"42",x"20"),
   545 => (x"42",x"20",x"42",x"20"),
   546 => (x"52",x"10",x"52",x"10"),
   547 => (x"4b",x"74",x"52",x"10"),
   548 => (x"00",x"17",x"14",x"27"),
   549 => (x"85",x"c1",x"5c",x"00"),
   550 => (x"c0",x"fe",x"4a",x"75"),
   551 => (x"04",x"b2",x"03",x"82"),
   552 => (x"19",x"27",x"07",x"ba"),
   553 => (x"97",x"00",x"00",x"17"),
   554 => (x"c0",x"fe",x"49",x"bf"),
   555 => (x"04",x"b1",x"03",x"81"),
   556 => (x"b7",x"71",x"07",x"b9"),
   557 => (x"ca",x"fe",x"06",x"aa"),
   558 => (x"71",x"93",x"6e",x"87"),
   559 => (x"73",x"1e",x"72",x"1e"),
   560 => (x"4a",x"66",x"d4",x"49"),
   561 => (x"00",x"05",x"f8",x"27"),
   562 => (x"4a",x"26",x"0f",x"00"),
   563 => (x"a6",x"c4",x"49",x"26"),
   564 => (x"cc",x"49",x"73",x"58"),
   565 => (x"91",x"c7",x"89",x"66"),
   566 => (x"8b",x"6e",x"4b",x"71"),
   567 => (x"6f",x"27",x"1e",x"76"),
   568 => (x"0f",x"00",x"00",x"0e"),
   569 => (x"84",x"c1",x"86",x"c4"),
   570 => (x"00",x"16",x"f4",x"27"),
   571 => (x"ac",x"b7",x"bf",x"00"),
   572 => (x"87",x"fd",x"f9",x"06"),
   573 => (x"00",x"06",x"3a",x"27"),
   574 => (x"00",x"27",x"0f",x"00"),
   575 => (x"58",x"00",x"00",x"3f"),
   576 => (x"00",x"11",x"69",x"27"),
   577 => (x"03",x"27",x"1e",x"00"),
   578 => (x"0f",x"00",x"00",x"03"),
   579 => (x"79",x"27",x"86",x"c4"),
   580 => (x"1e",x"00",x"00",x"11"),
   581 => (x"00",x"03",x"03",x"27"),
   582 => (x"86",x"c4",x"0f",x"00"),
   583 => (x"00",x"11",x"7b",x"27"),
   584 => (x"03",x"27",x"1e",x"00"),
   585 => (x"0f",x"00",x"00",x"03"),
   586 => (x"b1",x"27",x"86",x"c4"),
   587 => (x"1e",x"00",x"00",x"11"),
   588 => (x"00",x"03",x"03",x"27"),
   589 => (x"86",x"c4",x"0f",x"00"),
   590 => (x"00",x"17",x"10",x"27"),
   591 => (x"27",x"1e",x"bf",x"00"),
   592 => (x"00",x"00",x"11",x"b3"),
   593 => (x"03",x"03",x"27",x"1e"),
   594 => (x"c8",x"0f",x"00",x"00"),
   595 => (x"27",x"1e",x"c5",x"86"),
   596 => (x"00",x"00",x"11",x"cc"),
   597 => (x"03",x"03",x"27",x"1e"),
   598 => (x"c8",x"0f",x"00",x"00"),
   599 => (x"17",x"14",x"27",x"86"),
   600 => (x"1e",x"bf",x"00",x"00"),
   601 => (x"00",x"11",x"e5",x"27"),
   602 => (x"03",x"27",x"1e",x"00"),
   603 => (x"0f",x"00",x"00",x"03"),
   604 => (x"1e",x"c1",x"86",x"c8"),
   605 => (x"00",x"11",x"fe",x"27"),
   606 => (x"03",x"27",x"1e",x"00"),
   607 => (x"0f",x"00",x"00",x"03"),
   608 => (x"18",x"27",x"86",x"c8"),
   609 => (x"97",x"00",x"00",x"17"),
   610 => (x"c0",x"fe",x"49",x"bf"),
   611 => (x"04",x"b1",x"03",x"81"),
   612 => (x"1e",x"71",x"07",x"b9"),
   613 => (x"00",x"12",x"17",x"27"),
   614 => (x"03",x"27",x"1e",x"00"),
   615 => (x"0f",x"00",x"00",x"03"),
   616 => (x"c1",x"c1",x"86",x"c8"),
   617 => (x"12",x"30",x"27",x"1e"),
   618 => (x"27",x"1e",x"00",x"00"),
   619 => (x"00",x"00",x"03",x"03"),
   620 => (x"27",x"86",x"c8",x"0f"),
   621 => (x"00",x"00",x"17",x"19"),
   622 => (x"fe",x"49",x"bf",x"97"),
   623 => (x"b1",x"03",x"81",x"c0"),
   624 => (x"71",x"07",x"b9",x"04"),
   625 => (x"12",x"49",x"27",x"1e"),
   626 => (x"27",x"1e",x"00",x"00"),
   627 => (x"00",x"00",x"03",x"03"),
   628 => (x"c1",x"86",x"c8",x"0f"),
   629 => (x"62",x"27",x"1e",x"c2"),
   630 => (x"1e",x"00",x"00",x"12"),
   631 => (x"00",x"03",x"03",x"27"),
   632 => (x"86",x"c8",x"0f",x"00"),
   633 => (x"00",x"17",x"40",x"27"),
   634 => (x"27",x"1e",x"bf",x"00"),
   635 => (x"00",x"00",x"12",x"7b"),
   636 => (x"03",x"03",x"27",x"1e"),
   637 => (x"c8",x"0f",x"00",x"00"),
   638 => (x"27",x"1e",x"c7",x"86"),
   639 => (x"00",x"00",x"12",x"94"),
   640 => (x"03",x"03",x"27",x"1e"),
   641 => (x"c8",x"0f",x"00",x"00"),
   642 => (x"1e",x"44",x"27",x"86"),
   643 => (x"1e",x"bf",x"00",x"00"),
   644 => (x"00",x"12",x"ad",x"27"),
   645 => (x"03",x"27",x"1e",x"00"),
   646 => (x"0f",x"00",x"00",x"03"),
   647 => (x"c6",x"27",x"86",x"c8"),
   648 => (x"1e",x"00",x"00",x"12"),
   649 => (x"00",x"03",x"03",x"27"),
   650 => (x"86",x"c4",x"0f",x"00"),
   651 => (x"00",x"12",x"f0",x"27"),
   652 => (x"03",x"27",x"1e",x"00"),
   653 => (x"0f",x"00",x"00",x"03"),
   654 => (x"08",x"27",x"86",x"c4"),
   655 => (x"bf",x"00",x"00",x"17"),
   656 => (x"fc",x"27",x"1e",x"bf"),
   657 => (x"1e",x"00",x"00",x"12"),
   658 => (x"00",x"03",x"03",x"27"),
   659 => (x"86",x"c8",x"0f",x"00"),
   660 => (x"00",x"13",x"15",x"27"),
   661 => (x"03",x"27",x"1e",x"00"),
   662 => (x"0f",x"00",x"00",x"03"),
   663 => (x"08",x"27",x"86",x"c4"),
   664 => (x"bf",x"00",x"00",x"17"),
   665 => (x"69",x"81",x"c4",x"49"),
   666 => (x"13",x"46",x"27",x"1e"),
   667 => (x"27",x"1e",x"00",x"00"),
   668 => (x"00",x"00",x"03",x"03"),
   669 => (x"c0",x"86",x"c8",x"0f"),
   670 => (x"13",x"5f",x"27",x"1e"),
   671 => (x"27",x"1e",x"00",x"00"),
   672 => (x"00",x"00",x"03",x"03"),
   673 => (x"27",x"86",x"c8",x"0f"),
   674 => (x"00",x"00",x"17",x"08"),
   675 => (x"81",x"c8",x"49",x"bf"),
   676 => (x"78",x"27",x"1e",x"69"),
   677 => (x"1e",x"00",x"00",x"13"),
   678 => (x"00",x"03",x"03",x"27"),
   679 => (x"86",x"c8",x"0f",x"00"),
   680 => (x"91",x"27",x"1e",x"c2"),
   681 => (x"1e",x"00",x"00",x"13"),
   682 => (x"00",x"03",x"03",x"27"),
   683 => (x"86",x"c8",x"0f",x"00"),
   684 => (x"00",x"17",x"08",x"27"),
   685 => (x"cc",x"49",x"bf",x"00"),
   686 => (x"27",x"1e",x"69",x"81"),
   687 => (x"00",x"00",x"13",x"aa"),
   688 => (x"03",x"03",x"27",x"1e"),
   689 => (x"c8",x"0f",x"00",x"00"),
   690 => (x"27",x"1e",x"d1",x"86"),
   691 => (x"00",x"00",x"13",x"c3"),
   692 => (x"03",x"03",x"27",x"1e"),
   693 => (x"c8",x"0f",x"00",x"00"),
   694 => (x"17",x"08",x"27",x"86"),
   695 => (x"49",x"bf",x"00",x"00"),
   696 => (x"1e",x"71",x"81",x"d0"),
   697 => (x"00",x"13",x"dc",x"27"),
   698 => (x"03",x"27",x"1e",x"00"),
   699 => (x"0f",x"00",x"00",x"03"),
   700 => (x"f5",x"27",x"86",x"c8"),
   701 => (x"1e",x"00",x"00",x"13"),
   702 => (x"00",x"03",x"03",x"27"),
   703 => (x"86",x"c4",x"0f",x"00"),
   704 => (x"00",x"14",x"2a",x"27"),
   705 => (x"03",x"27",x"1e",x"00"),
   706 => (x"0f",x"00",x"00",x"03"),
   707 => (x"0c",x"27",x"86",x"c4"),
   708 => (x"bf",x"00",x"00",x"17"),
   709 => (x"3b",x"27",x"1e",x"bf"),
   710 => (x"1e",x"00",x"00",x"14"),
   711 => (x"00",x"03",x"03",x"27"),
   712 => (x"86",x"c8",x"0f",x"00"),
   713 => (x"00",x"14",x"54",x"27"),
   714 => (x"03",x"27",x"1e",x"00"),
   715 => (x"0f",x"00",x"00",x"03"),
   716 => (x"0c",x"27",x"86",x"c4"),
   717 => (x"bf",x"00",x"00",x"17"),
   718 => (x"69",x"81",x"c4",x"49"),
   719 => (x"14",x"94",x"27",x"1e"),
   720 => (x"27",x"1e",x"00",x"00"),
   721 => (x"00",x"00",x"03",x"03"),
   722 => (x"c0",x"86",x"c8",x"0f"),
   723 => (x"14",x"ad",x"27",x"1e"),
   724 => (x"27",x"1e",x"00",x"00"),
   725 => (x"00",x"00",x"03",x"03"),
   726 => (x"27",x"86",x"c8",x"0f"),
   727 => (x"00",x"00",x"17",x"0c"),
   728 => (x"81",x"c8",x"49",x"bf"),
   729 => (x"c6",x"27",x"1e",x"69"),
   730 => (x"1e",x"00",x"00",x"14"),
   731 => (x"00",x"03",x"03",x"27"),
   732 => (x"86",x"c8",x"0f",x"00"),
   733 => (x"df",x"27",x"1e",x"c1"),
   734 => (x"1e",x"00",x"00",x"14"),
   735 => (x"00",x"03",x"03",x"27"),
   736 => (x"86",x"c8",x"0f",x"00"),
   737 => (x"00",x"17",x"0c",x"27"),
   738 => (x"cc",x"49",x"bf",x"00"),
   739 => (x"27",x"1e",x"69",x"81"),
   740 => (x"00",x"00",x"14",x"f8"),
   741 => (x"03",x"03",x"27",x"1e"),
   742 => (x"c8",x"0f",x"00",x"00"),
   743 => (x"27",x"1e",x"d2",x"86"),
   744 => (x"00",x"00",x"15",x"11"),
   745 => (x"03",x"03",x"27",x"1e"),
   746 => (x"c8",x"0f",x"00",x"00"),
   747 => (x"17",x"0c",x"27",x"86"),
   748 => (x"49",x"bf",x"00",x"00"),
   749 => (x"1e",x"71",x"81",x"d0"),
   750 => (x"00",x"15",x"2a",x"27"),
   751 => (x"03",x"27",x"1e",x"00"),
   752 => (x"0f",x"00",x"00",x"03"),
   753 => (x"43",x"27",x"86",x"c8"),
   754 => (x"1e",x"00",x"00",x"15"),
   755 => (x"00",x"03",x"03",x"27"),
   756 => (x"86",x"c4",x"0f",x"00"),
   757 => (x"78",x"27",x"1e",x"6e"),
   758 => (x"1e",x"00",x"00",x"15"),
   759 => (x"00",x"03",x"03",x"27"),
   760 => (x"86",x"c8",x"0f",x"00"),
   761 => (x"91",x"27",x"1e",x"c5"),
   762 => (x"1e",x"00",x"00",x"15"),
   763 => (x"00",x"03",x"03",x"27"),
   764 => (x"86",x"c8",x"0f",x"00"),
   765 => (x"aa",x"27",x"1e",x"73"),
   766 => (x"1e",x"00",x"00",x"15"),
   767 => (x"00",x"03",x"03",x"27"),
   768 => (x"86",x"c8",x"0f",x"00"),
   769 => (x"c3",x"27",x"1e",x"cd"),
   770 => (x"1e",x"00",x"00",x"15"),
   771 => (x"00",x"03",x"03",x"27"),
   772 => (x"86",x"c8",x"0f",x"00"),
   773 => (x"27",x"1e",x"66",x"cc"),
   774 => (x"00",x"00",x"15",x"dc"),
   775 => (x"03",x"03",x"27",x"1e"),
   776 => (x"c8",x"0f",x"00",x"00"),
   777 => (x"27",x"1e",x"c7",x"86"),
   778 => (x"00",x"00",x"15",x"f5"),
   779 => (x"03",x"03",x"27",x"1e"),
   780 => (x"c8",x"0f",x"00",x"00"),
   781 => (x"1e",x"66",x"c8",x"86"),
   782 => (x"00",x"16",x"0e",x"27"),
   783 => (x"03",x"27",x"1e",x"00"),
   784 => (x"0f",x"00",x"00",x"03"),
   785 => (x"1e",x"c1",x"86",x"c8"),
   786 => (x"00",x"16",x"27",x"27"),
   787 => (x"03",x"27",x"1e",x"00"),
   788 => (x"0f",x"00",x"00",x"03"),
   789 => (x"70",x"27",x"86",x"c8"),
   790 => (x"1e",x"00",x"00",x"3f"),
   791 => (x"00",x"16",x"40",x"27"),
   792 => (x"03",x"27",x"1e",x"00"),
   793 => (x"0f",x"00",x"00",x"03"),
   794 => (x"59",x"27",x"86",x"c8"),
   795 => (x"1e",x"00",x"00",x"16"),
   796 => (x"00",x"03",x"03",x"27"),
   797 => (x"86",x"c4",x"0f",x"00"),
   798 => (x"00",x"3f",x"90",x"27"),
   799 => (x"8e",x"27",x"1e",x"00"),
   800 => (x"1e",x"00",x"00",x"16"),
   801 => (x"00",x"03",x"03",x"27"),
   802 => (x"86",x"c8",x"0f",x"00"),
   803 => (x"00",x"16",x"a7",x"27"),
   804 => (x"03",x"27",x"1e",x"00"),
   805 => (x"0f",x"00",x"00",x"03"),
   806 => (x"dc",x"27",x"86",x"c4"),
   807 => (x"1e",x"00",x"00",x"16"),
   808 => (x"00",x"03",x"03",x"27"),
   809 => (x"86",x"c4",x"0f",x"00"),
   810 => (x"00",x"3e",x"fc",x"27"),
   811 => (x"27",x"49",x"bf",x"00"),
   812 => (x"00",x"00",x"3e",x"f8"),
   813 => (x"04",x"27",x"89",x"bf"),
   814 => (x"59",x"00",x"00",x"3f"),
   815 => (x"de",x"27",x"1e",x"71"),
   816 => (x"1e",x"00",x"00",x"16"),
   817 => (x"00",x"03",x"03",x"27"),
   818 => (x"86",x"c8",x"0f",x"00"),
   819 => (x"00",x"3f",x"00",x"27"),
   820 => (x"c1",x"48",x"bf",x"00"),
   821 => (x"03",x"a8",x"b7",x"f8"),
   822 => (x"27",x"87",x"ea",x"c0"),
   823 => (x"00",x"00",x"0f",x"ee"),
   824 => (x"03",x"03",x"27",x"1e"),
   825 => (x"c4",x"0f",x"00",x"00"),
   826 => (x"10",x"24",x"27",x"86"),
   827 => (x"27",x"1e",x"00",x"00"),
   828 => (x"00",x"00",x"03",x"03"),
   829 => (x"27",x"86",x"c4",x"0f"),
   830 => (x"00",x"00",x"10",x"44"),
   831 => (x"03",x"03",x"27",x"1e"),
   832 => (x"c4",x"0f",x"00",x"00"),
   833 => (x"3f",x"00",x"27",x"86"),
   834 => (x"49",x"bf",x"00",x"00"),
   835 => (x"e8",x"cf",x"4a",x"71"),
   836 => (x"72",x"1e",x"71",x"92"),
   837 => (x"27",x"49",x"72",x"1e"),
   838 => (x"00",x"00",x"16",x"f4"),
   839 => (x"f8",x"27",x"4a",x"bf"),
   840 => (x"0f",x"00",x"00",x"05"),
   841 => (x"49",x"26",x"4a",x"26"),
   842 => (x"00",x"3f",x"08",x"27"),
   843 => (x"f4",x"27",x"58",x"00"),
   844 => (x"bf",x"00",x"00",x"16"),
   845 => (x"cf",x"4b",x"72",x"4a"),
   846 => (x"1e",x"71",x"93",x"e8"),
   847 => (x"09",x"73",x"1e",x"72"),
   848 => (x"05",x"f8",x"27",x"4a"),
   849 => (x"26",x"0f",x"00",x"00"),
   850 => (x"27",x"49",x"26",x"4a"),
   851 => (x"00",x"00",x"3f",x"0c"),
   852 => (x"92",x"f9",x"c8",x"58"),
   853 => (x"1e",x"72",x"1e",x"71"),
   854 => (x"27",x"4a",x"09",x"72"),
   855 => (x"00",x"00",x"05",x"f8"),
   856 => (x"26",x"4a",x"26",x"0f"),
   857 => (x"3f",x"10",x"27",x"49"),
   858 => (x"27",x"58",x"00",x"00"),
   859 => (x"00",x"00",x"10",x"46"),
   860 => (x"03",x"03",x"27",x"1e"),
   861 => (x"c4",x"0f",x"00",x"00"),
   862 => (x"3f",x"04",x"27",x"86"),
   863 => (x"1e",x"bf",x"00",x"00"),
   864 => (x"00",x"10",x"73",x"27"),
   865 => (x"03",x"27",x"1e",x"00"),
   866 => (x"0f",x"00",x"00",x"03"),
   867 => (x"78",x"27",x"86",x"c8"),
   868 => (x"1e",x"00",x"00",x"10"),
   869 => (x"00",x"03",x"03",x"27"),
   870 => (x"86",x"c4",x"0f",x"00"),
   871 => (x"00",x"3f",x"08",x"27"),
   872 => (x"27",x"1e",x"bf",x"00"),
   873 => (x"00",x"00",x"10",x"a5"),
   874 => (x"03",x"03",x"27",x"1e"),
   875 => (x"c8",x"0f",x"00",x"00"),
   876 => (x"3f",x"0c",x"27",x"86"),
   877 => (x"1e",x"bf",x"00",x"00"),
   878 => (x"00",x"10",x"aa",x"27"),
   879 => (x"03",x"27",x"1e",x"00"),
   880 => (x"0f",x"00",x"00",x"03"),
   881 => (x"c8",x"27",x"86",x"c8"),
   882 => (x"1e",x"00",x"00",x"10"),
   883 => (x"00",x"03",x"03",x"27"),
   884 => (x"86",x"c4",x"0f",x"00"),
   885 => (x"8e",x"f0",x"48",x"c0"),
   886 => (x"4c",x"26",x"4d",x"26"),
   887 => (x"4f",x"26",x"4b",x"26"),
   888 => (x"5c",x"5b",x"5e",x"0e"),
   889 => (x"66",x"d0",x"0e",x"5d"),
   890 => (x"73",x"4b",x"6d",x"4d"),
   891 => (x"27",x"1e",x"73",x"4c"),
   892 => (x"00",x"00",x"17",x"08"),
   893 => (x"f0",x"c0",x"48",x"bf"),
   894 => (x"43",x"20",x"4a",x"a3"),
   895 => (x"f9",x"05",x"aa",x"73"),
   896 => (x"75",x"4a",x"26",x"87"),
   897 => (x"c5",x"82",x"cc",x"4a"),
   898 => (x"cc",x"49",x"73",x"7a"),
   899 => (x"6d",x"79",x"6a",x"81"),
   900 => (x"27",x"1e",x"73",x"7b"),
   901 => (x"00",x"00",x"0e",x"bf"),
   902 => (x"73",x"86",x"c4",x"0f"),
   903 => (x"69",x"81",x"c4",x"49"),
   904 => (x"87",x"f3",x"c0",x"05"),
   905 => (x"81",x"c8",x"49",x"74"),
   906 => (x"83",x"cc",x"4b",x"74"),
   907 => (x"1e",x"71",x"7b",x"c6"),
   908 => (x"81",x"c8",x"49",x"75"),
   909 => (x"be",x"27",x"1e",x"69"),
   910 => (x"0f",x"00",x"00",x"03"),
   911 => (x"08",x"27",x"86",x"c8"),
   912 => (x"bf",x"00",x"00",x"17"),
   913 => (x"1e",x"73",x"7c",x"bf"),
   914 => (x"1e",x"6b",x"1e",x"ca"),
   915 => (x"00",x"04",x"26",x"27"),
   916 => (x"86",x"cc",x"0f",x"00"),
   917 => (x"6d",x"87",x"d0",x"c0"),
   918 => (x"48",x"4a",x"75",x"49"),
   919 => (x"4b",x"a2",x"f0",x"c0"),
   920 => (x"ab",x"72",x"42",x"20"),
   921 => (x"26",x"87",x"f9",x"05"),
   922 => (x"26",x"4c",x"26",x"4d"),
   923 => (x"0e",x"4f",x"26",x"4b"),
   924 => (x"5d",x"5c",x"5b",x"5e"),
   925 => (x"27",x"86",x"fc",x"0e"),
   926 => (x"00",x"00",x"17",x"18"),
   927 => (x"6e",x"4d",x"bf",x"97"),
   928 => (x"4b",x"66",x"d4",x"4c"),
   929 => (x"82",x"ca",x"4a",x"6b"),
   930 => (x"c0",x"fe",x"49",x"75"),
   931 => (x"04",x"b1",x"03",x"81"),
   932 => (x"c1",x"c1",x"07",x"b9"),
   933 => (x"cf",x"c0",x"05",x"a9"),
   934 => (x"72",x"8a",x"c1",x"87"),
   935 => (x"17",x"10",x"27",x"48"),
   936 => (x"88",x"bf",x"00",x"00"),
   937 => (x"4c",x"c0",x"7b",x"70"),
   938 => (x"ff",x"05",x"9c",x"74"),
   939 => (x"1c",x"27",x"87",x"da"),
   940 => (x"97",x"00",x"00",x"17"),
   941 => (x"26",x"8e",x"fc",x"5d"),
   942 => (x"26",x"4c",x"26",x"4d"),
   943 => (x"1e",x"4f",x"26",x"4b"),
   944 => (x"00",x"17",x"08",x"27"),
   945 => (x"c0",x"02",x"bf",x"00"),
   946 => (x"66",x"c4",x"87",x"cb"),
   947 => (x"17",x"08",x"27",x"48"),
   948 => (x"bf",x"bf",x"00",x"00"),
   949 => (x"17",x"08",x"27",x"78"),
   950 => (x"49",x"bf",x"00",x"00"),
   951 => (x"1e",x"71",x"81",x"cc"),
   952 => (x"00",x"17",x"10",x"27"),
   953 => (x"ca",x"1e",x"bf",x"00"),
   954 => (x"04",x"26",x"27",x"1e"),
   955 => (x"cc",x"0f",x"00",x"00"),
   956 => (x"1e",x"4f",x"26",x"86"),
   957 => (x"00",x"17",x"18",x"27"),
   958 => (x"49",x"bf",x"97",x"00"),
   959 => (x"03",x"81",x"c0",x"fe"),
   960 => (x"07",x"b9",x"04",x"b1"),
   961 => (x"02",x"a9",x"c1",x"c1"),
   962 => (x"c0",x"87",x"c5",x"c0"),
   963 => (x"87",x"c2",x"c0",x"49"),
   964 => (x"14",x"27",x"49",x"c1"),
   965 => (x"bf",x"00",x"00",x"17"),
   966 => (x"27",x"b0",x"71",x"48"),
   967 => (x"00",x"00",x"17",x"18"),
   968 => (x"17",x"19",x"27",x"58"),
   969 => (x"c1",x"48",x"00",x"00"),
   970 => (x"4f",x"26",x"50",x"c2"),
   971 => (x"17",x"18",x"27",x"1e"),
   972 => (x"c1",x"48",x"00",x"00"),
   973 => (x"14",x"27",x"50",x"c1"),
   974 => (x"48",x"00",x"00",x"17"),
   975 => (x"4f",x"26",x"78",x"c0"),
   976 => (x"33",x"32",x"31",x"30"),
   977 => (x"37",x"36",x"35",x"34"),
   978 => (x"42",x"41",x"39",x"38"),
   979 => (x"46",x"45",x"44",x"43"),
   980 => (x"6f",x"72",x"50",x"00"),
   981 => (x"6d",x"61",x"72",x"67"),
   982 => (x"6d",x"6f",x"63",x"20"),
   983 => (x"65",x"6c",x"69",x"70"),
   984 => (x"69",x"77",x"20",x"64"),
   985 => (x"27",x"20",x"68",x"74"),
   986 => (x"69",x"67",x"65",x"72"),
   987 => (x"72",x"65",x"74",x"73"),
   988 => (x"74",x"61",x"20",x"27"),
   989 => (x"62",x"69",x"72",x"74"),
   990 => (x"0a",x"65",x"74",x"75"),
   991 => (x"50",x"00",x"0a",x"00"),
   992 => (x"72",x"67",x"6f",x"72"),
   993 => (x"63",x"20",x"6d",x"61"),
   994 => (x"69",x"70",x"6d",x"6f"),
   995 => (x"20",x"64",x"65",x"6c"),
   996 => (x"68",x"74",x"69",x"77"),
   997 => (x"20",x"74",x"75",x"6f"),
   998 => (x"67",x"65",x"72",x"27"),
   999 => (x"65",x"74",x"73",x"69"),
  1000 => (x"61",x"20",x"27",x"72"),
  1001 => (x"69",x"72",x"74",x"74"),
  1002 => (x"65",x"74",x"75",x"62"),
  1003 => (x"00",x"0a",x"00",x"0a"),
  1004 => (x"59",x"52",x"48",x"44"),
  1005 => (x"4e",x"4f",x"54",x"53"),
  1006 => (x"52",x"50",x"20",x"45"),
  1007 => (x"41",x"52",x"47",x"4f"),
  1008 => (x"33",x"20",x"2c",x"4d"),
  1009 => (x"20",x"44",x"52",x"27"),
  1010 => (x"49",x"52",x"54",x"53"),
  1011 => (x"44",x"00",x"47",x"4e"),
  1012 => (x"53",x"59",x"52",x"48"),
  1013 => (x"45",x"4e",x"4f",x"54"),
  1014 => (x"4f",x"52",x"50",x"20"),
  1015 => (x"4d",x"41",x"52",x"47"),
  1016 => (x"27",x"32",x"20",x"2c"),
  1017 => (x"53",x"20",x"44",x"4e"),
  1018 => (x"4e",x"49",x"52",x"54"),
  1019 => (x"65",x"4d",x"00",x"47"),
  1020 => (x"72",x"75",x"73",x"61"),
  1021 => (x"74",x"20",x"64",x"65"),
  1022 => (x"20",x"65",x"6d",x"69"),
  1023 => (x"20",x"6f",x"6f",x"74"),
  1024 => (x"6c",x"61",x"6d",x"73"),
  1025 => (x"6f",x"74",x"20",x"6c"),
  1026 => (x"74",x"62",x"6f",x"20"),
  1027 => (x"20",x"6e",x"69",x"61"),
  1028 => (x"6e",x"61",x"65",x"6d"),
  1029 => (x"66",x"67",x"6e",x"69"),
  1030 => (x"72",x"20",x"6c",x"75"),
  1031 => (x"6c",x"75",x"73",x"65"),
  1032 => (x"00",x"0a",x"73",x"74"),
  1033 => (x"61",x"65",x"6c",x"50"),
  1034 => (x"69",x"20",x"65",x"73"),
  1035 => (x"65",x"72",x"63",x"6e"),
  1036 => (x"20",x"65",x"73",x"61"),
  1037 => (x"62",x"6d",x"75",x"6e"),
  1038 => (x"6f",x"20",x"72",x"65"),
  1039 => (x"75",x"72",x"20",x"66"),
  1040 => (x"00",x"0a",x"73",x"6e"),
  1041 => (x"69",x"4d",x"00",x"0a"),
  1042 => (x"73",x"6f",x"72",x"63"),
  1043 => (x"6e",x"6f",x"63",x"65"),
  1044 => (x"66",x"20",x"73",x"64"),
  1045 => (x"6f",x"20",x"72",x"6f"),
  1046 => (x"72",x"20",x"65",x"6e"),
  1047 => (x"74",x"20",x"6e",x"75"),
  1048 => (x"75",x"6f",x"72",x"68"),
  1049 => (x"44",x"20",x"68",x"67"),
  1050 => (x"73",x"79",x"72",x"68"),
  1051 => (x"65",x"6e",x"6f",x"74"),
  1052 => (x"25",x"00",x"20",x"3a"),
  1053 => (x"00",x"0a",x"20",x"64"),
  1054 => (x"79",x"72",x"68",x"44"),
  1055 => (x"6e",x"6f",x"74",x"73"),
  1056 => (x"70",x"20",x"73",x"65"),
  1057 => (x"53",x"20",x"72",x"65"),
  1058 => (x"6e",x"6f",x"63",x"65"),
  1059 => (x"20",x"20",x"3a",x"64"),
  1060 => (x"20",x"20",x"20",x"20"),
  1061 => (x"20",x"20",x"20",x"20"),
  1062 => (x"20",x"20",x"20",x"20"),
  1063 => (x"20",x"20",x"20",x"20"),
  1064 => (x"20",x"20",x"20",x"20"),
  1065 => (x"20",x"64",x"25",x"00"),
  1066 => (x"41",x"56",x"00",x"0a"),
  1067 => (x"49",x"4d",x"20",x"58"),
  1068 => (x"72",x"20",x"53",x"50"),
  1069 => (x"6e",x"69",x"74",x"61"),
  1070 => (x"20",x"2a",x"20",x"67"),
  1071 => (x"30",x"30",x"30",x"31"),
  1072 => (x"25",x"20",x"3d",x"20"),
  1073 => (x"00",x"0a",x"20",x"64"),
  1074 => (x"48",x"44",x"00",x"0a"),
  1075 => (x"54",x"53",x"59",x"52"),
  1076 => (x"20",x"45",x"4e",x"4f"),
  1077 => (x"47",x"4f",x"52",x"50"),
  1078 => (x"2c",x"4d",x"41",x"52"),
  1079 => (x"4d",x"4f",x"53",x"20"),
  1080 => (x"54",x"53",x"20",x"45"),
  1081 => (x"47",x"4e",x"49",x"52"),
  1082 => (x"52",x"48",x"44",x"00"),
  1083 => (x"4f",x"54",x"53",x"59"),
  1084 => (x"50",x"20",x"45",x"4e"),
  1085 => (x"52",x"47",x"4f",x"52"),
  1086 => (x"20",x"2c",x"4d",x"41"),
  1087 => (x"54",x"53",x"27",x"31"),
  1088 => (x"52",x"54",x"53",x"20"),
  1089 => (x"00",x"47",x"4e",x"49"),
  1090 => (x"68",x"44",x"00",x"0a"),
  1091 => (x"74",x"73",x"79",x"72"),
  1092 => (x"20",x"65",x"6e",x"6f"),
  1093 => (x"63",x"6e",x"65",x"42"),
  1094 => (x"72",x"61",x"6d",x"68"),
  1095 => (x"56",x"20",x"2c",x"6b"),
  1096 => (x"69",x"73",x"72",x"65"),
  1097 => (x"32",x"20",x"6e",x"6f"),
  1098 => (x"28",x"20",x"31",x"2e"),
  1099 => (x"67",x"6e",x"61",x"4c"),
  1100 => (x"65",x"67",x"61",x"75"),
  1101 => (x"29",x"43",x"20",x"3a"),
  1102 => (x"00",x"0a",x"00",x"0a"),
  1103 => (x"63",x"65",x"78",x"45"),
  1104 => (x"6f",x"69",x"74",x"75"),
  1105 => (x"74",x"73",x"20",x"6e"),
  1106 => (x"73",x"74",x"72",x"61"),
  1107 => (x"64",x"25",x"20",x"2c"),
  1108 => (x"6e",x"75",x"72",x"20"),
  1109 => (x"68",x"74",x"20",x"73"),
  1110 => (x"67",x"75",x"6f",x"72"),
  1111 => (x"68",x"44",x"20",x"68"),
  1112 => (x"74",x"73",x"79",x"72"),
  1113 => (x"0a",x"65",x"6e",x"6f"),
  1114 => (x"65",x"78",x"45",x"00"),
  1115 => (x"69",x"74",x"75",x"63"),
  1116 => (x"65",x"20",x"6e",x"6f"),
  1117 => (x"0a",x"73",x"64",x"6e"),
  1118 => (x"46",x"00",x"0a",x"00"),
  1119 => (x"6c",x"61",x"6e",x"69"),
  1120 => (x"6c",x"61",x"76",x"20"),
  1121 => (x"20",x"73",x"65",x"75"),
  1122 => (x"74",x"20",x"66",x"6f"),
  1123 => (x"76",x"20",x"65",x"68"),
  1124 => (x"61",x"69",x"72",x"61"),
  1125 => (x"73",x"65",x"6c",x"62"),
  1126 => (x"65",x"73",x"75",x"20"),
  1127 => (x"6e",x"69",x"20",x"64"),
  1128 => (x"65",x"68",x"74",x"20"),
  1129 => (x"6e",x"65",x"62",x"20"),
  1130 => (x"61",x"6d",x"68",x"63"),
  1131 => (x"0a",x"3a",x"6b",x"72"),
  1132 => (x"49",x"00",x"0a",x"00"),
  1133 => (x"47",x"5f",x"74",x"6e"),
  1134 => (x"3a",x"62",x"6f",x"6c"),
  1135 => (x"20",x"20",x"20",x"20"),
  1136 => (x"20",x"20",x"20",x"20"),
  1137 => (x"20",x"20",x"20",x"20"),
  1138 => (x"00",x"0a",x"64",x"25"),
  1139 => (x"20",x"20",x"20",x"20"),
  1140 => (x"20",x"20",x"20",x"20"),
  1141 => (x"75",x"6f",x"68",x"73"),
  1142 => (x"62",x"20",x"64",x"6c"),
  1143 => (x"20",x"20",x"3a",x"65"),
  1144 => (x"0a",x"64",x"25",x"20"),
  1145 => (x"6f",x"6f",x"42",x"00"),
  1146 => (x"6c",x"47",x"5f",x"6c"),
  1147 => (x"20",x"3a",x"62",x"6f"),
  1148 => (x"20",x"20",x"20",x"20"),
  1149 => (x"20",x"20",x"20",x"20"),
  1150 => (x"64",x"25",x"20",x"20"),
  1151 => (x"20",x"20",x"00",x"0a"),
  1152 => (x"20",x"20",x"20",x"20"),
  1153 => (x"68",x"73",x"20",x"20"),
  1154 => (x"64",x"6c",x"75",x"6f"),
  1155 => (x"3a",x"65",x"62",x"20"),
  1156 => (x"25",x"20",x"20",x"20"),
  1157 => (x"43",x"00",x"0a",x"64"),
  1158 => (x"5f",x"31",x"5f",x"68"),
  1159 => (x"62",x"6f",x"6c",x"47"),
  1160 => (x"20",x"20",x"20",x"3a"),
  1161 => (x"20",x"20",x"20",x"20"),
  1162 => (x"20",x"20",x"20",x"20"),
  1163 => (x"00",x"0a",x"63",x"25"),
  1164 => (x"20",x"20",x"20",x"20"),
  1165 => (x"20",x"20",x"20",x"20"),
  1166 => (x"75",x"6f",x"68",x"73"),
  1167 => (x"62",x"20",x"64",x"6c"),
  1168 => (x"20",x"20",x"3a",x"65"),
  1169 => (x"0a",x"63",x"25",x"20"),
  1170 => (x"5f",x"68",x"43",x"00"),
  1171 => (x"6c",x"47",x"5f",x"32"),
  1172 => (x"20",x"3a",x"62",x"6f"),
  1173 => (x"20",x"20",x"20",x"20"),
  1174 => (x"20",x"20",x"20",x"20"),
  1175 => (x"63",x"25",x"20",x"20"),
  1176 => (x"20",x"20",x"00",x"0a"),
  1177 => (x"20",x"20",x"20",x"20"),
  1178 => (x"68",x"73",x"20",x"20"),
  1179 => (x"64",x"6c",x"75",x"6f"),
  1180 => (x"3a",x"65",x"62",x"20"),
  1181 => (x"25",x"20",x"20",x"20"),
  1182 => (x"41",x"00",x"0a",x"63"),
  1183 => (x"31",x"5f",x"72",x"72"),
  1184 => (x"6f",x"6c",x"47",x"5f"),
  1185 => (x"5d",x"38",x"5b",x"62"),
  1186 => (x"20",x"20",x"20",x"3a"),
  1187 => (x"20",x"20",x"20",x"20"),
  1188 => (x"00",x"0a",x"64",x"25"),
  1189 => (x"20",x"20",x"20",x"20"),
  1190 => (x"20",x"20",x"20",x"20"),
  1191 => (x"75",x"6f",x"68",x"73"),
  1192 => (x"62",x"20",x"64",x"6c"),
  1193 => (x"20",x"20",x"3a",x"65"),
  1194 => (x"0a",x"64",x"25",x"20"),
  1195 => (x"72",x"72",x"41",x"00"),
  1196 => (x"47",x"5f",x"32",x"5f"),
  1197 => (x"5b",x"62",x"6f",x"6c"),
  1198 => (x"37",x"5b",x"5d",x"38"),
  1199 => (x"20",x"20",x"3a",x"5d"),
  1200 => (x"64",x"25",x"20",x"20"),
  1201 => (x"20",x"20",x"00",x"0a"),
  1202 => (x"20",x"20",x"20",x"20"),
  1203 => (x"68",x"73",x"20",x"20"),
  1204 => (x"64",x"6c",x"75",x"6f"),
  1205 => (x"3a",x"65",x"62",x"20"),
  1206 => (x"4e",x"20",x"20",x"20"),
  1207 => (x"65",x"62",x"6d",x"75"),
  1208 => (x"66",x"4f",x"5f",x"72"),
  1209 => (x"6e",x"75",x"52",x"5f"),
  1210 => (x"20",x"2b",x"20",x"73"),
  1211 => (x"00",x"0a",x"30",x"31"),
  1212 => (x"5f",x"72",x"74",x"50"),
  1213 => (x"62",x"6f",x"6c",x"47"),
  1214 => (x"00",x"0a",x"3e",x"2d"),
  1215 => (x"74",x"50",x"20",x"20"),
  1216 => (x"6f",x"43",x"5f",x"72"),
  1217 => (x"20",x"3a",x"70",x"6d"),
  1218 => (x"20",x"20",x"20",x"20"),
  1219 => (x"20",x"20",x"20",x"20"),
  1220 => (x"0a",x"64",x"25",x"20"),
  1221 => (x"20",x"20",x"20",x"00"),
  1222 => (x"20",x"20",x"20",x"20"),
  1223 => (x"6f",x"68",x"73",x"20"),
  1224 => (x"20",x"64",x"6c",x"75"),
  1225 => (x"20",x"3a",x"65",x"62"),
  1226 => (x"69",x"28",x"20",x"20"),
  1227 => (x"65",x"6c",x"70",x"6d"),
  1228 => (x"74",x"6e",x"65",x"6d"),
  1229 => (x"6f",x"69",x"74",x"61"),
  1230 => (x"65",x"64",x"2d",x"6e"),
  1231 => (x"64",x"6e",x"65",x"70"),
  1232 => (x"29",x"74",x"6e",x"65"),
  1233 => (x"20",x"20",x"00",x"0a"),
  1234 => (x"63",x"73",x"69",x"44"),
  1235 => (x"20",x"20",x"3a",x"72"),
  1236 => (x"20",x"20",x"20",x"20"),
  1237 => (x"20",x"20",x"20",x"20"),
  1238 => (x"25",x"20",x"20",x"20"),
  1239 => (x"20",x"00",x"0a",x"64"),
  1240 => (x"20",x"20",x"20",x"20"),
  1241 => (x"73",x"20",x"20",x"20"),
  1242 => (x"6c",x"75",x"6f",x"68"),
  1243 => (x"65",x"62",x"20",x"64"),
  1244 => (x"20",x"20",x"20",x"3a"),
  1245 => (x"00",x"0a",x"64",x"25"),
  1246 => (x"6e",x"45",x"20",x"20"),
  1247 => (x"43",x"5f",x"6d",x"75"),
  1248 => (x"3a",x"70",x"6d",x"6f"),
  1249 => (x"20",x"20",x"20",x"20"),
  1250 => (x"20",x"20",x"20",x"20"),
  1251 => (x"0a",x"64",x"25",x"20"),
  1252 => (x"20",x"20",x"20",x"00"),
  1253 => (x"20",x"20",x"20",x"20"),
  1254 => (x"6f",x"68",x"73",x"20"),
  1255 => (x"20",x"64",x"6c",x"75"),
  1256 => (x"20",x"3a",x"65",x"62"),
  1257 => (x"64",x"25",x"20",x"20"),
  1258 => (x"20",x"20",x"00",x"0a"),
  1259 => (x"5f",x"74",x"6e",x"49"),
  1260 => (x"70",x"6d",x"6f",x"43"),
  1261 => (x"20",x"20",x"20",x"3a"),
  1262 => (x"20",x"20",x"20",x"20"),
  1263 => (x"25",x"20",x"20",x"20"),
  1264 => (x"20",x"00",x"0a",x"64"),
  1265 => (x"20",x"20",x"20",x"20"),
  1266 => (x"73",x"20",x"20",x"20"),
  1267 => (x"6c",x"75",x"6f",x"68"),
  1268 => (x"65",x"62",x"20",x"64"),
  1269 => (x"20",x"20",x"20",x"3a"),
  1270 => (x"00",x"0a",x"64",x"25"),
  1271 => (x"74",x"53",x"20",x"20"),
  1272 => (x"6f",x"43",x"5f",x"72"),
  1273 => (x"20",x"3a",x"70",x"6d"),
  1274 => (x"20",x"20",x"20",x"20"),
  1275 => (x"20",x"20",x"20",x"20"),
  1276 => (x"0a",x"73",x"25",x"20"),
  1277 => (x"20",x"20",x"20",x"00"),
  1278 => (x"20",x"20",x"20",x"20"),
  1279 => (x"6f",x"68",x"73",x"20"),
  1280 => (x"20",x"64",x"6c",x"75"),
  1281 => (x"20",x"3a",x"65",x"62"),
  1282 => (x"48",x"44",x"20",x"20"),
  1283 => (x"54",x"53",x"59",x"52"),
  1284 => (x"20",x"45",x"4e",x"4f"),
  1285 => (x"47",x"4f",x"52",x"50"),
  1286 => (x"2c",x"4d",x"41",x"52"),
  1287 => (x"4d",x"4f",x"53",x"20"),
  1288 => (x"54",x"53",x"20",x"45"),
  1289 => (x"47",x"4e",x"49",x"52"),
  1290 => (x"65",x"4e",x"00",x"0a"),
  1291 => (x"50",x"5f",x"74",x"78"),
  1292 => (x"47",x"5f",x"72",x"74"),
  1293 => (x"2d",x"62",x"6f",x"6c"),
  1294 => (x"20",x"00",x"0a",x"3e"),
  1295 => (x"72",x"74",x"50",x"20"),
  1296 => (x"6d",x"6f",x"43",x"5f"),
  1297 => (x"20",x"20",x"3a",x"70"),
  1298 => (x"20",x"20",x"20",x"20"),
  1299 => (x"20",x"20",x"20",x"20"),
  1300 => (x"00",x"0a",x"64",x"25"),
  1301 => (x"20",x"20",x"20",x"20"),
  1302 => (x"20",x"20",x"20",x"20"),
  1303 => (x"75",x"6f",x"68",x"73"),
  1304 => (x"62",x"20",x"64",x"6c"),
  1305 => (x"20",x"20",x"3a",x"65"),
  1306 => (x"6d",x"69",x"28",x"20"),
  1307 => (x"6d",x"65",x"6c",x"70"),
  1308 => (x"61",x"74",x"6e",x"65"),
  1309 => (x"6e",x"6f",x"69",x"74"),
  1310 => (x"70",x"65",x"64",x"2d"),
  1311 => (x"65",x"64",x"6e",x"65"),
  1312 => (x"2c",x"29",x"74",x"6e"),
  1313 => (x"6d",x"61",x"73",x"20"),
  1314 => (x"73",x"61",x"20",x"65"),
  1315 => (x"6f",x"62",x"61",x"20"),
  1316 => (x"00",x"0a",x"65",x"76"),
  1317 => (x"69",x"44",x"20",x"20"),
  1318 => (x"3a",x"72",x"63",x"73"),
  1319 => (x"20",x"20",x"20",x"20"),
  1320 => (x"20",x"20",x"20",x"20"),
  1321 => (x"20",x"20",x"20",x"20"),
  1322 => (x"0a",x"64",x"25",x"20"),
  1323 => (x"20",x"20",x"20",x"00"),
  1324 => (x"20",x"20",x"20",x"20"),
  1325 => (x"6f",x"68",x"73",x"20"),
  1326 => (x"20",x"64",x"6c",x"75"),
  1327 => (x"20",x"3a",x"65",x"62"),
  1328 => (x"64",x"25",x"20",x"20"),
  1329 => (x"20",x"20",x"00",x"0a"),
  1330 => (x"6d",x"75",x"6e",x"45"),
  1331 => (x"6d",x"6f",x"43",x"5f"),
  1332 => (x"20",x"20",x"3a",x"70"),
  1333 => (x"20",x"20",x"20",x"20"),
  1334 => (x"25",x"20",x"20",x"20"),
  1335 => (x"20",x"00",x"0a",x"64"),
  1336 => (x"20",x"20",x"20",x"20"),
  1337 => (x"73",x"20",x"20",x"20"),
  1338 => (x"6c",x"75",x"6f",x"68"),
  1339 => (x"65",x"62",x"20",x"64"),
  1340 => (x"20",x"20",x"20",x"3a"),
  1341 => (x"00",x"0a",x"64",x"25"),
  1342 => (x"6e",x"49",x"20",x"20"),
  1343 => (x"6f",x"43",x"5f",x"74"),
  1344 => (x"20",x"3a",x"70",x"6d"),
  1345 => (x"20",x"20",x"20",x"20"),
  1346 => (x"20",x"20",x"20",x"20"),
  1347 => (x"0a",x"64",x"25",x"20"),
  1348 => (x"20",x"20",x"20",x"00"),
  1349 => (x"20",x"20",x"20",x"20"),
  1350 => (x"6f",x"68",x"73",x"20"),
  1351 => (x"20",x"64",x"6c",x"75"),
  1352 => (x"20",x"3a",x"65",x"62"),
  1353 => (x"64",x"25",x"20",x"20"),
  1354 => (x"20",x"20",x"00",x"0a"),
  1355 => (x"5f",x"72",x"74",x"53"),
  1356 => (x"70",x"6d",x"6f",x"43"),
  1357 => (x"20",x"20",x"20",x"3a"),
  1358 => (x"20",x"20",x"20",x"20"),
  1359 => (x"25",x"20",x"20",x"20"),
  1360 => (x"20",x"00",x"0a",x"73"),
  1361 => (x"20",x"20",x"20",x"20"),
  1362 => (x"73",x"20",x"20",x"20"),
  1363 => (x"6c",x"75",x"6f",x"68"),
  1364 => (x"65",x"62",x"20",x"64"),
  1365 => (x"20",x"20",x"20",x"3a"),
  1366 => (x"59",x"52",x"48",x"44"),
  1367 => (x"4e",x"4f",x"54",x"53"),
  1368 => (x"52",x"50",x"20",x"45"),
  1369 => (x"41",x"52",x"47",x"4f"),
  1370 => (x"53",x"20",x"2c",x"4d"),
  1371 => (x"20",x"45",x"4d",x"4f"),
  1372 => (x"49",x"52",x"54",x"53"),
  1373 => (x"00",x"0a",x"47",x"4e"),
  1374 => (x"5f",x"74",x"6e",x"49"),
  1375 => (x"6f",x"4c",x"5f",x"31"),
  1376 => (x"20",x"20",x"3a",x"63"),
  1377 => (x"20",x"20",x"20",x"20"),
  1378 => (x"20",x"20",x"20",x"20"),
  1379 => (x"0a",x"64",x"25",x"20"),
  1380 => (x"20",x"20",x"20",x"00"),
  1381 => (x"20",x"20",x"20",x"20"),
  1382 => (x"6f",x"68",x"73",x"20"),
  1383 => (x"20",x"64",x"6c",x"75"),
  1384 => (x"20",x"3a",x"65",x"62"),
  1385 => (x"64",x"25",x"20",x"20"),
  1386 => (x"6e",x"49",x"00",x"0a"),
  1387 => (x"5f",x"32",x"5f",x"74"),
  1388 => (x"3a",x"63",x"6f",x"4c"),
  1389 => (x"20",x"20",x"20",x"20"),
  1390 => (x"20",x"20",x"20",x"20"),
  1391 => (x"25",x"20",x"20",x"20"),
  1392 => (x"20",x"00",x"0a",x"64"),
  1393 => (x"20",x"20",x"20",x"20"),
  1394 => (x"73",x"20",x"20",x"20"),
  1395 => (x"6c",x"75",x"6f",x"68"),
  1396 => (x"65",x"62",x"20",x"64"),
  1397 => (x"20",x"20",x"20",x"3a"),
  1398 => (x"00",x"0a",x"64",x"25"),
  1399 => (x"5f",x"74",x"6e",x"49"),
  1400 => (x"6f",x"4c",x"5f",x"33"),
  1401 => (x"20",x"20",x"3a",x"63"),
  1402 => (x"20",x"20",x"20",x"20"),
  1403 => (x"20",x"20",x"20",x"20"),
  1404 => (x"0a",x"64",x"25",x"20"),
  1405 => (x"20",x"20",x"20",x"00"),
  1406 => (x"20",x"20",x"20",x"20"),
  1407 => (x"6f",x"68",x"73",x"20"),
  1408 => (x"20",x"64",x"6c",x"75"),
  1409 => (x"20",x"3a",x"65",x"62"),
  1410 => (x"64",x"25",x"20",x"20"),
  1411 => (x"6e",x"45",x"00",x"0a"),
  1412 => (x"4c",x"5f",x"6d",x"75"),
  1413 => (x"20",x"3a",x"63",x"6f"),
  1414 => (x"20",x"20",x"20",x"20"),
  1415 => (x"20",x"20",x"20",x"20"),
  1416 => (x"25",x"20",x"20",x"20"),
  1417 => (x"20",x"00",x"0a",x"64"),
  1418 => (x"20",x"20",x"20",x"20"),
  1419 => (x"73",x"20",x"20",x"20"),
  1420 => (x"6c",x"75",x"6f",x"68"),
  1421 => (x"65",x"62",x"20",x"64"),
  1422 => (x"20",x"20",x"20",x"3a"),
  1423 => (x"00",x"0a",x"64",x"25"),
  1424 => (x"5f",x"72",x"74",x"53"),
  1425 => (x"6f",x"4c",x"5f",x"31"),
  1426 => (x"20",x"20",x"3a",x"63"),
  1427 => (x"20",x"20",x"20",x"20"),
  1428 => (x"20",x"20",x"20",x"20"),
  1429 => (x"0a",x"73",x"25",x"20"),
  1430 => (x"20",x"20",x"20",x"00"),
  1431 => (x"20",x"20",x"20",x"20"),
  1432 => (x"6f",x"68",x"73",x"20"),
  1433 => (x"20",x"64",x"6c",x"75"),
  1434 => (x"20",x"3a",x"65",x"62"),
  1435 => (x"48",x"44",x"20",x"20"),
  1436 => (x"54",x"53",x"59",x"52"),
  1437 => (x"20",x"45",x"4e",x"4f"),
  1438 => (x"47",x"4f",x"52",x"50"),
  1439 => (x"2c",x"4d",x"41",x"52"),
  1440 => (x"53",x"27",x"31",x"20"),
  1441 => (x"54",x"53",x"20",x"54"),
  1442 => (x"47",x"4e",x"49",x"52"),
  1443 => (x"74",x"53",x"00",x"0a"),
  1444 => (x"5f",x"32",x"5f",x"72"),
  1445 => (x"3a",x"63",x"6f",x"4c"),
  1446 => (x"20",x"20",x"20",x"20"),
  1447 => (x"20",x"20",x"20",x"20"),
  1448 => (x"25",x"20",x"20",x"20"),
  1449 => (x"20",x"00",x"0a",x"73"),
  1450 => (x"20",x"20",x"20",x"20"),
  1451 => (x"73",x"20",x"20",x"20"),
  1452 => (x"6c",x"75",x"6f",x"68"),
  1453 => (x"65",x"62",x"20",x"64"),
  1454 => (x"20",x"20",x"20",x"3a"),
  1455 => (x"59",x"52",x"48",x"44"),
  1456 => (x"4e",x"4f",x"54",x"53"),
  1457 => (x"52",x"50",x"20",x"45"),
  1458 => (x"41",x"52",x"47",x"4f"),
  1459 => (x"32",x"20",x"2c",x"4d"),
  1460 => (x"20",x"44",x"4e",x"27"),
  1461 => (x"49",x"52",x"54",x"53"),
  1462 => (x"00",x"0a",x"47",x"4e"),
  1463 => (x"73",x"55",x"00",x"0a"),
  1464 => (x"74",x"20",x"72",x"65"),
  1465 => (x"3a",x"65",x"6d",x"69"),
  1466 => (x"0a",x"64",x"25",x"20"),
  1467 => (x"00",x"00",x"00",x"00"),
  1468 => (x"00",x"00",x"00",x"00"),
  1469 => (x"00",x"00",x"61",x"a8"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
