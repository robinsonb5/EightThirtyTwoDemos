
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"46",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"38"),
    10 => (x"41",x"98",x"27",x"4f"),
    11 => (x"27",x"4e",x"00",x"00"),
    12 => (x"00",x"00",x"06",x"22"),
    13 => (x"87",x"fd",x"00",x"0f"),
    14 => (x"4e",x"c0",x"f0",x"c1"),
    15 => (x"00",x"00",x"45",x"27"),
    16 => (x"fd",x"00",x"0f",x"00"),
    17 => (x"1e",x"4f",x"4f",x"87"),
    18 => (x"c0",x"ff",x"86",x"fc"),
    19 => (x"c4",x"48",x"69",x"49"),
    20 => (x"a6",x"c4",x"98",x"c0"),
    21 => (x"ff",x"02",x"6e",x"58"),
    22 => (x"66",x"c8",x"87",x"f3"),
    23 => (x"8e",x"fc",x"48",x"79"),
    24 => (x"5e",x"0e",x"4f",x"26"),
    25 => (x"cc",x"0e",x"5c",x"5b"),
    26 => (x"4c",x"c0",x"4b",x"66"),
    27 => (x"ff",x"c3",x"4a",x"13"),
    28 => (x"02",x"9a",x"72",x"9a"),
    29 => (x"72",x"87",x"d9",x"c0"),
    30 => (x"27",x"1e",x"71",x"49"),
    31 => (x"00",x"00",x"00",x"47"),
    32 => (x"c1",x"86",x"c4",x"0f"),
    33 => (x"c3",x"4a",x"13",x"84"),
    34 => (x"9a",x"72",x"9a",x"ff"),
    35 => (x"87",x"e7",x"ff",x"05"),
    36 => (x"4c",x"26",x"48",x"74"),
    37 => (x"4f",x"26",x"4b",x"26"),
    38 => (x"5c",x"5b",x"5e",x"0e"),
    39 => (x"66",x"d0",x"0e",x"5d"),
    40 => (x"16",x"e0",x"27",x"4a"),
    41 => (x"27",x"4b",x"00",x"00"),
    42 => (x"00",x"00",x"0f",x"28"),
    43 => (x"72",x"4c",x"c0",x"4d"),
    44 => (x"c6",x"c0",x"05",x"9a"),
    45 => (x"53",x"f0",x"c0",x"87"),
    46 => (x"72",x"87",x"f0",x"c0"),
    47 => (x"ea",x"c0",x"02",x"9a"),
    48 => (x"72",x"1e",x"72",x"87"),
    49 => (x"4a",x"66",x"d8",x"49"),
    50 => (x"00",x"05",x"a6",x"27"),
    51 => (x"4a",x"26",x"0f",x"00"),
    52 => (x"53",x"11",x"81",x"75"),
    53 => (x"49",x"72",x"1e",x"71"),
    54 => (x"27",x"4a",x"66",x"d8"),
    55 => (x"00",x"00",x"05",x"a6"),
    56 => (x"26",x"4a",x"70",x"0f"),
    57 => (x"05",x"9a",x"72",x"49"),
    58 => (x"27",x"87",x"d6",x"ff"),
    59 => (x"00",x"00",x"16",x"e0"),
    60 => (x"e1",x"c0",x"02",x"ab"),
    61 => (x"4d",x"66",x"d8",x"87"),
    62 => (x"c1",x"1e",x"66",x"dc"),
    63 => (x"49",x"6b",x"97",x"8b"),
    64 => (x"b9",x"81",x"c0",x"fe"),
    65 => (x"0f",x"75",x"1e",x"71"),
    66 => (x"84",x"c1",x"86",x"c8"),
    67 => (x"00",x"16",x"e0",x"27"),
    68 => (x"ff",x"05",x"ab",x"00"),
    69 => (x"48",x"74",x"87",x"e2"),
    70 => (x"4c",x"26",x"4d",x"26"),
    71 => (x"4f",x"26",x"4b",x"26"),
    72 => (x"5c",x"5b",x"5e",x"0e"),
    73 => (x"66",x"d0",x"0e",x"5d"),
    74 => (x"14",x"4d",x"ff",x"4c"),
    75 => (x"83",x"c0",x"fe",x"4b"),
    76 => (x"02",x"9b",x"73",x"bb"),
    77 => (x"c1",x"87",x"de",x"c0"),
    78 => (x"1e",x"66",x"d8",x"85"),
    79 => (x"66",x"dc",x"1e",x"73"),
    80 => (x"73",x"86",x"c8",x"0f"),
    81 => (x"cc",x"c0",x"05",x"a8"),
    82 => (x"fe",x"4b",x"14",x"87"),
    83 => (x"73",x"bb",x"83",x"c0"),
    84 => (x"e2",x"ff",x"05",x"9b"),
    85 => (x"26",x"48",x"75",x"87"),
    86 => (x"26",x"4c",x"26",x"4d"),
    87 => (x"0e",x"4f",x"26",x"4b"),
    88 => (x"5d",x"5c",x"5b",x"5e"),
    89 => (x"c0",x"86",x"f4",x"0e"),
    90 => (x"c0",x"4b",x"66",x"e4"),
    91 => (x"48",x"a6",x"c4",x"4c"),
    92 => (x"66",x"dc",x"78",x"c0"),
    93 => (x"fe",x"4d",x"bf",x"97"),
    94 => (x"dc",x"bd",x"85",x"c0"),
    95 => (x"80",x"c1",x"48",x"66"),
    96 => (x"58",x"a6",x"e0",x"c0"),
    97 => (x"c5",x"02",x"9d",x"75"),
    98 => (x"66",x"c4",x"87",x"c3"),
    99 => (x"87",x"cc",x"c4",x"02"),
   100 => (x"c0",x"48",x"a6",x"c8"),
   101 => (x"48",x"a6",x"c4",x"78"),
   102 => (x"49",x"75",x"78",x"c0"),
   103 => (x"02",x"ad",x"f0",x"c0"),
   104 => (x"c1",x"87",x"e7",x"c1"),
   105 => (x"c1",x"02",x"a9",x"e3"),
   106 => (x"e4",x"c1",x"87",x"e8"),
   107 => (x"e6",x"c0",x"02",x"a9"),
   108 => (x"a9",x"ec",x"c1",x"87"),
   109 => (x"87",x"d2",x"c1",x"02"),
   110 => (x"02",x"a9",x"f0",x"c1"),
   111 => (x"c1",x"87",x"e0",x"c0"),
   112 => (x"c0",x"02",x"a9",x"f3"),
   113 => (x"f5",x"c1",x"87",x"e1"),
   114 => (x"ca",x"c0",x"02",x"a9"),
   115 => (x"a9",x"f8",x"c1",x"87"),
   116 => (x"87",x"cb",x"c0",x"02"),
   117 => (x"c8",x"87",x"da",x"c1"),
   118 => (x"78",x"ca",x"48",x"a6"),
   119 => (x"c8",x"87",x"e9",x"c1"),
   120 => (x"78",x"d0",x"48",x"a6"),
   121 => (x"c0",x"87",x"e1",x"c1"),
   122 => (x"73",x"1e",x"66",x"e8"),
   123 => (x"66",x"e8",x"c0",x"1e"),
   124 => (x"c0",x"80",x"c4",x"48"),
   125 => (x"c0",x"58",x"a6",x"ec"),
   126 => (x"c4",x"49",x"66",x"e8"),
   127 => (x"fc",x"1e",x"69",x"89"),
   128 => (x"86",x"cc",x"87",x"de"),
   129 => (x"c0",x"84",x"49",x"70"),
   130 => (x"a6",x"c4",x"87",x"fe"),
   131 => (x"c0",x"78",x"c1",x"48"),
   132 => (x"e8",x"c0",x"87",x"f6"),
   133 => (x"e4",x"c0",x"1e",x"66"),
   134 => (x"80",x"c4",x"48",x"66"),
   135 => (x"58",x"a6",x"e8",x"c0"),
   136 => (x"49",x"66",x"e4",x"c0"),
   137 => (x"1e",x"69",x"89",x"c4"),
   138 => (x"86",x"c8",x"0f",x"73"),
   139 => (x"d7",x"c0",x"84",x"c1"),
   140 => (x"66",x"e8",x"c0",x"87"),
   141 => (x"1e",x"e5",x"c0",x"1e"),
   142 => (x"86",x"c8",x"0f",x"73"),
   143 => (x"1e",x"66",x"e8",x"c0"),
   144 => (x"0f",x"73",x"1e",x"75"),
   145 => (x"84",x"c1",x"86",x"c8"),
   146 => (x"c1",x"02",x"66",x"c8"),
   147 => (x"e0",x"c0",x"87",x"e7"),
   148 => (x"80",x"c4",x"48",x"66"),
   149 => (x"58",x"a6",x"e4",x"c0"),
   150 => (x"49",x"66",x"e0",x"c0"),
   151 => (x"48",x"76",x"89",x"c4"),
   152 => (x"e4",x"c1",x"78",x"69"),
   153 => (x"dc",x"c0",x"05",x"ad"),
   154 => (x"c0",x"48",x"6e",x"87"),
   155 => (x"c0",x"03",x"a8",x"b7"),
   156 => (x"ed",x"c0",x"87",x"d3"),
   157 => (x"00",x"47",x"27",x"1e"),
   158 => (x"c4",x"0f",x"00",x"00"),
   159 => (x"c0",x"48",x"6e",x"86"),
   160 => (x"a6",x"c4",x"88",x"08"),
   161 => (x"66",x"e8",x"c0",x"58"),
   162 => (x"d0",x"1e",x"73",x"1e"),
   163 => (x"66",x"cc",x"1e",x"66"),
   164 => (x"87",x"c4",x"f8",x"1e"),
   165 => (x"49",x"70",x"86",x"d0"),
   166 => (x"87",x"d9",x"c0",x"84"),
   167 => (x"05",x"ad",x"e5",x"c0"),
   168 => (x"c4",x"87",x"c8",x"c0"),
   169 => (x"78",x"c1",x"48",x"a6"),
   170 => (x"c0",x"87",x"ca",x"c0"),
   171 => (x"75",x"1e",x"66",x"e8"),
   172 => (x"c8",x"0f",x"73",x"1e"),
   173 => (x"97",x"66",x"dc",x"86"),
   174 => (x"c0",x"fe",x"4d",x"bf"),
   175 => (x"66",x"dc",x"bd",x"85"),
   176 => (x"c0",x"80",x"c1",x"48"),
   177 => (x"75",x"58",x"a6",x"e0"),
   178 => (x"fd",x"fa",x"05",x"9d"),
   179 => (x"f4",x"48",x"74",x"87"),
   180 => (x"26",x"4d",x"26",x"8e"),
   181 => (x"26",x"4b",x"26",x"4c"),
   182 => (x"1e",x"c0",x"1e",x"4f"),
   183 => (x"00",x"00",x"47",x"27"),
   184 => (x"66",x"d0",x"1e",x"00"),
   185 => (x"1e",x"66",x"d0",x"1e"),
   186 => (x"00",x"01",x"5f",x"27"),
   187 => (x"86",x"d0",x"0f",x"00"),
   188 => (x"c0",x"1e",x"4f",x"26"),
   189 => (x"00",x"47",x"27",x"1e"),
   190 => (x"d0",x"1e",x"00",x"00"),
   191 => (x"66",x"d0",x"1e",x"a6"),
   192 => (x"01",x"5f",x"27",x"1e"),
   193 => (x"d0",x"0f",x"00",x"00"),
   194 => (x"1e",x"4f",x"26",x"86"),
   195 => (x"49",x"4a",x"66",x"c8"),
   196 => (x"02",x"69",x"81",x"c4"),
   197 => (x"72",x"87",x"df",x"c0"),
   198 => (x"69",x"81",x"c4",x"49"),
   199 => (x"70",x"88",x"c1",x"48"),
   200 => (x"71",x"49",x"6a",x"79"),
   201 => (x"70",x"80",x"c1",x"48"),
   202 => (x"66",x"c4",x"97",x"7a"),
   203 => (x"98",x"ff",x"c3",x"51"),
   204 => (x"c0",x"48",x"66",x"c4"),
   205 => (x"48",x"c0",x"87",x"c2"),
   206 => (x"f8",x"1e",x"4f",x"26"),
   207 => (x"cc",x"48",x"76",x"86"),
   208 => (x"a6",x"c4",x"78",x"66"),
   209 => (x"76",x"78",x"ff",x"48"),
   210 => (x"03",x"0b",x"27",x"1e"),
   211 => (x"dc",x"1e",x"00",x"00"),
   212 => (x"66",x"dc",x"1e",x"a6"),
   213 => (x"01",x"5f",x"27",x"1e"),
   214 => (x"d0",x"0f",x"00",x"00"),
   215 => (x"26",x"8e",x"f8",x"86"),
   216 => (x"86",x"f8",x"1e",x"4f"),
   217 => (x"66",x"cc",x"48",x"76"),
   218 => (x"48",x"a6",x"c4",x"78"),
   219 => (x"76",x"78",x"66",x"d0"),
   220 => (x"03",x"0b",x"27",x"1e"),
   221 => (x"c0",x"1e",x"00",x"00"),
   222 => (x"c0",x"1e",x"a6",x"e0"),
   223 => (x"27",x"1e",x"66",x"e0"),
   224 => (x"00",x"00",x"01",x"5f"),
   225 => (x"f8",x"86",x"d0",x"0f"),
   226 => (x"1e",x"4f",x"26",x"8e"),
   227 => (x"48",x"76",x"86",x"f8"),
   228 => (x"c4",x"78",x"66",x"cc"),
   229 => (x"78",x"ff",x"48",x"a6"),
   230 => (x"0b",x"27",x"1e",x"76"),
   231 => (x"1e",x"00",x"00",x"03"),
   232 => (x"dc",x"1e",x"66",x"dc"),
   233 => (x"5f",x"27",x"1e",x"66"),
   234 => (x"0f",x"00",x"00",x"01"),
   235 => (x"8e",x"f8",x"86",x"d0"),
   236 => (x"73",x"1e",x"4f",x"26"),
   237 => (x"4b",x"66",x"cc",x"1e"),
   238 => (x"1e",x"7b",x"66",x"c8"),
   239 => (x"00",x"05",x"93",x"27"),
   240 => (x"86",x"c4",x"0f",x"00"),
   241 => (x"c0",x"05",x"98",x"70"),
   242 => (x"7b",x"c3",x"87",x"c2"),
   243 => (x"48",x"49",x"66",x"c8"),
   244 => (x"c0",x"02",x"a8",x"c0"),
   245 => (x"a9",x"c1",x"87",x"db"),
   246 => (x"87",x"da",x"c0",x"02"),
   247 => (x"c0",x"02",x"a9",x"c2"),
   248 => (x"a9",x"c3",x"87",x"ed"),
   249 => (x"87",x"ee",x"c0",x"02"),
   250 => (x"c0",x"02",x"a9",x"c4"),
   251 => (x"e5",x"c0",x"87",x"e6"),
   252 => (x"c0",x"7b",x"c0",x"87"),
   253 => (x"f8",x"27",x"87",x"e0"),
   254 => (x"bf",x"00",x"00",x"16"),
   255 => (x"b7",x"e4",x"c1",x"48"),
   256 => (x"c5",x"c0",x"06",x"a8"),
   257 => (x"c0",x"7b",x"c0",x"87"),
   258 => (x"7b",x"c3",x"87",x"cc"),
   259 => (x"c1",x"87",x"c7",x"c0"),
   260 => (x"87",x"c2",x"c0",x"7b"),
   261 => (x"4b",x"26",x"7b",x"c2"),
   262 => (x"c4",x"1e",x"4f",x"26"),
   263 => (x"81",x"c2",x"49",x"66"),
   264 => (x"71",x"48",x"66",x"c8"),
   265 => (x"08",x"66",x"cc",x"80"),
   266 => (x"4f",x"26",x"08",x"78"),
   267 => (x"5c",x"5b",x"5e",x"0e"),
   268 => (x"66",x"d8",x"0e",x"5d"),
   269 => (x"74",x"84",x"c5",x"4c"),
   270 => (x"93",x"b7",x"c4",x"4b"),
   271 => (x"dc",x"83",x"66",x"d0"),
   272 => (x"49",x"74",x"7b",x"66"),
   273 => (x"4a",x"71",x"81",x"c1"),
   274 => (x"d0",x"92",x"b7",x"c4"),
   275 => (x"7a",x"6b",x"82",x"66"),
   276 => (x"82",x"de",x"4a",x"74"),
   277 => (x"d0",x"92",x"b7",x"c4"),
   278 => (x"7a",x"74",x"82",x"66"),
   279 => (x"ac",x"b7",x"71",x"4d"),
   280 => (x"87",x"df",x"c0",x"01"),
   281 => (x"c8",x"c3",x"4a",x"74"),
   282 => (x"66",x"d4",x"92",x"b7"),
   283 => (x"c4",x"49",x"75",x"82"),
   284 => (x"81",x"72",x"91",x"b7"),
   285 => (x"85",x"c1",x"79",x"74"),
   286 => (x"81",x"c1",x"49",x"74"),
   287 => (x"06",x"ad",x"b7",x"71"),
   288 => (x"74",x"87",x"e1",x"ff"),
   289 => (x"b7",x"c8",x"c3",x"4a"),
   290 => (x"82",x"66",x"d4",x"92"),
   291 => (x"89",x"c1",x"49",x"74"),
   292 => (x"72",x"91",x"b7",x"c4"),
   293 => (x"c1",x"48",x"69",x"81"),
   294 => (x"74",x"79",x"70",x"80"),
   295 => (x"91",x"b7",x"c4",x"49"),
   296 => (x"71",x"4a",x"66",x"d0"),
   297 => (x"d4",x"4b",x"74",x"82"),
   298 => (x"b7",x"c8",x"c3",x"83"),
   299 => (x"83",x"66",x"d4",x"93"),
   300 => (x"79",x"6a",x"81",x"73"),
   301 => (x"00",x"16",x"f8",x"27"),
   302 => (x"78",x"c5",x"48",x"00"),
   303 => (x"4c",x"26",x"4d",x"26"),
   304 => (x"4f",x"26",x"4b",x"26"),
   305 => (x"0e",x"5b",x"5e",x"0e"),
   306 => (x"4b",x"66",x"c8",x"97"),
   307 => (x"c0",x"fe",x"4a",x"73"),
   308 => (x"cc",x"97",x"ba",x"82"),
   309 => (x"c0",x"fe",x"49",x"66"),
   310 => (x"b7",x"71",x"b9",x"81"),
   311 => (x"c5",x"c0",x"02",x"aa"),
   312 => (x"c0",x"48",x"c0",x"87"),
   313 => (x"04",x"27",x"87",x"c9"),
   314 => (x"97",x"00",x"00",x"17"),
   315 => (x"26",x"48",x"c1",x"5b"),
   316 => (x"0e",x"4f",x"26",x"4b"),
   317 => (x"0e",x"5c",x"5b",x"5e"),
   318 => (x"6e",x"97",x"86",x"fc"),
   319 => (x"d4",x"4b",x"c2",x"4c"),
   320 => (x"81",x"c1",x"49",x"66"),
   321 => (x"69",x"97",x"81",x"73"),
   322 => (x"81",x"c0",x"fe",x"49"),
   323 => (x"d4",x"1e",x"71",x"b9"),
   324 => (x"81",x"73",x"49",x"66"),
   325 => (x"fe",x"49",x"69",x"97"),
   326 => (x"71",x"b9",x"81",x"c0"),
   327 => (x"04",x"c4",x"27",x"1e"),
   328 => (x"c8",x"0f",x"00",x"00"),
   329 => (x"05",x"98",x"70",x"86"),
   330 => (x"c1",x"87",x"c5",x"c0"),
   331 => (x"83",x"c1",x"4c",x"c1"),
   332 => (x"06",x"ab",x"b7",x"c2"),
   333 => (x"74",x"87",x"c8",x"ff"),
   334 => (x"81",x"c0",x"fe",x"49"),
   335 => (x"b7",x"d7",x"c1",x"b9"),
   336 => (x"d0",x"c0",x"04",x"a9"),
   337 => (x"fe",x"49",x"74",x"87"),
   338 => (x"c1",x"b9",x"81",x"c0"),
   339 => (x"03",x"a9",x"b7",x"da"),
   340 => (x"c7",x"87",x"c2",x"c0"),
   341 => (x"fe",x"49",x"74",x"4b"),
   342 => (x"c1",x"b9",x"81",x"c0"),
   343 => (x"c0",x"05",x"a9",x"d2"),
   344 => (x"48",x"c1",x"87",x"c5"),
   345 => (x"d0",x"87",x"e4",x"c0"),
   346 => (x"66",x"d4",x"4a",x"66"),
   347 => (x"06",x"0a",x"27",x"49"),
   348 => (x"c0",x"0f",x"00",x"00"),
   349 => (x"c0",x"06",x"a8",x"b7"),
   350 => (x"48",x"73",x"87",x"cf"),
   351 => (x"fc",x"27",x"80",x"c7"),
   352 => (x"58",x"00",x"00",x"16"),
   353 => (x"c2",x"c0",x"48",x"c1"),
   354 => (x"fc",x"48",x"c0",x"87"),
   355 => (x"26",x"4c",x"26",x"8e"),
   356 => (x"1e",x"4f",x"26",x"4b"),
   357 => (x"c2",x"48",x"66",x"c4"),
   358 => (x"c5",x"c0",x"05",x"a8"),
   359 => (x"c0",x"48",x"c1",x"87"),
   360 => (x"48",x"c0",x"87",x"c2"),
   361 => (x"73",x"1e",x"4f",x"26"),
   362 => (x"02",x"9a",x"72",x"1e"),
   363 => (x"48",x"c0",x"87",x"e7"),
   364 => (x"a9",x"72",x"4b",x"c1"),
   365 => (x"72",x"87",x"d1",x"06"),
   366 => (x"87",x"c9",x"06",x"82"),
   367 => (x"a9",x"72",x"83",x"73"),
   368 => (x"c3",x"87",x"f4",x"01"),
   369 => (x"3a",x"b2",x"c1",x"87"),
   370 => (x"89",x"03",x"a9",x"72"),
   371 => (x"c1",x"07",x"80",x"73"),
   372 => (x"f3",x"05",x"2b",x"2a"),
   373 => (x"26",x"4b",x"26",x"87"),
   374 => (x"1e",x"75",x"1e",x"4f"),
   375 => (x"b7",x"71",x"4d",x"c4"),
   376 => (x"b9",x"ff",x"04",x"a1"),
   377 => (x"bd",x"c3",x"81",x"c1"),
   378 => (x"a2",x"b7",x"72",x"07"),
   379 => (x"c1",x"ba",x"ff",x"04"),
   380 => (x"07",x"bd",x"c1",x"82"),
   381 => (x"c1",x"87",x"ef",x"fe"),
   382 => (x"b8",x"ff",x"04",x"2d"),
   383 => (x"2d",x"07",x"80",x"c1"),
   384 => (x"c1",x"b9",x"ff",x"04"),
   385 => (x"4d",x"26",x"07",x"81"),
   386 => (x"72",x"1e",x"4f",x"26"),
   387 => (x"11",x"48",x"12",x"1e"),
   388 => (x"88",x"87",x"c4",x"02"),
   389 => (x"26",x"87",x"f6",x"02"),
   390 => (x"1e",x"4f",x"26",x"4a"),
   391 => (x"48",x"bf",x"c8",x"ff"),
   392 => (x"5e",x"0e",x"4f",x"26"),
   393 => (x"0e",x"5d",x"5c",x"5b"),
   394 => (x"66",x"c4",x"86",x"f0"),
   395 => (x"16",x"f4",x"27",x"4b"),
   396 => (x"27",x"48",x"00",x"00"),
   397 => (x"00",x"00",x"3e",x"f8"),
   398 => (x"16",x"f0",x"27",x"78"),
   399 => (x"27",x"48",x"00",x"00"),
   400 => (x"00",x"00",x"3f",x"28"),
   401 => (x"3f",x"28",x"27",x"78"),
   402 => (x"27",x"48",x"00",x"00"),
   403 => (x"00",x"00",x"3e",x"f8"),
   404 => (x"3f",x"2c",x"27",x"78"),
   405 => (x"c0",x"48",x"00",x"00"),
   406 => (x"3f",x"30",x"27",x"78"),
   407 => (x"c2",x"48",x"00",x"00"),
   408 => (x"3f",x"34",x"27",x"78"),
   409 => (x"c0",x"48",x"00",x"00"),
   410 => (x"1e",x"71",x"78",x"e8"),
   411 => (x"00",x"3f",x"38",x"27"),
   412 => (x"b2",x"27",x"49",x"00"),
   413 => (x"48",x"00",x"00",x"10"),
   414 => (x"41",x"20",x"41",x"20"),
   415 => (x"41",x"20",x"41",x"20"),
   416 => (x"41",x"20",x"41",x"20"),
   417 => (x"51",x"10",x"41",x"20"),
   418 => (x"51",x"10",x"51",x"10"),
   419 => (x"1e",x"71",x"49",x"26"),
   420 => (x"00",x"3f",x"58",x"27"),
   421 => (x"d1",x"27",x"49",x"00"),
   422 => (x"48",x"00",x"00",x"10"),
   423 => (x"41",x"20",x"41",x"20"),
   424 => (x"41",x"20",x"41",x"20"),
   425 => (x"41",x"20",x"41",x"20"),
   426 => (x"51",x"10",x"41",x"20"),
   427 => (x"51",x"10",x"51",x"10"),
   428 => (x"2c",x"27",x"49",x"26"),
   429 => (x"48",x"00",x"00",x"1e"),
   430 => (x"f0",x"27",x"78",x"ca"),
   431 => (x"1e",x"00",x"00",x"10"),
   432 => (x"00",x"02",x"f2",x"27"),
   433 => (x"86",x"c4",x"0f",x"00"),
   434 => (x"00",x"10",x"f2",x"27"),
   435 => (x"f2",x"27",x"1e",x"00"),
   436 => (x"0f",x"00",x"00",x"02"),
   437 => (x"22",x"27",x"86",x"c4"),
   438 => (x"1e",x"00",x"00",x"11"),
   439 => (x"00",x"02",x"f2",x"27"),
   440 => (x"86",x"c4",x"0f",x"00"),
   441 => (x"00",x"16",x"d8",x"27"),
   442 => (x"c0",x"02",x"bf",x"00"),
   443 => (x"39",x"27",x"87",x"df"),
   444 => (x"1e",x"00",x"00",x"0f"),
   445 => (x"00",x"02",x"f2",x"27"),
   446 => (x"86",x"c4",x"0f",x"00"),
   447 => (x"00",x"0f",x"65",x"27"),
   448 => (x"f2",x"27",x"1e",x"00"),
   449 => (x"0f",x"00",x"00",x"02"),
   450 => (x"dc",x"c0",x"86",x"c4"),
   451 => (x"0f",x"67",x"27",x"87"),
   452 => (x"27",x"1e",x"00",x"00"),
   453 => (x"00",x"00",x"02",x"f2"),
   454 => (x"27",x"86",x"c4",x"0f"),
   455 => (x"00",x"00",x"0f",x"96"),
   456 => (x"02",x"f2",x"27",x"1e"),
   457 => (x"c4",x"0f",x"00",x"00"),
   458 => (x"16",x"dc",x"27",x"86"),
   459 => (x"1e",x"bf",x"00",x"00"),
   460 => (x"00",x"11",x"24",x"27"),
   461 => (x"f2",x"27",x"1e",x"00"),
   462 => (x"0f",x"00",x"00",x"02"),
   463 => (x"1b",x"27",x"86",x"c8"),
   464 => (x"0f",x"00",x"00",x"06"),
   465 => (x"00",x"3e",x"e4",x"27"),
   466 => (x"4c",x"c1",x"58",x"00"),
   467 => (x"00",x"16",x"dc",x"27"),
   468 => (x"c0",x"48",x"bf",x"00"),
   469 => (x"c5",x"06",x"a8",x"b7"),
   470 => (x"11",x"27",x"87",x"fe"),
   471 => (x"0f",x"00",x"00",x"0f"),
   472 => (x"00",x"0e",x"dc",x"27"),
   473 => (x"48",x"76",x"0f",x"00"),
   474 => (x"4b",x"c3",x"78",x"c2"),
   475 => (x"78",x"27",x"1e",x"71"),
   476 => (x"49",x"00",x"00",x"3f"),
   477 => (x"00",x"0f",x"b7",x"27"),
   478 => (x"41",x"20",x"48",x"00"),
   479 => (x"41",x"20",x"41",x"20"),
   480 => (x"41",x"20",x"41",x"20"),
   481 => (x"41",x"20",x"41",x"20"),
   482 => (x"51",x"10",x"51",x"10"),
   483 => (x"49",x"26",x"51",x"10"),
   484 => (x"c1",x"48",x"a6",x"c8"),
   485 => (x"3f",x"78",x"27",x"78"),
   486 => (x"27",x"1e",x"00",x"00"),
   487 => (x"00",x"00",x"3f",x"58"),
   488 => (x"04",x"f3",x"27",x"1e"),
   489 => (x"c8",x"0f",x"00",x"00"),
   490 => (x"05",x"98",x"70",x"86"),
   491 => (x"c1",x"87",x"c5",x"c0"),
   492 => (x"87",x"c2",x"c0",x"49"),
   493 => (x"00",x"27",x"49",x"c0"),
   494 => (x"59",x"00",x"00",x"17"),
   495 => (x"06",x"ab",x"b7",x"6e"),
   496 => (x"6e",x"87",x"ea",x"c0"),
   497 => (x"91",x"b7",x"c5",x"49"),
   498 => (x"88",x"73",x"48",x"71"),
   499 => (x"cc",x"58",x"a6",x"d0"),
   500 => (x"1e",x"73",x"1e",x"a6"),
   501 => (x"27",x"1e",x"66",x"c8"),
   502 => (x"00",x"00",x"04",x"1a"),
   503 => (x"6e",x"86",x"cc",x"0f"),
   504 => (x"c4",x"80",x"c1",x"48"),
   505 => (x"b7",x"6e",x"58",x"a6"),
   506 => (x"d6",x"ff",x"01",x"ab"),
   507 => (x"1e",x"66",x"cc",x"87"),
   508 => (x"27",x"1e",x"66",x"c4"),
   509 => (x"00",x"00",x"17",x"d0"),
   510 => (x"17",x"08",x"27",x"1e"),
   511 => (x"27",x"1e",x"00",x"00"),
   512 => (x"00",x"00",x"04",x"2c"),
   513 => (x"27",x"86",x"d0",x"0f"),
   514 => (x"00",x"00",x"16",x"f0"),
   515 => (x"bf",x"27",x"1e",x"bf"),
   516 => (x"0f",x"00",x"00",x"0d"),
   517 => (x"c1",x"c1",x"86",x"c4"),
   518 => (x"17",x"01",x"27",x"4d"),
   519 => (x"bf",x"97",x"00",x"00"),
   520 => (x"81",x"c0",x"fe",x"49"),
   521 => (x"b7",x"c1",x"c1",x"b9"),
   522 => (x"ee",x"c1",x"04",x"a9"),
   523 => (x"1e",x"c3",x"c1",x"87"),
   524 => (x"c0",x"fe",x"49",x"75"),
   525 => (x"1e",x"71",x"b9",x"81"),
   526 => (x"00",x"04",x"c4",x"27"),
   527 => (x"86",x"c8",x"0f",x"00"),
   528 => (x"05",x"a8",x"66",x"c8"),
   529 => (x"c8",x"87",x"f9",x"c0"),
   530 => (x"1e",x"c0",x"1e",x"a6"),
   531 => (x"00",x"03",x"b2",x"27"),
   532 => (x"86",x"c8",x"0f",x"00"),
   533 => (x"78",x"27",x"1e",x"71"),
   534 => (x"49",x"00",x"00",x"3f"),
   535 => (x"00",x"0f",x"98",x"27"),
   536 => (x"41",x"20",x"48",x"00"),
   537 => (x"41",x"20",x"41",x"20"),
   538 => (x"41",x"20",x"41",x"20"),
   539 => (x"41",x"20",x"41",x"20"),
   540 => (x"51",x"10",x"51",x"10"),
   541 => (x"49",x"26",x"51",x"10"),
   542 => (x"fc",x"27",x"4b",x"74"),
   543 => (x"5c",x"00",x"00",x"16"),
   544 => (x"4a",x"75",x"85",x"c1"),
   545 => (x"ba",x"82",x"c0",x"fe"),
   546 => (x"00",x"17",x"01",x"27"),
   547 => (x"49",x"bf",x"97",x"00"),
   548 => (x"b9",x"81",x"c0",x"fe"),
   549 => (x"06",x"aa",x"b7",x"71"),
   550 => (x"6e",x"87",x"d2",x"fe"),
   551 => (x"1e",x"71",x"93",x"b7"),
   552 => (x"49",x"73",x"1e",x"72"),
   553 => (x"27",x"4a",x"66",x"d4"),
   554 => (x"00",x"00",x"05",x"d9"),
   555 => (x"26",x"4a",x"26",x"0f"),
   556 => (x"58",x"a6",x"c4",x"49"),
   557 => (x"66",x"cc",x"49",x"73"),
   558 => (x"91",x"b7",x"c7",x"89"),
   559 => (x"8b",x"6e",x"4b",x"71"),
   560 => (x"5c",x"27",x"1e",x"76"),
   561 => (x"0f",x"00",x"00",x"0e"),
   562 => (x"84",x"c1",x"86",x"c4"),
   563 => (x"00",x"16",x"dc",x"27"),
   564 => (x"ac",x"b7",x"bf",x"00"),
   565 => (x"87",x"c2",x"fa",x"06"),
   566 => (x"00",x"06",x"1b",x"27"),
   567 => (x"e8",x"27",x"0f",x"00"),
   568 => (x"58",x"00",x"00",x"3e"),
   569 => (x"00",x"11",x"51",x"27"),
   570 => (x"f2",x"27",x"1e",x"00"),
   571 => (x"0f",x"00",x"00",x"02"),
   572 => (x"61",x"27",x"86",x"c4"),
   573 => (x"1e",x"00",x"00",x"11"),
   574 => (x"00",x"02",x"f2",x"27"),
   575 => (x"86",x"c4",x"0f",x"00"),
   576 => (x"00",x"11",x"63",x"27"),
   577 => (x"f2",x"27",x"1e",x"00"),
   578 => (x"0f",x"00",x"00",x"02"),
   579 => (x"99",x"27",x"86",x"c4"),
   580 => (x"1e",x"00",x"00",x"11"),
   581 => (x"00",x"02",x"f2",x"27"),
   582 => (x"86",x"c4",x"0f",x"00"),
   583 => (x"00",x"16",x"f8",x"27"),
   584 => (x"27",x"1e",x"bf",x"00"),
   585 => (x"00",x"00",x"11",x"9b"),
   586 => (x"02",x"f2",x"27",x"1e"),
   587 => (x"c8",x"0f",x"00",x"00"),
   588 => (x"27",x"1e",x"c5",x"86"),
   589 => (x"00",x"00",x"11",x"b4"),
   590 => (x"02",x"f2",x"27",x"1e"),
   591 => (x"c8",x"0f",x"00",x"00"),
   592 => (x"16",x"fc",x"27",x"86"),
   593 => (x"1e",x"bf",x"00",x"00"),
   594 => (x"00",x"11",x"cd",x"27"),
   595 => (x"f2",x"27",x"1e",x"00"),
   596 => (x"0f",x"00",x"00",x"02"),
   597 => (x"1e",x"c1",x"86",x"c8"),
   598 => (x"00",x"11",x"e6",x"27"),
   599 => (x"f2",x"27",x"1e",x"00"),
   600 => (x"0f",x"00",x"00",x"02"),
   601 => (x"00",x"27",x"86",x"c8"),
   602 => (x"97",x"00",x"00",x"17"),
   603 => (x"c0",x"fe",x"49",x"bf"),
   604 => (x"1e",x"71",x"b9",x"81"),
   605 => (x"00",x"11",x"ff",x"27"),
   606 => (x"f2",x"27",x"1e",x"00"),
   607 => (x"0f",x"00",x"00",x"02"),
   608 => (x"c1",x"c1",x"86",x"c8"),
   609 => (x"12",x"18",x"27",x"1e"),
   610 => (x"27",x"1e",x"00",x"00"),
   611 => (x"00",x"00",x"02",x"f2"),
   612 => (x"27",x"86",x"c8",x"0f"),
   613 => (x"00",x"00",x"17",x"01"),
   614 => (x"fe",x"49",x"bf",x"97"),
   615 => (x"71",x"b9",x"81",x"c0"),
   616 => (x"12",x"31",x"27",x"1e"),
   617 => (x"27",x"1e",x"00",x"00"),
   618 => (x"00",x"00",x"02",x"f2"),
   619 => (x"c1",x"86",x"c8",x"0f"),
   620 => (x"4a",x"27",x"1e",x"c2"),
   621 => (x"1e",x"00",x"00",x"12"),
   622 => (x"00",x"02",x"f2",x"27"),
   623 => (x"86",x"c8",x"0f",x"00"),
   624 => (x"00",x"17",x"28",x"27"),
   625 => (x"27",x"1e",x"bf",x"00"),
   626 => (x"00",x"00",x"12",x"63"),
   627 => (x"02",x"f2",x"27",x"1e"),
   628 => (x"c8",x"0f",x"00",x"00"),
   629 => (x"27",x"1e",x"c7",x"86"),
   630 => (x"00",x"00",x"12",x"7c"),
   631 => (x"02",x"f2",x"27",x"1e"),
   632 => (x"c8",x"0f",x"00",x"00"),
   633 => (x"1e",x"2c",x"27",x"86"),
   634 => (x"1e",x"bf",x"00",x"00"),
   635 => (x"00",x"12",x"95",x"27"),
   636 => (x"f2",x"27",x"1e",x"00"),
   637 => (x"0f",x"00",x"00",x"02"),
   638 => (x"ae",x"27",x"86",x"c8"),
   639 => (x"1e",x"00",x"00",x"12"),
   640 => (x"00",x"02",x"f2",x"27"),
   641 => (x"86",x"c4",x"0f",x"00"),
   642 => (x"00",x"12",x"d8",x"27"),
   643 => (x"f2",x"27",x"1e",x"00"),
   644 => (x"0f",x"00",x"00",x"02"),
   645 => (x"f0",x"27",x"86",x"c4"),
   646 => (x"bf",x"00",x"00",x"16"),
   647 => (x"e4",x"27",x"1e",x"bf"),
   648 => (x"1e",x"00",x"00",x"12"),
   649 => (x"00",x"02",x"f2",x"27"),
   650 => (x"86",x"c8",x"0f",x"00"),
   651 => (x"00",x"12",x"fd",x"27"),
   652 => (x"f2",x"27",x"1e",x"00"),
   653 => (x"0f",x"00",x"00",x"02"),
   654 => (x"f0",x"27",x"86",x"c4"),
   655 => (x"bf",x"00",x"00",x"16"),
   656 => (x"69",x"81",x"c4",x"49"),
   657 => (x"13",x"2e",x"27",x"1e"),
   658 => (x"27",x"1e",x"00",x"00"),
   659 => (x"00",x"00",x"02",x"f2"),
   660 => (x"c0",x"86",x"c8",x"0f"),
   661 => (x"13",x"47",x"27",x"1e"),
   662 => (x"27",x"1e",x"00",x"00"),
   663 => (x"00",x"00",x"02",x"f2"),
   664 => (x"27",x"86",x"c8",x"0f"),
   665 => (x"00",x"00",x"16",x"f0"),
   666 => (x"81",x"c8",x"49",x"bf"),
   667 => (x"60",x"27",x"1e",x"69"),
   668 => (x"1e",x"00",x"00",x"13"),
   669 => (x"00",x"02",x"f2",x"27"),
   670 => (x"86",x"c8",x"0f",x"00"),
   671 => (x"79",x"27",x"1e",x"c2"),
   672 => (x"1e",x"00",x"00",x"13"),
   673 => (x"00",x"02",x"f2",x"27"),
   674 => (x"86",x"c8",x"0f",x"00"),
   675 => (x"00",x"16",x"f0",x"27"),
   676 => (x"cc",x"49",x"bf",x"00"),
   677 => (x"27",x"1e",x"69",x"81"),
   678 => (x"00",x"00",x"13",x"92"),
   679 => (x"02",x"f2",x"27",x"1e"),
   680 => (x"c8",x"0f",x"00",x"00"),
   681 => (x"27",x"1e",x"d1",x"86"),
   682 => (x"00",x"00",x"13",x"ab"),
   683 => (x"02",x"f2",x"27",x"1e"),
   684 => (x"c8",x"0f",x"00",x"00"),
   685 => (x"16",x"f0",x"27",x"86"),
   686 => (x"49",x"bf",x"00",x"00"),
   687 => (x"1e",x"71",x"81",x"d0"),
   688 => (x"00",x"13",x"c4",x"27"),
   689 => (x"f2",x"27",x"1e",x"00"),
   690 => (x"0f",x"00",x"00",x"02"),
   691 => (x"dd",x"27",x"86",x"c8"),
   692 => (x"1e",x"00",x"00",x"13"),
   693 => (x"00",x"02",x"f2",x"27"),
   694 => (x"86",x"c4",x"0f",x"00"),
   695 => (x"00",x"14",x"12",x"27"),
   696 => (x"f2",x"27",x"1e",x"00"),
   697 => (x"0f",x"00",x"00",x"02"),
   698 => (x"f4",x"27",x"86",x"c4"),
   699 => (x"bf",x"00",x"00",x"16"),
   700 => (x"23",x"27",x"1e",x"bf"),
   701 => (x"1e",x"00",x"00",x"14"),
   702 => (x"00",x"02",x"f2",x"27"),
   703 => (x"86",x"c8",x"0f",x"00"),
   704 => (x"00",x"14",x"3c",x"27"),
   705 => (x"f2",x"27",x"1e",x"00"),
   706 => (x"0f",x"00",x"00",x"02"),
   707 => (x"f4",x"27",x"86",x"c4"),
   708 => (x"bf",x"00",x"00",x"16"),
   709 => (x"69",x"81",x"c4",x"49"),
   710 => (x"14",x"7c",x"27",x"1e"),
   711 => (x"27",x"1e",x"00",x"00"),
   712 => (x"00",x"00",x"02",x"f2"),
   713 => (x"c0",x"86",x"c8",x"0f"),
   714 => (x"14",x"95",x"27",x"1e"),
   715 => (x"27",x"1e",x"00",x"00"),
   716 => (x"00",x"00",x"02",x"f2"),
   717 => (x"27",x"86",x"c8",x"0f"),
   718 => (x"00",x"00",x"16",x"f4"),
   719 => (x"81",x"c8",x"49",x"bf"),
   720 => (x"ae",x"27",x"1e",x"69"),
   721 => (x"1e",x"00",x"00",x"14"),
   722 => (x"00",x"02",x"f2",x"27"),
   723 => (x"86",x"c8",x"0f",x"00"),
   724 => (x"c7",x"27",x"1e",x"c1"),
   725 => (x"1e",x"00",x"00",x"14"),
   726 => (x"00",x"02",x"f2",x"27"),
   727 => (x"86",x"c8",x"0f",x"00"),
   728 => (x"00",x"16",x"f4",x"27"),
   729 => (x"cc",x"49",x"bf",x"00"),
   730 => (x"27",x"1e",x"69",x"81"),
   731 => (x"00",x"00",x"14",x"e0"),
   732 => (x"02",x"f2",x"27",x"1e"),
   733 => (x"c8",x"0f",x"00",x"00"),
   734 => (x"27",x"1e",x"d2",x"86"),
   735 => (x"00",x"00",x"14",x"f9"),
   736 => (x"02",x"f2",x"27",x"1e"),
   737 => (x"c8",x"0f",x"00",x"00"),
   738 => (x"16",x"f4",x"27",x"86"),
   739 => (x"49",x"bf",x"00",x"00"),
   740 => (x"1e",x"71",x"81",x"d0"),
   741 => (x"00",x"15",x"12",x"27"),
   742 => (x"f2",x"27",x"1e",x"00"),
   743 => (x"0f",x"00",x"00",x"02"),
   744 => (x"2b",x"27",x"86",x"c8"),
   745 => (x"1e",x"00",x"00",x"15"),
   746 => (x"00",x"02",x"f2",x"27"),
   747 => (x"86",x"c4",x"0f",x"00"),
   748 => (x"60",x"27",x"1e",x"6e"),
   749 => (x"1e",x"00",x"00",x"15"),
   750 => (x"00",x"02",x"f2",x"27"),
   751 => (x"86",x"c8",x"0f",x"00"),
   752 => (x"79",x"27",x"1e",x"c5"),
   753 => (x"1e",x"00",x"00",x"15"),
   754 => (x"00",x"02",x"f2",x"27"),
   755 => (x"86",x"c8",x"0f",x"00"),
   756 => (x"92",x"27",x"1e",x"73"),
   757 => (x"1e",x"00",x"00",x"15"),
   758 => (x"00",x"02",x"f2",x"27"),
   759 => (x"86",x"c8",x"0f",x"00"),
   760 => (x"ab",x"27",x"1e",x"cd"),
   761 => (x"1e",x"00",x"00",x"15"),
   762 => (x"00",x"02",x"f2",x"27"),
   763 => (x"86",x"c8",x"0f",x"00"),
   764 => (x"27",x"1e",x"66",x"cc"),
   765 => (x"00",x"00",x"15",x"c4"),
   766 => (x"02",x"f2",x"27",x"1e"),
   767 => (x"c8",x"0f",x"00",x"00"),
   768 => (x"27",x"1e",x"c7",x"86"),
   769 => (x"00",x"00",x"15",x"dd"),
   770 => (x"02",x"f2",x"27",x"1e"),
   771 => (x"c8",x"0f",x"00",x"00"),
   772 => (x"1e",x"66",x"c8",x"86"),
   773 => (x"00",x"15",x"f6",x"27"),
   774 => (x"f2",x"27",x"1e",x"00"),
   775 => (x"0f",x"00",x"00",x"02"),
   776 => (x"1e",x"c1",x"86",x"c8"),
   777 => (x"00",x"16",x"0f",x"27"),
   778 => (x"f2",x"27",x"1e",x"00"),
   779 => (x"0f",x"00",x"00",x"02"),
   780 => (x"58",x"27",x"86",x"c8"),
   781 => (x"1e",x"00",x"00",x"3f"),
   782 => (x"00",x"16",x"28",x"27"),
   783 => (x"f2",x"27",x"1e",x"00"),
   784 => (x"0f",x"00",x"00",x"02"),
   785 => (x"41",x"27",x"86",x"c8"),
   786 => (x"1e",x"00",x"00",x"16"),
   787 => (x"00",x"02",x"f2",x"27"),
   788 => (x"86",x"c4",x"0f",x"00"),
   789 => (x"00",x"3f",x"78",x"27"),
   790 => (x"76",x"27",x"1e",x"00"),
   791 => (x"1e",x"00",x"00",x"16"),
   792 => (x"00",x"02",x"f2",x"27"),
   793 => (x"86",x"c8",x"0f",x"00"),
   794 => (x"00",x"16",x"8f",x"27"),
   795 => (x"f2",x"27",x"1e",x"00"),
   796 => (x"0f",x"00",x"00",x"02"),
   797 => (x"c4",x"27",x"86",x"c4"),
   798 => (x"1e",x"00",x"00",x"16"),
   799 => (x"00",x"02",x"f2",x"27"),
   800 => (x"86",x"c4",x"0f",x"00"),
   801 => (x"00",x"3e",x"e4",x"27"),
   802 => (x"27",x"49",x"bf",x"00"),
   803 => (x"00",x"00",x"3e",x"e0"),
   804 => (x"ec",x"27",x"89",x"bf"),
   805 => (x"59",x"00",x"00",x"3e"),
   806 => (x"c6",x"27",x"1e",x"71"),
   807 => (x"1e",x"00",x"00",x"16"),
   808 => (x"00",x"02",x"f2",x"27"),
   809 => (x"86",x"c8",x"0f",x"00"),
   810 => (x"00",x"3e",x"e8",x"27"),
   811 => (x"c1",x"48",x"bf",x"00"),
   812 => (x"03",x"a8",x"b7",x"f8"),
   813 => (x"27",x"87",x"ea",x"c0"),
   814 => (x"00",x"00",x"0f",x"d6"),
   815 => (x"02",x"f2",x"27",x"1e"),
   816 => (x"c4",x"0f",x"00",x"00"),
   817 => (x"10",x"0c",x"27",x"86"),
   818 => (x"27",x"1e",x"00",x"00"),
   819 => (x"00",x"00",x"02",x"f2"),
   820 => (x"27",x"86",x"c4",x"0f"),
   821 => (x"00",x"00",x"10",x"2c"),
   822 => (x"02",x"f2",x"27",x"1e"),
   823 => (x"c4",x"0f",x"00",x"00"),
   824 => (x"3e",x"e8",x"27",x"86"),
   825 => (x"49",x"bf",x"00",x"00"),
   826 => (x"e8",x"cf",x"4a",x"71"),
   827 => (x"1e",x"71",x"92",x"b7"),
   828 => (x"49",x"72",x"1e",x"72"),
   829 => (x"00",x"16",x"dc",x"27"),
   830 => (x"27",x"4a",x"bf",x"00"),
   831 => (x"00",x"00",x"05",x"d9"),
   832 => (x"26",x"4a",x"26",x"0f"),
   833 => (x"3e",x"f0",x"27",x"49"),
   834 => (x"27",x"58",x"00",x"00"),
   835 => (x"00",x"00",x"16",x"dc"),
   836 => (x"4b",x"72",x"4a",x"bf"),
   837 => (x"93",x"b7",x"e8",x"cf"),
   838 => (x"1e",x"72",x"1e",x"71"),
   839 => (x"27",x"4a",x"09",x"73"),
   840 => (x"00",x"00",x"05",x"d9"),
   841 => (x"26",x"4a",x"26",x"0f"),
   842 => (x"3e",x"f4",x"27",x"49"),
   843 => (x"c8",x"58",x"00",x"00"),
   844 => (x"71",x"92",x"b7",x"f9"),
   845 => (x"72",x"1e",x"72",x"1e"),
   846 => (x"d9",x"27",x"4a",x"09"),
   847 => (x"0f",x"00",x"00",x"05"),
   848 => (x"49",x"26",x"4a",x"26"),
   849 => (x"00",x"3e",x"f8",x"27"),
   850 => (x"2e",x"27",x"58",x"00"),
   851 => (x"1e",x"00",x"00",x"10"),
   852 => (x"00",x"02",x"f2",x"27"),
   853 => (x"86",x"c4",x"0f",x"00"),
   854 => (x"00",x"3e",x"ec",x"27"),
   855 => (x"27",x"1e",x"bf",x"00"),
   856 => (x"00",x"00",x"10",x"5b"),
   857 => (x"02",x"f2",x"27",x"1e"),
   858 => (x"c8",x"0f",x"00",x"00"),
   859 => (x"10",x"60",x"27",x"86"),
   860 => (x"27",x"1e",x"00",x"00"),
   861 => (x"00",x"00",x"02",x"f2"),
   862 => (x"27",x"86",x"c4",x"0f"),
   863 => (x"00",x"00",x"3e",x"f0"),
   864 => (x"8d",x"27",x"1e",x"bf"),
   865 => (x"1e",x"00",x"00",x"10"),
   866 => (x"00",x"02",x"f2",x"27"),
   867 => (x"86",x"c8",x"0f",x"00"),
   868 => (x"00",x"3e",x"f4",x"27"),
   869 => (x"27",x"1e",x"bf",x"00"),
   870 => (x"00",x"00",x"10",x"92"),
   871 => (x"02",x"f2",x"27",x"1e"),
   872 => (x"c8",x"0f",x"00",x"00"),
   873 => (x"10",x"b0",x"27",x"86"),
   874 => (x"27",x"1e",x"00",x"00"),
   875 => (x"00",x"00",x"02",x"f2"),
   876 => (x"c0",x"86",x"c4",x"0f"),
   877 => (x"26",x"8e",x"f0",x"48"),
   878 => (x"26",x"4c",x"26",x"4d"),
   879 => (x"0e",x"4f",x"26",x"4b"),
   880 => (x"5d",x"5c",x"5b",x"5e"),
   881 => (x"4d",x"66",x"d0",x"0e"),
   882 => (x"4c",x"73",x"4b",x"6d"),
   883 => (x"1e",x"72",x"1e",x"71"),
   884 => (x"f0",x"27",x"49",x"73"),
   885 => (x"bf",x"00",x"00",x"16"),
   886 => (x"a1",x"f0",x"c0",x"48"),
   887 => (x"71",x"41",x"20",x"4a"),
   888 => (x"87",x"f9",x"05",x"aa"),
   889 => (x"49",x"26",x"4a",x"26"),
   890 => (x"82",x"cc",x"4a",x"75"),
   891 => (x"49",x"73",x"7a",x"c5"),
   892 => (x"79",x"6a",x"81",x"cc"),
   893 => (x"1e",x"73",x"7b",x"6d"),
   894 => (x"00",x"0e",x"a8",x"27"),
   895 => (x"86",x"c4",x"0f",x"00"),
   896 => (x"81",x"c4",x"49",x"73"),
   897 => (x"f3",x"c0",x"05",x"69"),
   898 => (x"c8",x"49",x"74",x"87"),
   899 => (x"cc",x"4b",x"74",x"81"),
   900 => (x"71",x"7b",x"c6",x"83"),
   901 => (x"c8",x"49",x"75",x"1e"),
   902 => (x"27",x"1e",x"69",x"81"),
   903 => (x"00",x"00",x"03",x"b2"),
   904 => (x"27",x"86",x"c8",x"0f"),
   905 => (x"00",x"00",x"16",x"f0"),
   906 => (x"73",x"7c",x"bf",x"bf"),
   907 => (x"6b",x"1e",x"ca",x"1e"),
   908 => (x"04",x"1a",x"27",x"1e"),
   909 => (x"cc",x"0f",x"00",x"00"),
   910 => (x"87",x"d8",x"c0",x"86"),
   911 => (x"1e",x"71",x"49",x"6d"),
   912 => (x"49",x"75",x"1e",x"72"),
   913 => (x"a1",x"f0",x"c0",x"48"),
   914 => (x"71",x"41",x"20",x"4a"),
   915 => (x"87",x"f9",x"05",x"aa"),
   916 => (x"49",x"26",x"4a",x"26"),
   917 => (x"4c",x"26",x"4d",x"26"),
   918 => (x"4f",x"26",x"4b",x"26"),
   919 => (x"5c",x"5b",x"5e",x"0e"),
   920 => (x"86",x"fc",x"0e",x"5d"),
   921 => (x"00",x"17",x"00",x"27"),
   922 => (x"4d",x"bf",x"97",x"00"),
   923 => (x"66",x"d4",x"4c",x"6e"),
   924 => (x"ca",x"4a",x"6b",x"4b"),
   925 => (x"fe",x"49",x"75",x"82"),
   926 => (x"c1",x"b9",x"81",x"c0"),
   927 => (x"c0",x"05",x"a9",x"c1"),
   928 => (x"8a",x"c1",x"87",x"cf"),
   929 => (x"f8",x"27",x"48",x"72"),
   930 => (x"bf",x"00",x"00",x"16"),
   931 => (x"c0",x"7b",x"70",x"88"),
   932 => (x"05",x"9c",x"74",x"4c"),
   933 => (x"27",x"87",x"de",x"ff"),
   934 => (x"00",x"00",x"17",x"04"),
   935 => (x"8e",x"fc",x"5d",x"97"),
   936 => (x"4c",x"26",x"4d",x"26"),
   937 => (x"4f",x"26",x"4b",x"26"),
   938 => (x"16",x"f0",x"27",x"1e"),
   939 => (x"02",x"bf",x"00",x"00"),
   940 => (x"c4",x"87",x"cb",x"c0"),
   941 => (x"f0",x"27",x"48",x"66"),
   942 => (x"bf",x"00",x"00",x"16"),
   943 => (x"f0",x"27",x"78",x"bf"),
   944 => (x"bf",x"00",x"00",x"16"),
   945 => (x"71",x"81",x"cc",x"49"),
   946 => (x"16",x"f8",x"27",x"1e"),
   947 => (x"1e",x"bf",x"00",x"00"),
   948 => (x"1a",x"27",x"1e",x"ca"),
   949 => (x"0f",x"00",x"00",x"04"),
   950 => (x"4f",x"26",x"86",x"cc"),
   951 => (x"17",x"00",x"27",x"1e"),
   952 => (x"bf",x"97",x"00",x"00"),
   953 => (x"81",x"c0",x"fe",x"49"),
   954 => (x"a9",x"c1",x"c1",x"b9"),
   955 => (x"87",x"c5",x"c0",x"02"),
   956 => (x"c2",x"c0",x"49",x"c0"),
   957 => (x"27",x"49",x"c1",x"87"),
   958 => (x"00",x"00",x"16",x"fc"),
   959 => (x"b0",x"71",x"48",x"bf"),
   960 => (x"00",x"17",x"00",x"27"),
   961 => (x"01",x"27",x"58",x"00"),
   962 => (x"48",x"00",x"00",x"17"),
   963 => (x"26",x"50",x"c2",x"c1"),
   964 => (x"00",x"27",x"1e",x"4f"),
   965 => (x"48",x"00",x"00",x"17"),
   966 => (x"27",x"50",x"c1",x"c1"),
   967 => (x"00",x"00",x"16",x"fc"),
   968 => (x"26",x"78",x"c0",x"48"),
   969 => (x"00",x"00",x"00",x"4f"),
   970 => (x"33",x"32",x"31",x"30"),
   971 => (x"37",x"36",x"35",x"34"),
   972 => (x"42",x"41",x"39",x"38"),
   973 => (x"46",x"45",x"44",x"43"),
   974 => (x"6f",x"72",x"50",x"00"),
   975 => (x"6d",x"61",x"72",x"67"),
   976 => (x"6d",x"6f",x"63",x"20"),
   977 => (x"65",x"6c",x"69",x"70"),
   978 => (x"69",x"77",x"20",x"64"),
   979 => (x"27",x"20",x"68",x"74"),
   980 => (x"69",x"67",x"65",x"72"),
   981 => (x"72",x"65",x"74",x"73"),
   982 => (x"74",x"61",x"20",x"27"),
   983 => (x"62",x"69",x"72",x"74"),
   984 => (x"0a",x"65",x"74",x"75"),
   985 => (x"50",x"00",x"0a",x"00"),
   986 => (x"72",x"67",x"6f",x"72"),
   987 => (x"63",x"20",x"6d",x"61"),
   988 => (x"69",x"70",x"6d",x"6f"),
   989 => (x"20",x"64",x"65",x"6c"),
   990 => (x"68",x"74",x"69",x"77"),
   991 => (x"20",x"74",x"75",x"6f"),
   992 => (x"67",x"65",x"72",x"27"),
   993 => (x"65",x"74",x"73",x"69"),
   994 => (x"61",x"20",x"27",x"72"),
   995 => (x"69",x"72",x"74",x"74"),
   996 => (x"65",x"74",x"75",x"62"),
   997 => (x"00",x"0a",x"00",x"0a"),
   998 => (x"59",x"52",x"48",x"44"),
   999 => (x"4e",x"4f",x"54",x"53"),
  1000 => (x"52",x"50",x"20",x"45"),
  1001 => (x"41",x"52",x"47",x"4f"),
  1002 => (x"33",x"20",x"2c",x"4d"),
  1003 => (x"20",x"44",x"52",x"27"),
  1004 => (x"49",x"52",x"54",x"53"),
  1005 => (x"44",x"00",x"47",x"4e"),
  1006 => (x"53",x"59",x"52",x"48"),
  1007 => (x"45",x"4e",x"4f",x"54"),
  1008 => (x"4f",x"52",x"50",x"20"),
  1009 => (x"4d",x"41",x"52",x"47"),
  1010 => (x"27",x"32",x"20",x"2c"),
  1011 => (x"53",x"20",x"44",x"4e"),
  1012 => (x"4e",x"49",x"52",x"54"),
  1013 => (x"65",x"4d",x"00",x"47"),
  1014 => (x"72",x"75",x"73",x"61"),
  1015 => (x"74",x"20",x"64",x"65"),
  1016 => (x"20",x"65",x"6d",x"69"),
  1017 => (x"20",x"6f",x"6f",x"74"),
  1018 => (x"6c",x"61",x"6d",x"73"),
  1019 => (x"6f",x"74",x"20",x"6c"),
  1020 => (x"74",x"62",x"6f",x"20"),
  1021 => (x"20",x"6e",x"69",x"61"),
  1022 => (x"6e",x"61",x"65",x"6d"),
  1023 => (x"66",x"67",x"6e",x"69"),
  1024 => (x"72",x"20",x"6c",x"75"),
  1025 => (x"6c",x"75",x"73",x"65"),
  1026 => (x"00",x"0a",x"73",x"74"),
  1027 => (x"61",x"65",x"6c",x"50"),
  1028 => (x"69",x"20",x"65",x"73"),
  1029 => (x"65",x"72",x"63",x"6e"),
  1030 => (x"20",x"65",x"73",x"61"),
  1031 => (x"62",x"6d",x"75",x"6e"),
  1032 => (x"6f",x"20",x"72",x"65"),
  1033 => (x"75",x"72",x"20",x"66"),
  1034 => (x"00",x"0a",x"73",x"6e"),
  1035 => (x"69",x"4d",x"00",x"0a"),
  1036 => (x"73",x"6f",x"72",x"63"),
  1037 => (x"6e",x"6f",x"63",x"65"),
  1038 => (x"66",x"20",x"73",x"64"),
  1039 => (x"6f",x"20",x"72",x"6f"),
  1040 => (x"72",x"20",x"65",x"6e"),
  1041 => (x"74",x"20",x"6e",x"75"),
  1042 => (x"75",x"6f",x"72",x"68"),
  1043 => (x"44",x"20",x"68",x"67"),
  1044 => (x"73",x"79",x"72",x"68"),
  1045 => (x"65",x"6e",x"6f",x"74"),
  1046 => (x"25",x"00",x"20",x"3a"),
  1047 => (x"00",x"0a",x"20",x"64"),
  1048 => (x"79",x"72",x"68",x"44"),
  1049 => (x"6e",x"6f",x"74",x"73"),
  1050 => (x"70",x"20",x"73",x"65"),
  1051 => (x"53",x"20",x"72",x"65"),
  1052 => (x"6e",x"6f",x"63",x"65"),
  1053 => (x"20",x"20",x"3a",x"64"),
  1054 => (x"20",x"20",x"20",x"20"),
  1055 => (x"20",x"20",x"20",x"20"),
  1056 => (x"20",x"20",x"20",x"20"),
  1057 => (x"20",x"20",x"20",x"20"),
  1058 => (x"20",x"20",x"20",x"20"),
  1059 => (x"20",x"64",x"25",x"00"),
  1060 => (x"41",x"56",x"00",x"0a"),
  1061 => (x"49",x"4d",x"20",x"58"),
  1062 => (x"72",x"20",x"53",x"50"),
  1063 => (x"6e",x"69",x"74",x"61"),
  1064 => (x"20",x"2a",x"20",x"67"),
  1065 => (x"30",x"30",x"30",x"31"),
  1066 => (x"25",x"20",x"3d",x"20"),
  1067 => (x"00",x"0a",x"20",x"64"),
  1068 => (x"48",x"44",x"00",x"0a"),
  1069 => (x"54",x"53",x"59",x"52"),
  1070 => (x"20",x"45",x"4e",x"4f"),
  1071 => (x"47",x"4f",x"52",x"50"),
  1072 => (x"2c",x"4d",x"41",x"52"),
  1073 => (x"4d",x"4f",x"53",x"20"),
  1074 => (x"54",x"53",x"20",x"45"),
  1075 => (x"47",x"4e",x"49",x"52"),
  1076 => (x"52",x"48",x"44",x"00"),
  1077 => (x"4f",x"54",x"53",x"59"),
  1078 => (x"50",x"20",x"45",x"4e"),
  1079 => (x"52",x"47",x"4f",x"52"),
  1080 => (x"20",x"2c",x"4d",x"41"),
  1081 => (x"54",x"53",x"27",x"31"),
  1082 => (x"52",x"54",x"53",x"20"),
  1083 => (x"00",x"47",x"4e",x"49"),
  1084 => (x"68",x"44",x"00",x"0a"),
  1085 => (x"74",x"73",x"79",x"72"),
  1086 => (x"20",x"65",x"6e",x"6f"),
  1087 => (x"63",x"6e",x"65",x"42"),
  1088 => (x"72",x"61",x"6d",x"68"),
  1089 => (x"56",x"20",x"2c",x"6b"),
  1090 => (x"69",x"73",x"72",x"65"),
  1091 => (x"32",x"20",x"6e",x"6f"),
  1092 => (x"28",x"20",x"31",x"2e"),
  1093 => (x"67",x"6e",x"61",x"4c"),
  1094 => (x"65",x"67",x"61",x"75"),
  1095 => (x"29",x"43",x"20",x"3a"),
  1096 => (x"00",x"0a",x"00",x"0a"),
  1097 => (x"63",x"65",x"78",x"45"),
  1098 => (x"6f",x"69",x"74",x"75"),
  1099 => (x"74",x"73",x"20",x"6e"),
  1100 => (x"73",x"74",x"72",x"61"),
  1101 => (x"64",x"25",x"20",x"2c"),
  1102 => (x"6e",x"75",x"72",x"20"),
  1103 => (x"68",x"74",x"20",x"73"),
  1104 => (x"67",x"75",x"6f",x"72"),
  1105 => (x"68",x"44",x"20",x"68"),
  1106 => (x"74",x"73",x"79",x"72"),
  1107 => (x"0a",x"65",x"6e",x"6f"),
  1108 => (x"65",x"78",x"45",x"00"),
  1109 => (x"69",x"74",x"75",x"63"),
  1110 => (x"65",x"20",x"6e",x"6f"),
  1111 => (x"0a",x"73",x"64",x"6e"),
  1112 => (x"46",x"00",x"0a",x"00"),
  1113 => (x"6c",x"61",x"6e",x"69"),
  1114 => (x"6c",x"61",x"76",x"20"),
  1115 => (x"20",x"73",x"65",x"75"),
  1116 => (x"74",x"20",x"66",x"6f"),
  1117 => (x"76",x"20",x"65",x"68"),
  1118 => (x"61",x"69",x"72",x"61"),
  1119 => (x"73",x"65",x"6c",x"62"),
  1120 => (x"65",x"73",x"75",x"20"),
  1121 => (x"6e",x"69",x"20",x"64"),
  1122 => (x"65",x"68",x"74",x"20"),
  1123 => (x"6e",x"65",x"62",x"20"),
  1124 => (x"61",x"6d",x"68",x"63"),
  1125 => (x"0a",x"3a",x"6b",x"72"),
  1126 => (x"49",x"00",x"0a",x"00"),
  1127 => (x"47",x"5f",x"74",x"6e"),
  1128 => (x"3a",x"62",x"6f",x"6c"),
  1129 => (x"20",x"20",x"20",x"20"),
  1130 => (x"20",x"20",x"20",x"20"),
  1131 => (x"20",x"20",x"20",x"20"),
  1132 => (x"00",x"0a",x"64",x"25"),
  1133 => (x"20",x"20",x"20",x"20"),
  1134 => (x"20",x"20",x"20",x"20"),
  1135 => (x"75",x"6f",x"68",x"73"),
  1136 => (x"62",x"20",x"64",x"6c"),
  1137 => (x"20",x"20",x"3a",x"65"),
  1138 => (x"0a",x"64",x"25",x"20"),
  1139 => (x"6f",x"6f",x"42",x"00"),
  1140 => (x"6c",x"47",x"5f",x"6c"),
  1141 => (x"20",x"3a",x"62",x"6f"),
  1142 => (x"20",x"20",x"20",x"20"),
  1143 => (x"20",x"20",x"20",x"20"),
  1144 => (x"64",x"25",x"20",x"20"),
  1145 => (x"20",x"20",x"00",x"0a"),
  1146 => (x"20",x"20",x"20",x"20"),
  1147 => (x"68",x"73",x"20",x"20"),
  1148 => (x"64",x"6c",x"75",x"6f"),
  1149 => (x"3a",x"65",x"62",x"20"),
  1150 => (x"25",x"20",x"20",x"20"),
  1151 => (x"43",x"00",x"0a",x"64"),
  1152 => (x"5f",x"31",x"5f",x"68"),
  1153 => (x"62",x"6f",x"6c",x"47"),
  1154 => (x"20",x"20",x"20",x"3a"),
  1155 => (x"20",x"20",x"20",x"20"),
  1156 => (x"20",x"20",x"20",x"20"),
  1157 => (x"00",x"0a",x"63",x"25"),
  1158 => (x"20",x"20",x"20",x"20"),
  1159 => (x"20",x"20",x"20",x"20"),
  1160 => (x"75",x"6f",x"68",x"73"),
  1161 => (x"62",x"20",x"64",x"6c"),
  1162 => (x"20",x"20",x"3a",x"65"),
  1163 => (x"0a",x"63",x"25",x"20"),
  1164 => (x"5f",x"68",x"43",x"00"),
  1165 => (x"6c",x"47",x"5f",x"32"),
  1166 => (x"20",x"3a",x"62",x"6f"),
  1167 => (x"20",x"20",x"20",x"20"),
  1168 => (x"20",x"20",x"20",x"20"),
  1169 => (x"63",x"25",x"20",x"20"),
  1170 => (x"20",x"20",x"00",x"0a"),
  1171 => (x"20",x"20",x"20",x"20"),
  1172 => (x"68",x"73",x"20",x"20"),
  1173 => (x"64",x"6c",x"75",x"6f"),
  1174 => (x"3a",x"65",x"62",x"20"),
  1175 => (x"25",x"20",x"20",x"20"),
  1176 => (x"41",x"00",x"0a",x"63"),
  1177 => (x"31",x"5f",x"72",x"72"),
  1178 => (x"6f",x"6c",x"47",x"5f"),
  1179 => (x"5d",x"38",x"5b",x"62"),
  1180 => (x"20",x"20",x"20",x"3a"),
  1181 => (x"20",x"20",x"20",x"20"),
  1182 => (x"00",x"0a",x"64",x"25"),
  1183 => (x"20",x"20",x"20",x"20"),
  1184 => (x"20",x"20",x"20",x"20"),
  1185 => (x"75",x"6f",x"68",x"73"),
  1186 => (x"62",x"20",x"64",x"6c"),
  1187 => (x"20",x"20",x"3a",x"65"),
  1188 => (x"0a",x"64",x"25",x"20"),
  1189 => (x"72",x"72",x"41",x"00"),
  1190 => (x"47",x"5f",x"32",x"5f"),
  1191 => (x"5b",x"62",x"6f",x"6c"),
  1192 => (x"37",x"5b",x"5d",x"38"),
  1193 => (x"20",x"20",x"3a",x"5d"),
  1194 => (x"64",x"25",x"20",x"20"),
  1195 => (x"20",x"20",x"00",x"0a"),
  1196 => (x"20",x"20",x"20",x"20"),
  1197 => (x"68",x"73",x"20",x"20"),
  1198 => (x"64",x"6c",x"75",x"6f"),
  1199 => (x"3a",x"65",x"62",x"20"),
  1200 => (x"4e",x"20",x"20",x"20"),
  1201 => (x"65",x"62",x"6d",x"75"),
  1202 => (x"66",x"4f",x"5f",x"72"),
  1203 => (x"6e",x"75",x"52",x"5f"),
  1204 => (x"20",x"2b",x"20",x"73"),
  1205 => (x"00",x"0a",x"30",x"31"),
  1206 => (x"5f",x"72",x"74",x"50"),
  1207 => (x"62",x"6f",x"6c",x"47"),
  1208 => (x"00",x"0a",x"3e",x"2d"),
  1209 => (x"74",x"50",x"20",x"20"),
  1210 => (x"6f",x"43",x"5f",x"72"),
  1211 => (x"20",x"3a",x"70",x"6d"),
  1212 => (x"20",x"20",x"20",x"20"),
  1213 => (x"20",x"20",x"20",x"20"),
  1214 => (x"0a",x"64",x"25",x"20"),
  1215 => (x"20",x"20",x"20",x"00"),
  1216 => (x"20",x"20",x"20",x"20"),
  1217 => (x"6f",x"68",x"73",x"20"),
  1218 => (x"20",x"64",x"6c",x"75"),
  1219 => (x"20",x"3a",x"65",x"62"),
  1220 => (x"69",x"28",x"20",x"20"),
  1221 => (x"65",x"6c",x"70",x"6d"),
  1222 => (x"74",x"6e",x"65",x"6d"),
  1223 => (x"6f",x"69",x"74",x"61"),
  1224 => (x"65",x"64",x"2d",x"6e"),
  1225 => (x"64",x"6e",x"65",x"70"),
  1226 => (x"29",x"74",x"6e",x"65"),
  1227 => (x"20",x"20",x"00",x"0a"),
  1228 => (x"63",x"73",x"69",x"44"),
  1229 => (x"20",x"20",x"3a",x"72"),
  1230 => (x"20",x"20",x"20",x"20"),
  1231 => (x"20",x"20",x"20",x"20"),
  1232 => (x"25",x"20",x"20",x"20"),
  1233 => (x"20",x"00",x"0a",x"64"),
  1234 => (x"20",x"20",x"20",x"20"),
  1235 => (x"73",x"20",x"20",x"20"),
  1236 => (x"6c",x"75",x"6f",x"68"),
  1237 => (x"65",x"62",x"20",x"64"),
  1238 => (x"20",x"20",x"20",x"3a"),
  1239 => (x"00",x"0a",x"64",x"25"),
  1240 => (x"6e",x"45",x"20",x"20"),
  1241 => (x"43",x"5f",x"6d",x"75"),
  1242 => (x"3a",x"70",x"6d",x"6f"),
  1243 => (x"20",x"20",x"20",x"20"),
  1244 => (x"20",x"20",x"20",x"20"),
  1245 => (x"0a",x"64",x"25",x"20"),
  1246 => (x"20",x"20",x"20",x"00"),
  1247 => (x"20",x"20",x"20",x"20"),
  1248 => (x"6f",x"68",x"73",x"20"),
  1249 => (x"20",x"64",x"6c",x"75"),
  1250 => (x"20",x"3a",x"65",x"62"),
  1251 => (x"64",x"25",x"20",x"20"),
  1252 => (x"20",x"20",x"00",x"0a"),
  1253 => (x"5f",x"74",x"6e",x"49"),
  1254 => (x"70",x"6d",x"6f",x"43"),
  1255 => (x"20",x"20",x"20",x"3a"),
  1256 => (x"20",x"20",x"20",x"20"),
  1257 => (x"25",x"20",x"20",x"20"),
  1258 => (x"20",x"00",x"0a",x"64"),
  1259 => (x"20",x"20",x"20",x"20"),
  1260 => (x"73",x"20",x"20",x"20"),
  1261 => (x"6c",x"75",x"6f",x"68"),
  1262 => (x"65",x"62",x"20",x"64"),
  1263 => (x"20",x"20",x"20",x"3a"),
  1264 => (x"00",x"0a",x"64",x"25"),
  1265 => (x"74",x"53",x"20",x"20"),
  1266 => (x"6f",x"43",x"5f",x"72"),
  1267 => (x"20",x"3a",x"70",x"6d"),
  1268 => (x"20",x"20",x"20",x"20"),
  1269 => (x"20",x"20",x"20",x"20"),
  1270 => (x"0a",x"73",x"25",x"20"),
  1271 => (x"20",x"20",x"20",x"00"),
  1272 => (x"20",x"20",x"20",x"20"),
  1273 => (x"6f",x"68",x"73",x"20"),
  1274 => (x"20",x"64",x"6c",x"75"),
  1275 => (x"20",x"3a",x"65",x"62"),
  1276 => (x"48",x"44",x"20",x"20"),
  1277 => (x"54",x"53",x"59",x"52"),
  1278 => (x"20",x"45",x"4e",x"4f"),
  1279 => (x"47",x"4f",x"52",x"50"),
  1280 => (x"2c",x"4d",x"41",x"52"),
  1281 => (x"4d",x"4f",x"53",x"20"),
  1282 => (x"54",x"53",x"20",x"45"),
  1283 => (x"47",x"4e",x"49",x"52"),
  1284 => (x"65",x"4e",x"00",x"0a"),
  1285 => (x"50",x"5f",x"74",x"78"),
  1286 => (x"47",x"5f",x"72",x"74"),
  1287 => (x"2d",x"62",x"6f",x"6c"),
  1288 => (x"20",x"00",x"0a",x"3e"),
  1289 => (x"72",x"74",x"50",x"20"),
  1290 => (x"6d",x"6f",x"43",x"5f"),
  1291 => (x"20",x"20",x"3a",x"70"),
  1292 => (x"20",x"20",x"20",x"20"),
  1293 => (x"20",x"20",x"20",x"20"),
  1294 => (x"00",x"0a",x"64",x"25"),
  1295 => (x"20",x"20",x"20",x"20"),
  1296 => (x"20",x"20",x"20",x"20"),
  1297 => (x"75",x"6f",x"68",x"73"),
  1298 => (x"62",x"20",x"64",x"6c"),
  1299 => (x"20",x"20",x"3a",x"65"),
  1300 => (x"6d",x"69",x"28",x"20"),
  1301 => (x"6d",x"65",x"6c",x"70"),
  1302 => (x"61",x"74",x"6e",x"65"),
  1303 => (x"6e",x"6f",x"69",x"74"),
  1304 => (x"70",x"65",x"64",x"2d"),
  1305 => (x"65",x"64",x"6e",x"65"),
  1306 => (x"2c",x"29",x"74",x"6e"),
  1307 => (x"6d",x"61",x"73",x"20"),
  1308 => (x"73",x"61",x"20",x"65"),
  1309 => (x"6f",x"62",x"61",x"20"),
  1310 => (x"00",x"0a",x"65",x"76"),
  1311 => (x"69",x"44",x"20",x"20"),
  1312 => (x"3a",x"72",x"63",x"73"),
  1313 => (x"20",x"20",x"20",x"20"),
  1314 => (x"20",x"20",x"20",x"20"),
  1315 => (x"20",x"20",x"20",x"20"),
  1316 => (x"0a",x"64",x"25",x"20"),
  1317 => (x"20",x"20",x"20",x"00"),
  1318 => (x"20",x"20",x"20",x"20"),
  1319 => (x"6f",x"68",x"73",x"20"),
  1320 => (x"20",x"64",x"6c",x"75"),
  1321 => (x"20",x"3a",x"65",x"62"),
  1322 => (x"64",x"25",x"20",x"20"),
  1323 => (x"20",x"20",x"00",x"0a"),
  1324 => (x"6d",x"75",x"6e",x"45"),
  1325 => (x"6d",x"6f",x"43",x"5f"),
  1326 => (x"20",x"20",x"3a",x"70"),
  1327 => (x"20",x"20",x"20",x"20"),
  1328 => (x"25",x"20",x"20",x"20"),
  1329 => (x"20",x"00",x"0a",x"64"),
  1330 => (x"20",x"20",x"20",x"20"),
  1331 => (x"73",x"20",x"20",x"20"),
  1332 => (x"6c",x"75",x"6f",x"68"),
  1333 => (x"65",x"62",x"20",x"64"),
  1334 => (x"20",x"20",x"20",x"3a"),
  1335 => (x"00",x"0a",x"64",x"25"),
  1336 => (x"6e",x"49",x"20",x"20"),
  1337 => (x"6f",x"43",x"5f",x"74"),
  1338 => (x"20",x"3a",x"70",x"6d"),
  1339 => (x"20",x"20",x"20",x"20"),
  1340 => (x"20",x"20",x"20",x"20"),
  1341 => (x"0a",x"64",x"25",x"20"),
  1342 => (x"20",x"20",x"20",x"00"),
  1343 => (x"20",x"20",x"20",x"20"),
  1344 => (x"6f",x"68",x"73",x"20"),
  1345 => (x"20",x"64",x"6c",x"75"),
  1346 => (x"20",x"3a",x"65",x"62"),
  1347 => (x"64",x"25",x"20",x"20"),
  1348 => (x"20",x"20",x"00",x"0a"),
  1349 => (x"5f",x"72",x"74",x"53"),
  1350 => (x"70",x"6d",x"6f",x"43"),
  1351 => (x"20",x"20",x"20",x"3a"),
  1352 => (x"20",x"20",x"20",x"20"),
  1353 => (x"25",x"20",x"20",x"20"),
  1354 => (x"20",x"00",x"0a",x"73"),
  1355 => (x"20",x"20",x"20",x"20"),
  1356 => (x"73",x"20",x"20",x"20"),
  1357 => (x"6c",x"75",x"6f",x"68"),
  1358 => (x"65",x"62",x"20",x"64"),
  1359 => (x"20",x"20",x"20",x"3a"),
  1360 => (x"59",x"52",x"48",x"44"),
  1361 => (x"4e",x"4f",x"54",x"53"),
  1362 => (x"52",x"50",x"20",x"45"),
  1363 => (x"41",x"52",x"47",x"4f"),
  1364 => (x"53",x"20",x"2c",x"4d"),
  1365 => (x"20",x"45",x"4d",x"4f"),
  1366 => (x"49",x"52",x"54",x"53"),
  1367 => (x"00",x"0a",x"47",x"4e"),
  1368 => (x"5f",x"74",x"6e",x"49"),
  1369 => (x"6f",x"4c",x"5f",x"31"),
  1370 => (x"20",x"20",x"3a",x"63"),
  1371 => (x"20",x"20",x"20",x"20"),
  1372 => (x"20",x"20",x"20",x"20"),
  1373 => (x"0a",x"64",x"25",x"20"),
  1374 => (x"20",x"20",x"20",x"00"),
  1375 => (x"20",x"20",x"20",x"20"),
  1376 => (x"6f",x"68",x"73",x"20"),
  1377 => (x"20",x"64",x"6c",x"75"),
  1378 => (x"20",x"3a",x"65",x"62"),
  1379 => (x"64",x"25",x"20",x"20"),
  1380 => (x"6e",x"49",x"00",x"0a"),
  1381 => (x"5f",x"32",x"5f",x"74"),
  1382 => (x"3a",x"63",x"6f",x"4c"),
  1383 => (x"20",x"20",x"20",x"20"),
  1384 => (x"20",x"20",x"20",x"20"),
  1385 => (x"25",x"20",x"20",x"20"),
  1386 => (x"20",x"00",x"0a",x"64"),
  1387 => (x"20",x"20",x"20",x"20"),
  1388 => (x"73",x"20",x"20",x"20"),
  1389 => (x"6c",x"75",x"6f",x"68"),
  1390 => (x"65",x"62",x"20",x"64"),
  1391 => (x"20",x"20",x"20",x"3a"),
  1392 => (x"00",x"0a",x"64",x"25"),
  1393 => (x"5f",x"74",x"6e",x"49"),
  1394 => (x"6f",x"4c",x"5f",x"33"),
  1395 => (x"20",x"20",x"3a",x"63"),
  1396 => (x"20",x"20",x"20",x"20"),
  1397 => (x"20",x"20",x"20",x"20"),
  1398 => (x"0a",x"64",x"25",x"20"),
  1399 => (x"20",x"20",x"20",x"00"),
  1400 => (x"20",x"20",x"20",x"20"),
  1401 => (x"6f",x"68",x"73",x"20"),
  1402 => (x"20",x"64",x"6c",x"75"),
  1403 => (x"20",x"3a",x"65",x"62"),
  1404 => (x"64",x"25",x"20",x"20"),
  1405 => (x"6e",x"45",x"00",x"0a"),
  1406 => (x"4c",x"5f",x"6d",x"75"),
  1407 => (x"20",x"3a",x"63",x"6f"),
  1408 => (x"20",x"20",x"20",x"20"),
  1409 => (x"20",x"20",x"20",x"20"),
  1410 => (x"25",x"20",x"20",x"20"),
  1411 => (x"20",x"00",x"0a",x"64"),
  1412 => (x"20",x"20",x"20",x"20"),
  1413 => (x"73",x"20",x"20",x"20"),
  1414 => (x"6c",x"75",x"6f",x"68"),
  1415 => (x"65",x"62",x"20",x"64"),
  1416 => (x"20",x"20",x"20",x"3a"),
  1417 => (x"00",x"0a",x"64",x"25"),
  1418 => (x"5f",x"72",x"74",x"53"),
  1419 => (x"6f",x"4c",x"5f",x"31"),
  1420 => (x"20",x"20",x"3a",x"63"),
  1421 => (x"20",x"20",x"20",x"20"),
  1422 => (x"20",x"20",x"20",x"20"),
  1423 => (x"0a",x"73",x"25",x"20"),
  1424 => (x"20",x"20",x"20",x"00"),
  1425 => (x"20",x"20",x"20",x"20"),
  1426 => (x"6f",x"68",x"73",x"20"),
  1427 => (x"20",x"64",x"6c",x"75"),
  1428 => (x"20",x"3a",x"65",x"62"),
  1429 => (x"48",x"44",x"20",x"20"),
  1430 => (x"54",x"53",x"59",x"52"),
  1431 => (x"20",x"45",x"4e",x"4f"),
  1432 => (x"47",x"4f",x"52",x"50"),
  1433 => (x"2c",x"4d",x"41",x"52"),
  1434 => (x"53",x"27",x"31",x"20"),
  1435 => (x"54",x"53",x"20",x"54"),
  1436 => (x"47",x"4e",x"49",x"52"),
  1437 => (x"74",x"53",x"00",x"0a"),
  1438 => (x"5f",x"32",x"5f",x"72"),
  1439 => (x"3a",x"63",x"6f",x"4c"),
  1440 => (x"20",x"20",x"20",x"20"),
  1441 => (x"20",x"20",x"20",x"20"),
  1442 => (x"25",x"20",x"20",x"20"),
  1443 => (x"20",x"00",x"0a",x"73"),
  1444 => (x"20",x"20",x"20",x"20"),
  1445 => (x"73",x"20",x"20",x"20"),
  1446 => (x"6c",x"75",x"6f",x"68"),
  1447 => (x"65",x"62",x"20",x"64"),
  1448 => (x"20",x"20",x"20",x"3a"),
  1449 => (x"59",x"52",x"48",x"44"),
  1450 => (x"4e",x"4f",x"54",x"53"),
  1451 => (x"52",x"50",x"20",x"45"),
  1452 => (x"41",x"52",x"47",x"4f"),
  1453 => (x"32",x"20",x"2c",x"4d"),
  1454 => (x"20",x"44",x"4e",x"27"),
  1455 => (x"49",x"52",x"54",x"53"),
  1456 => (x"00",x"0a",x"47",x"4e"),
  1457 => (x"73",x"55",x"00",x"0a"),
  1458 => (x"74",x"20",x"72",x"65"),
  1459 => (x"3a",x"65",x"6d",x"69"),
  1460 => (x"0a",x"64",x"25",x"20"),
  1461 => (x"00",x"00",x"00",x"00"),
  1462 => (x"00",x"00",x"00",x"00"),
  1463 => (x"00",x"00",x"61",x"a8"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
