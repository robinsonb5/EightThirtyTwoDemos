
package Toplevel_Config is
	constant Toplevel_UseSDRAM : boolean := false;
	constant Toplevel_UseUART : boolean := true;
	constant Toplevel_UseVGA : boolean := false;
	constant Toplevel_UseAudio : boolean := false;
end package;
