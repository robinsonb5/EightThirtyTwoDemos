
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of OSDBoot_832_ROM is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"d4",x"01"),
     1 => (x"18",x"0e",x"87",x"d7"),
     2 => (x"3e",x"27",x"0e",x"1e"),
     3 => (x"0f",x"00",x"00",x"00"),
     4 => (x"80",x"ff",x"48",x"26"),
     5 => (x"27",x"4f",x"08",x"26"),
     6 => (x"00",x"00",x"00",x"23"),
     7 => (x"00",x"30",x"27",x"4f"),
     8 => (x"c2",x"4f",x"00",x"00"),
     9 => (x"27",x"4e",x"c0",x"c0"),
    10 => (x"00",x"00",x"05",x"90"),
    11 => (x"87",x"fd",x"00",x"0f"),
    12 => (x"4e",x"c0",x"f0",x"c1"),
    13 => (x"00",x"00",x"3d",x"27"),
    14 => (x"fd",x"00",x"0f",x"00"),
    15 => (x"0e",x"4f",x"4f",x"87"),
    16 => (x"5c",x"5b",x"5a",x"5e"),
    17 => (x"8e",x"d0",x"0e",x"5d"),
    18 => (x"a6",x"c4",x"4c",x"c0"),
    19 => (x"c0",x"79",x"c0",x"49"),
    20 => (x"c0",x"4b",x"a6",x"e8"),
    21 => (x"c0",x"4a",x"66",x"e4"),
    22 => (x"c1",x"48",x"66",x"e4"),
    23 => (x"a6",x"e8",x"c0",x"80"),
    24 => (x"c1",x"48",x"12",x"58"),
    25 => (x"c0",x"c0",x"c0",x"c0"),
    26 => (x"b7",x"c0",x"c4",x"90"),
    27 => (x"a6",x"c4",x"48",x"90"),
    28 => (x"c5",x"02",x"6e",x"58"),
    29 => (x"66",x"c4",x"87",x"c3"),
    30 => (x"87",x"ff",x"c3",x"02"),
    31 => (x"c0",x"49",x"a6",x"c4"),
    32 => (x"6e",x"4a",x"6e",x"79"),
    33 => (x"a9",x"f0",x"c0",x"49"),
    34 => (x"87",x"c5",x"c3",x"02"),
    35 => (x"02",x"aa",x"e3",x"c1"),
    36 => (x"c1",x"87",x"c6",x"c3"),
    37 => (x"c0",x"02",x"aa",x"e4"),
    38 => (x"ec",x"c1",x"87",x"e3"),
    39 => (x"f0",x"c2",x"02",x"aa"),
    40 => (x"aa",x"f0",x"c1",x"87"),
    41 => (x"87",x"d5",x"c0",x"02"),
    42 => (x"02",x"aa",x"f3",x"c1"),
    43 => (x"c1",x"87",x"c9",x"c2"),
    44 => (x"c0",x"02",x"aa",x"f5"),
    45 => (x"f8",x"c1",x"87",x"c7"),
    46 => (x"f1",x"c2",x"05",x"aa"),
    47 => (x"73",x"83",x"c4",x"87"),
    48 => (x"76",x"8a",x"c4",x"4a"),
    49 => (x"6e",x"79",x"6a",x"49"),
    50 => (x"87",x"dc",x"c1",x"02"),
    51 => (x"c0",x"49",x"a6",x"c8"),
    52 => (x"49",x"a6",x"cc",x"79"),
    53 => (x"4a",x"6e",x"79",x"c0"),
    54 => (x"72",x"2a",x"b7",x"dc"),
    55 => (x"6e",x"9d",x"cf",x"4d"),
    56 => (x"c4",x"30",x"c4",x"48"),
    57 => (x"9d",x"75",x"58",x"a6"),
    58 => (x"87",x"c5",x"c0",x"02"),
    59 => (x"c1",x"49",x"a6",x"c8"),
    60 => (x"ad",x"b7",x"c9",x"79"),
    61 => (x"87",x"c6",x"c0",x"06"),
    62 => (x"c0",x"85",x"f7",x"c0"),
    63 => (x"f0",x"c0",x"87",x"c3"),
    64 => (x"02",x"66",x"c8",x"85"),
    65 => (x"75",x"87",x"cc",x"c0"),
    66 => (x"16",x"e0",x"27",x"1e"),
    67 => (x"c4",x"0f",x"00",x"00"),
    68 => (x"cc",x"84",x"c1",x"86"),
    69 => (x"80",x"c1",x"48",x"66"),
    70 => (x"cc",x"58",x"a6",x"d0"),
    71 => (x"b7",x"c8",x"49",x"66"),
    72 => (x"f1",x"fe",x"04",x"a9"),
    73 => (x"87",x"ee",x"c1",x"87"),
    74 => (x"27",x"1e",x"f0",x"c0"),
    75 => (x"00",x"00",x"16",x"e0"),
    76 => (x"c1",x"86",x"c4",x"0f"),
    77 => (x"87",x"de",x"c1",x"84"),
    78 => (x"4a",x"73",x"83",x"c4"),
    79 => (x"1e",x"6a",x"8a",x"c4"),
    80 => (x"00",x"17",x"0f",x"27"),
    81 => (x"86",x"c4",x"0f",x"00"),
    82 => (x"4c",x"74",x"4a",x"70"),
    83 => (x"c5",x"c1",x"84",x"72"),
    84 => (x"49",x"a6",x"c4",x"87"),
    85 => (x"fd",x"c0",x"79",x"c1"),
    86 => (x"73",x"83",x"c4",x"87"),
    87 => (x"6a",x"8a",x"c4",x"4a"),
    88 => (x"16",x"e0",x"27",x"1e"),
    89 => (x"c4",x"0f",x"00",x"00"),
    90 => (x"c0",x"84",x"c1",x"86"),
    91 => (x"1e",x"6e",x"87",x"e8"),
    92 => (x"00",x"16",x"e0",x"27"),
    93 => (x"86",x"c4",x"0f",x"00"),
    94 => (x"6e",x"87",x"db",x"c0"),
    95 => (x"a9",x"e5",x"c0",x"49"),
    96 => (x"87",x"c8",x"c0",x"05"),
    97 => (x"c1",x"49",x"a6",x"c4"),
    98 => (x"87",x"ca",x"c0",x"79"),
    99 => (x"e0",x"27",x"1e",x"6e"),
   100 => (x"0f",x"00",x"00",x"16"),
   101 => (x"e4",x"c0",x"86",x"c4"),
   102 => (x"e4",x"c0",x"4a",x"66"),
   103 => (x"80",x"c1",x"48",x"66"),
   104 => (x"58",x"a6",x"e8",x"c0"),
   105 => (x"c0",x"c1",x"48",x"12"),
   106 => (x"90",x"c0",x"c0",x"c0"),
   107 => (x"90",x"b7",x"c0",x"c4"),
   108 => (x"58",x"a6",x"c4",x"48"),
   109 => (x"fd",x"fa",x"05",x"6e"),
   110 => (x"d0",x"48",x"74",x"87"),
   111 => (x"26",x"4d",x"26",x"86"),
   112 => (x"26",x"4b",x"26",x"4c"),
   113 => (x"0e",x"4f",x"26",x"4a"),
   114 => (x"0e",x"5b",x"5a",x"5e"),
   115 => (x"d8",x"4a",x"66",x"cc"),
   116 => (x"9a",x"ff",x"c3",x"2a"),
   117 => (x"c8",x"4b",x"66",x"cc"),
   118 => (x"c0",x"fc",x"cf",x"2b"),
   119 => (x"73",x"4a",x"72",x"9b"),
   120 => (x"4b",x"66",x"cc",x"b2"),
   121 => (x"ff",x"c0",x"33",x"c8"),
   122 => (x"9b",x"c0",x"c0",x"f0"),
   123 => (x"b2",x"73",x"4a",x"72"),
   124 => (x"d8",x"4b",x"66",x"cc"),
   125 => (x"c0",x"fc",x"cf",x"33"),
   126 => (x"72",x"9b",x"c0",x"c0"),
   127 => (x"72",x"b2",x"73",x"4a"),
   128 => (x"26",x"4b",x"26",x"48"),
   129 => (x"0e",x"4f",x"26",x"4a"),
   130 => (x"0e",x"5b",x"5a",x"5e"),
   131 => (x"c8",x"4a",x"66",x"cc"),
   132 => (x"9a",x"ff",x"c3",x"2a"),
   133 => (x"c8",x"4b",x"66",x"cc"),
   134 => (x"c0",x"fc",x"cf",x"33"),
   135 => (x"73",x"4a",x"72",x"9b"),
   136 => (x"26",x"48",x"72",x"b2"),
   137 => (x"26",x"4a",x"26",x"4b"),
   138 => (x"5a",x"5e",x"0e",x"4f"),
   139 => (x"66",x"cc",x"0e",x"5b"),
   140 => (x"cf",x"2a",x"d0",x"4a"),
   141 => (x"4a",x"9a",x"ff",x"ff"),
   142 => (x"d0",x"4b",x"66",x"cc"),
   143 => (x"c0",x"c0",x"f0",x"33"),
   144 => (x"73",x"4a",x"72",x"9b"),
   145 => (x"26",x"48",x"72",x"b2"),
   146 => (x"26",x"4a",x"26",x"4b"),
   147 => (x"fd",x"ff",x"1e",x"4f"),
   148 => (x"1e",x"4f",x"26",x"87"),
   149 => (x"66",x"cc",x"1e",x"72"),
   150 => (x"9a",x"df",x"c3",x"4a"),
   151 => (x"c0",x"8a",x"f7",x"c0"),
   152 => (x"c0",x"03",x"aa",x"b7"),
   153 => (x"e7",x"c0",x"87",x"c3"),
   154 => (x"48",x"66",x"c8",x"82"),
   155 => (x"a6",x"cc",x"30",x"c4"),
   156 => (x"48",x"66",x"c8",x"58"),
   157 => (x"a6",x"cc",x"b0",x"72"),
   158 => (x"48",x"66",x"c8",x"58"),
   159 => (x"4f",x"26",x"4a",x"26"),
   160 => (x"5b",x"5a",x"5e",x"0e"),
   161 => (x"c0",x"0e",x"5d",x"5c"),
   162 => (x"c0",x"c0",x"e8",x"f6"),
   163 => (x"19",x"80",x"27",x"4c"),
   164 => (x"48",x"bf",x"00",x"00"),
   165 => (x"84",x"27",x"80",x"c1"),
   166 => (x"58",x"00",x"00",x"19"),
   167 => (x"4a",x"66",x"d4",x"97"),
   168 => (x"c0",x"c0",x"c0",x"c1"),
   169 => (x"c0",x"c4",x"92",x"c0"),
   170 => (x"c1",x"4a",x"92",x"b7"),
   171 => (x"05",x"aa",x"b7",x"d3"),
   172 => (x"27",x"87",x"e6",x"c0"),
   173 => (x"00",x"00",x"19",x"80"),
   174 => (x"27",x"79",x"c0",x"49"),
   175 => (x"00",x"00",x"19",x"84"),
   176 => (x"27",x"79",x"c0",x"49"),
   177 => (x"00",x"00",x"19",x"8c"),
   178 => (x"27",x"79",x"c0",x"49"),
   179 => (x"00",x"00",x"19",x"90"),
   180 => (x"c1",x"79",x"c0",x"49"),
   181 => (x"e7",x"c9",x"7c",x"d3"),
   182 => (x"19",x"80",x"27",x"87"),
   183 => (x"49",x"bf",x"00",x"00"),
   184 => (x"05",x"a9",x"b7",x"c1"),
   185 => (x"c1",x"87",x"d5",x"c1"),
   186 => (x"d4",x"97",x"7c",x"f4"),
   187 => (x"c0",x"c1",x"4a",x"66"),
   188 => (x"92",x"c0",x"c0",x"c0"),
   189 => (x"92",x"b7",x"c0",x"c4"),
   190 => (x"27",x"1e",x"72",x"4a"),
   191 => (x"00",x"00",x"19",x"90"),
   192 => (x"53",x"27",x"1e",x"bf"),
   193 => (x"0f",x"00",x"00",x"02"),
   194 => (x"94",x"27",x"86",x"c8"),
   195 => (x"58",x"00",x"00",x"19"),
   196 => (x"00",x"19",x"90",x"27"),
   197 => (x"c3",x"4d",x"bf",x"00"),
   198 => (x"c0",x"06",x"ad",x"b7"),
   199 => (x"48",x"ca",x"87",x"c6"),
   200 => (x"4d",x"70",x"88",x"75"),
   201 => (x"82",x"c1",x"4a",x"75"),
   202 => (x"30",x"c1",x"48",x"72"),
   203 => (x"00",x"19",x"8c",x"27"),
   204 => (x"48",x"75",x"58",x"00"),
   205 => (x"70",x"80",x"f0",x"c0"),
   206 => (x"87",x"c4",x"c8",x"7c"),
   207 => (x"00",x"19",x"90",x"27"),
   208 => (x"c9",x"49",x"bf",x"00"),
   209 => (x"c7",x"01",x"a9",x"b7"),
   210 => (x"90",x"27",x"87",x"f6"),
   211 => (x"bf",x"00",x"00",x"19"),
   212 => (x"a9",x"b7",x"c0",x"49"),
   213 => (x"87",x"e8",x"c7",x"06"),
   214 => (x"00",x"19",x"90",x"27"),
   215 => (x"c0",x"48",x"bf",x"00"),
   216 => (x"7c",x"70",x"80",x"f0"),
   217 => (x"00",x"19",x"80",x"27"),
   218 => (x"c3",x"49",x"bf",x"00"),
   219 => (x"c0",x"01",x"a9",x"b7"),
   220 => (x"d4",x"97",x"87",x"e9"),
   221 => (x"c0",x"c1",x"4a",x"66"),
   222 => (x"92",x"c0",x"c0",x"c0"),
   223 => (x"92",x"b7",x"c0",x"c4"),
   224 => (x"27",x"1e",x"72",x"4a"),
   225 => (x"00",x"00",x"19",x"8c"),
   226 => (x"53",x"27",x"1e",x"bf"),
   227 => (x"0f",x"00",x"00",x"02"),
   228 => (x"90",x"27",x"86",x"c8"),
   229 => (x"58",x"00",x"00",x"19"),
   230 => (x"27",x"87",x"e5",x"c6"),
   231 => (x"00",x"00",x"19",x"88"),
   232 => (x"82",x"c3",x"4a",x"bf"),
   233 => (x"00",x"19",x"80",x"27"),
   234 => (x"72",x"49",x"bf",x"00"),
   235 => (x"c0",x"01",x"a9",x"b7"),
   236 => (x"d4",x"97",x"87",x"f1"),
   237 => (x"c0",x"c1",x"4a",x"66"),
   238 => (x"92",x"c0",x"c0",x"c0"),
   239 => (x"92",x"b7",x"c0",x"c4"),
   240 => (x"27",x"1e",x"72",x"4a"),
   241 => (x"00",x"00",x"19",x"84"),
   242 => (x"53",x"27",x"1e",x"bf"),
   243 => (x"0f",x"00",x"00",x"02"),
   244 => (x"88",x"27",x"86",x"c8"),
   245 => (x"58",x"00",x"00",x"19"),
   246 => (x"00",x"19",x"94",x"27"),
   247 => (x"79",x"c1",x"49",x"00"),
   248 => (x"27",x"87",x"dd",x"c5"),
   249 => (x"00",x"00",x"19",x"90"),
   250 => (x"b7",x"c0",x"49",x"bf"),
   251 => (x"d0",x"c3",x"06",x"a9"),
   252 => (x"19",x"90",x"27",x"87"),
   253 => (x"49",x"bf",x"00",x"00"),
   254 => (x"01",x"a9",x"b7",x"c3"),
   255 => (x"27",x"87",x"c2",x"c3"),
   256 => (x"00",x"00",x"19",x"8c"),
   257 => (x"32",x"c1",x"4a",x"bf"),
   258 => (x"80",x"27",x"82",x"c1"),
   259 => (x"bf",x"00",x"00",x"19"),
   260 => (x"a9",x"b7",x"72",x"49"),
   261 => (x"87",x"c2",x"c2",x"01"),
   262 => (x"4a",x"66",x"d4",x"97"),
   263 => (x"c0",x"c0",x"c0",x"c1"),
   264 => (x"c0",x"c4",x"92",x"c0"),
   265 => (x"72",x"4a",x"92",x"b7"),
   266 => (x"19",x"98",x"27",x"1e"),
   267 => (x"1e",x"bf",x"00",x"00"),
   268 => (x"00",x"02",x"53",x"27"),
   269 => (x"86",x"c8",x"0f",x"00"),
   270 => (x"00",x"19",x"9c",x"27"),
   271 => (x"94",x"27",x"58",x"00"),
   272 => (x"bf",x"00",x"00",x"19"),
   273 => (x"27",x"8a",x"c1",x"4a"),
   274 => (x"00",x"00",x"19",x"94"),
   275 => (x"c0",x"79",x"72",x"49"),
   276 => (x"c3",x"03",x"aa",x"b7"),
   277 => (x"84",x"27",x"87",x"ea"),
   278 => (x"bf",x"00",x"00",x"19"),
   279 => (x"19",x"98",x"27",x"4a"),
   280 => (x"bf",x"97",x"00",x"00"),
   281 => (x"19",x"84",x"27",x"52"),
   282 => (x"4a",x"bf",x"00",x"00"),
   283 => (x"84",x"27",x"82",x"c1"),
   284 => (x"49",x"00",x"00",x"19"),
   285 => (x"9c",x"27",x"79",x"72"),
   286 => (x"bf",x"00",x"00",x"19"),
   287 => (x"c0",x"06",x"aa",x"b7"),
   288 => (x"9c",x"27",x"87",x"cd"),
   289 => (x"49",x"00",x"00",x"19"),
   290 => (x"00",x"19",x"84",x"27"),
   291 => (x"27",x"79",x"bf",x"00"),
   292 => (x"00",x"00",x"19",x"94"),
   293 => (x"c2",x"79",x"c1",x"49"),
   294 => (x"94",x"27",x"87",x"e6"),
   295 => (x"bf",x"00",x"00",x"19"),
   296 => (x"87",x"dc",x"c2",x"05"),
   297 => (x"00",x"19",x"98",x"27"),
   298 => (x"c4",x"4b",x"bf",x"00"),
   299 => (x"19",x"98",x"27",x"33"),
   300 => (x"73",x"49",x"00",x"00"),
   301 => (x"19",x"84",x"27",x"79"),
   302 => (x"4a",x"bf",x"00",x"00"),
   303 => (x"ff",x"c1",x"52",x"73"),
   304 => (x"19",x"90",x"27",x"87"),
   305 => (x"49",x"bf",x"00",x"00"),
   306 => (x"04",x"a9",x"b7",x"c7"),
   307 => (x"c0",x"87",x"e5",x"c1"),
   308 => (x"49",x"f4",x"fe",x"4b"),
   309 => (x"84",x"27",x"79",x"c1"),
   310 => (x"49",x"00",x"00",x"19"),
   311 => (x"9c",x"27",x"79",x"c0"),
   312 => (x"bf",x"00",x"00",x"19"),
   313 => (x"a9",x"b7",x"c0",x"49"),
   314 => (x"87",x"e5",x"c0",x"06"),
   315 => (x"00",x"19",x"84",x"27"),
   316 => (x"83",x"bf",x"bf",x"00"),
   317 => (x"00",x"19",x"84",x"27"),
   318 => (x"c4",x"4a",x"bf",x"00"),
   319 => (x"19",x"84",x"27",x"82"),
   320 => (x"72",x"49",x"00",x"00"),
   321 => (x"19",x"9c",x"27",x"79"),
   322 => (x"b7",x"bf",x"00",x"00"),
   323 => (x"db",x"ff",x"04",x"aa"),
   324 => (x"27",x"1e",x"73",x"87"),
   325 => (x"00",x"00",x"19",x"9c"),
   326 => (x"ce",x"27",x"1e",x"bf"),
   327 => (x"1e",x"00",x"00",x"17"),
   328 => (x"00",x"00",x"3f",x"27"),
   329 => (x"86",x"cc",x"0f",x"00"),
   330 => (x"27",x"7c",x"c2",x"c1"),
   331 => (x"00",x"00",x"02",x"4d"),
   332 => (x"87",x"cc",x"c0",x"0f"),
   333 => (x"00",x"19",x"90",x"27"),
   334 => (x"c0",x"48",x"bf",x"00"),
   335 => (x"7c",x"70",x"80",x"f0"),
   336 => (x"4c",x"26",x"4d",x"26"),
   337 => (x"4a",x"26",x"4b",x"26"),
   338 => (x"5e",x"0e",x"4f",x"26"),
   339 => (x"5d",x"5c",x"5b",x"5a"),
   340 => (x"4d",x"66",x"d8",x"0e"),
   341 => (x"66",x"d4",x"4c",x"c0"),
   342 => (x"2a",x"b7",x"dc",x"4a"),
   343 => (x"9b",x"cf",x"4b",x"72"),
   344 => (x"c4",x"48",x"66",x"d4"),
   345 => (x"58",x"a6",x"d8",x"30"),
   346 => (x"06",x"ab",x"b7",x"c9"),
   347 => (x"c0",x"87",x"c6",x"c0"),
   348 => (x"c3",x"c0",x"83",x"f7"),
   349 => (x"83",x"f0",x"c0",x"87"),
   350 => (x"c1",x"7d",x"97",x"73"),
   351 => (x"c8",x"84",x"c1",x"85"),
   352 => (x"ff",x"04",x"ac",x"b7"),
   353 => (x"4d",x"26",x"87",x"d0"),
   354 => (x"4b",x"26",x"4c",x"26"),
   355 => (x"4f",x"26",x"4a",x"26"),
   356 => (x"5b",x"5a",x"5e",x"0e"),
   357 => (x"cc",x"0e",x"5d",x"5c"),
   358 => (x"07",x"1e",x"27",x"8e"),
   359 => (x"27",x"1e",x"00",x"00"),
   360 => (x"00",x"00",x"17",x"0f"),
   361 => (x"27",x"86",x"c4",x"0f"),
   362 => (x"00",x"00",x"15",x"43"),
   363 => (x"72",x"4a",x"70",x"0f"),
   364 => (x"cf",x"c4",x"02",x"9a"),
   365 => (x"07",x"07",x"27",x"87"),
   366 => (x"27",x"1e",x"00",x"00"),
   367 => (x"00",x"00",x"17",x"0f"),
   368 => (x"27",x"86",x"c4",x"0f"),
   369 => (x"00",x"00",x"07",x"91"),
   370 => (x"72",x"4a",x"70",x"0f"),
   371 => (x"e5",x"c3",x"02",x"9a"),
   372 => (x"20",x"00",x"27",x"87"),
   373 => (x"27",x"1e",x"00",x"00"),
   374 => (x"00",x"00",x"06",x"df"),
   375 => (x"0e",x"50",x"27",x"1e"),
   376 => (x"c8",x"0f",x"00",x"00"),
   377 => (x"73",x"4b",x"70",x"86"),
   378 => (x"d7",x"c3",x"02",x"9b"),
   379 => (x"49",x"a6",x"c4",x"87"),
   380 => (x"00",x"20",x"00",x"27"),
   381 => (x"4d",x"c0",x"79",x"00"),
   382 => (x"9b",x"fc",x"83",x"c3"),
   383 => (x"00",x"20",x"00",x"27"),
   384 => (x"84",x"73",x"4c",x"00"),
   385 => (x"d3",x"27",x"1e",x"74"),
   386 => (x"1e",x"00",x"00",x"06"),
   387 => (x"00",x"0e",x"50",x"27"),
   388 => (x"86",x"c8",x"0f",x"00"),
   389 => (x"9a",x"72",x"4a",x"70"),
   390 => (x"87",x"e8",x"c2",x"02"),
   391 => (x"ab",x"b7",x"ff",x"c7"),
   392 => (x"87",x"e0",x"c2",x"06"),
   393 => (x"c8",x"1e",x"c0",x"c8"),
   394 => (x"82",x"75",x"4a",x"66"),
   395 => (x"43",x"27",x"1e",x"72"),
   396 => (x"0f",x"00",x"00",x"17"),
   397 => (x"4a",x"70",x"86",x"c8"),
   398 => (x"72",x"49",x"a6",x"c8"),
   399 => (x"24",x"49",x"76",x"79"),
   400 => (x"85",x"c0",x"c8",x"79"),
   401 => (x"c8",x"8b",x"c0",x"c8"),
   402 => (x"b7",x"6e",x"49",x"66"),
   403 => (x"da",x"c1",x"02",x"a9"),
   404 => (x"19",x"60",x"27",x"87"),
   405 => (x"75",x"1e",x"00",x"00"),
   406 => (x"05",x"4a",x"27",x"1e"),
   407 => (x"c8",x"0f",x"00",x"00"),
   408 => (x"19",x"68",x"27",x"86"),
   409 => (x"c0",x"49",x"00",x"00"),
   410 => (x"69",x"27",x"51",x"e0"),
   411 => (x"1e",x"00",x"00",x"19"),
   412 => (x"27",x"1e",x"66",x"cc"),
   413 => (x"00",x"00",x"05",x"4a"),
   414 => (x"27",x"86",x"c8",x"0f"),
   415 => (x"00",x"00",x"19",x"71"),
   416 => (x"51",x"e0",x"c0",x"49"),
   417 => (x"00",x"19",x"72",x"27"),
   418 => (x"66",x"c4",x"1e",x"00"),
   419 => (x"05",x"4a",x"27",x"1e"),
   420 => (x"c8",x"0f",x"00",x"00"),
   421 => (x"19",x"7a",x"27",x"86"),
   422 => (x"c0",x"49",x"00",x"00"),
   423 => (x"19",x"60",x"27",x"51"),
   424 => (x"27",x"1e",x"00",x"00"),
   425 => (x"00",x"00",x"0f",x"b6"),
   426 => (x"c7",x"86",x"c4",x"0f"),
   427 => (x"01",x"ab",x"b7",x"ff"),
   428 => (x"c0",x"87",x"f1",x"fd"),
   429 => (x"eb",x"27",x"87",x"ce"),
   430 => (x"1e",x"00",x"00",x"06"),
   431 => (x"00",x"17",x"0f",x"27"),
   432 => (x"86",x"c4",x"0f",x"00"),
   433 => (x"cc",x"87",x"fd",x"ff"),
   434 => (x"26",x"4d",x"26",x"86"),
   435 => (x"26",x"4b",x"26",x"4c"),
   436 => (x"43",x"4f",x"26",x"4a"),
   437 => (x"4b",x"43",x"45",x"48"),
   438 => (x"42",x"4d",x"55",x"53"),
   439 => (x"4f",x"00",x"4e",x"49"),
   440 => (x"33",x"38",x"44",x"53"),
   441 => (x"53",x"31",x"30",x"32"),
   442 => (x"55",x"00",x"53",x"59"),
   443 => (x"6c",x"62",x"61",x"6e"),
   444 => (x"6f",x"74",x"20",x"65"),
   445 => (x"63",x"6f",x"6c",x"20"),
   446 => (x"20",x"65",x"74",x"61"),
   447 => (x"74",x"72",x"61",x"70"),
   448 => (x"6f",x"69",x"74",x"69"),
   449 => (x"48",x"00",x"0a",x"6e"),
   450 => (x"69",x"74",x"6e",x"75"),
   451 => (x"66",x"20",x"67",x"6e"),
   452 => (x"70",x"20",x"72",x"6f"),
   453 => (x"69",x"74",x"72",x"61"),
   454 => (x"6e",x"6f",x"69",x"74"),
   455 => (x"6e",x"49",x"00",x"0a"),
   456 => (x"61",x"69",x"74",x"69"),
   457 => (x"69",x"7a",x"69",x"6c"),
   458 => (x"53",x"20",x"67",x"6e"),
   459 => (x"61",x"63",x"20",x"44"),
   460 => (x"00",x"0a",x"64",x"72"),
   461 => (x"5b",x"5a",x"5e",x"0e"),
   462 => (x"d4",x"0e",x"5d",x"5c"),
   463 => (x"4c",x"c0",x"4d",x"66"),
   464 => (x"c0",x"49",x"66",x"dc"),
   465 => (x"c0",x"06",x"a9",x"b7"),
   466 => (x"4b",x"15",x"87",x"fb"),
   467 => (x"c0",x"c0",x"c0",x"c1"),
   468 => (x"c0",x"c4",x"93",x"c0"),
   469 => (x"d8",x"4b",x"93",x"b7"),
   470 => (x"4a",x"bf",x"97",x"66"),
   471 => (x"c0",x"c0",x"c0",x"c1"),
   472 => (x"c0",x"c4",x"92",x"c0"),
   473 => (x"d8",x"4a",x"92",x"b7"),
   474 => (x"80",x"c1",x"48",x"66"),
   475 => (x"72",x"58",x"a6",x"dc"),
   476 => (x"c0",x"02",x"ab",x"b7"),
   477 => (x"48",x"c1",x"87",x"c5"),
   478 => (x"c1",x"87",x"cc",x"c0"),
   479 => (x"b7",x"66",x"dc",x"84"),
   480 => (x"c5",x"ff",x"04",x"ac"),
   481 => (x"26",x"48",x"c0",x"87"),
   482 => (x"26",x"4c",x"26",x"4d"),
   483 => (x"26",x"4a",x"26",x"4b"),
   484 => (x"5a",x"5e",x"0e",x"4f"),
   485 => (x"0e",x"5d",x"5c",x"5b"),
   486 => (x"00",x"1b",x"a8",x"27"),
   487 => (x"79",x"c0",x"49",x"00"),
   488 => (x"00",x"18",x"b6",x"27"),
   489 => (x"0f",x"27",x"1e",x"00"),
   490 => (x"0f",x"00",x"00",x"17"),
   491 => (x"a0",x"27",x"86",x"c4"),
   492 => (x"1e",x"00",x"00",x"19"),
   493 => (x"e4",x"27",x"1e",x"c0"),
   494 => (x"0f",x"00",x"00",x"15"),
   495 => (x"4a",x"70",x"86",x"c8"),
   496 => (x"c0",x"05",x"9a",x"72"),
   497 => (x"e2",x"27",x"87",x"d3"),
   498 => (x"1e",x"00",x"00",x"17"),
   499 => (x"00",x"17",x"0f",x"27"),
   500 => (x"86",x"c4",x"0f",x"00"),
   501 => (x"d8",x"cf",x"48",x"c0"),
   502 => (x"18",x"c3",x"27",x"87"),
   503 => (x"27",x"1e",x"00",x"00"),
   504 => (x"00",x"00",x"17",x"0f"),
   505 => (x"c0",x"86",x"c4",x"0f"),
   506 => (x"1b",x"d4",x"27",x"4c"),
   507 => (x"c1",x"49",x"00",x"00"),
   508 => (x"27",x"1e",x"c8",x"79"),
   509 => (x"00",x"00",x"18",x"da"),
   510 => (x"19",x"d6",x"27",x"1e"),
   511 => (x"27",x"1e",x"00",x"00"),
   512 => (x"00",x"00",x"07",x"34"),
   513 => (x"70",x"86",x"cc",x"0f"),
   514 => (x"05",x"9a",x"72",x"4a"),
   515 => (x"27",x"87",x"c8",x"c0"),
   516 => (x"00",x"00",x"1b",x"d4"),
   517 => (x"c8",x"79",x"c0",x"49"),
   518 => (x"18",x"e3",x"27",x"1e"),
   519 => (x"27",x"1e",x"00",x"00"),
   520 => (x"00",x"00",x"19",x"f2"),
   521 => (x"07",x"34",x"27",x"1e"),
   522 => (x"cc",x"0f",x"00",x"00"),
   523 => (x"72",x"4a",x"70",x"86"),
   524 => (x"c8",x"c0",x"05",x"9a"),
   525 => (x"1b",x"d4",x"27",x"87"),
   526 => (x"c0",x"49",x"00",x"00"),
   527 => (x"1b",x"d4",x"27",x"79"),
   528 => (x"1e",x"bf",x"00",x"00"),
   529 => (x"00",x"18",x"ec",x"27"),
   530 => (x"3f",x"27",x"1e",x"00"),
   531 => (x"0f",x"00",x"00",x"00"),
   532 => (x"d4",x"27",x"86",x"c8"),
   533 => (x"bf",x"00",x"00",x"1b"),
   534 => (x"87",x"c0",x"c3",x"02"),
   535 => (x"00",x"19",x"a0",x"27"),
   536 => (x"5e",x"27",x"4d",x"00"),
   537 => (x"4b",x"00",x"00",x"1b"),
   538 => (x"00",x"1b",x"9e",x"27"),
   539 => (x"4a",x"bf",x"9f",x"00"),
   540 => (x"9e",x"27",x"1e",x"72"),
   541 => (x"4a",x"00",x"00",x"1b"),
   542 => (x"00",x"19",x"a0",x"27"),
   543 => (x"1e",x"72",x"8a",x"00"),
   544 => (x"c0",x"c8",x"1e",x"d0"),
   545 => (x"18",x"14",x"27",x"1e"),
   546 => (x"27",x"1e",x"00",x"00"),
   547 => (x"00",x"00",x"00",x"3f"),
   548 => (x"73",x"86",x"d4",x"0f"),
   549 => (x"6a",x"82",x"c8",x"4a"),
   550 => (x"1b",x"9e",x"27",x"4c"),
   551 => (x"bf",x"9f",x"00",x"00"),
   552 => (x"ea",x"d6",x"c5",x"4a"),
   553 => (x"c0",x"05",x"aa",x"b7"),
   554 => (x"4a",x"73",x"87",x"d3"),
   555 => (x"1e",x"6a",x"82",x"c8"),
   556 => (x"00",x"01",x"c7",x"27"),
   557 => (x"86",x"c4",x"0f",x"00"),
   558 => (x"e4",x"c0",x"4c",x"70"),
   559 => (x"c7",x"4a",x"75",x"87"),
   560 => (x"6a",x"9f",x"82",x"fe"),
   561 => (x"d5",x"e9",x"ca",x"4a"),
   562 => (x"c0",x"02",x"aa",x"b7"),
   563 => (x"f6",x"27",x"87",x"d3"),
   564 => (x"1e",x"00",x"00",x"17"),
   565 => (x"00",x"17",x"0f",x"27"),
   566 => (x"86",x"c4",x"0f",x"00"),
   567 => (x"d0",x"cb",x"48",x"c0"),
   568 => (x"27",x"1e",x"74",x"87"),
   569 => (x"00",x"00",x"18",x"51"),
   570 => (x"00",x"3f",x"27",x"1e"),
   571 => (x"c8",x"0f",x"00",x"00"),
   572 => (x"19",x"a0",x"27",x"86"),
   573 => (x"74",x"1e",x"00",x"00"),
   574 => (x"15",x"e4",x"27",x"1e"),
   575 => (x"c8",x"0f",x"00",x"00"),
   576 => (x"72",x"4a",x"70",x"86"),
   577 => (x"c5",x"c0",x"05",x"9a"),
   578 => (x"ca",x"48",x"c0",x"87"),
   579 => (x"69",x"27",x"87",x"e3"),
   580 => (x"1e",x"00",x"00",x"18"),
   581 => (x"00",x"17",x"0f",x"27"),
   582 => (x"86",x"c4",x"0f",x"00"),
   583 => (x"00",x"18",x"ff",x"27"),
   584 => (x"3f",x"27",x"1e",x"00"),
   585 => (x"0f",x"00",x"00",x"00"),
   586 => (x"1e",x"c8",x"86",x"c4"),
   587 => (x"00",x"19",x"17",x"27"),
   588 => (x"f2",x"27",x"1e",x"00"),
   589 => (x"1e",x"00",x"00",x"19"),
   590 => (x"00",x"07",x"34",x"27"),
   591 => (x"86",x"cc",x"0f",x"00"),
   592 => (x"9a",x"72",x"4a",x"70"),
   593 => (x"87",x"cb",x"c0",x"05"),
   594 => (x"00",x"1b",x"a8",x"27"),
   595 => (x"79",x"c1",x"49",x"00"),
   596 => (x"c8",x"87",x"f1",x"c0"),
   597 => (x"19",x"20",x"27",x"1e"),
   598 => (x"27",x"1e",x"00",x"00"),
   599 => (x"00",x"00",x"19",x"d6"),
   600 => (x"07",x"34",x"27",x"1e"),
   601 => (x"cc",x"0f",x"00",x"00"),
   602 => (x"72",x"4a",x"70",x"86"),
   603 => (x"d3",x"c0",x"02",x"9a"),
   604 => (x"18",x"90",x"27",x"87"),
   605 => (x"27",x"1e",x"00",x"00"),
   606 => (x"00",x"00",x"00",x"3f"),
   607 => (x"c0",x"86",x"c4",x"0f"),
   608 => (x"87",x"ed",x"c8",x"48"),
   609 => (x"00",x"1b",x"9e",x"27"),
   610 => (x"4a",x"bf",x"97",x"00"),
   611 => (x"aa",x"b7",x"d5",x"c1"),
   612 => (x"87",x"d0",x"c0",x"05"),
   613 => (x"00",x"1b",x"9f",x"27"),
   614 => (x"4a",x"bf",x"97",x"00"),
   615 => (x"aa",x"b7",x"ea",x"c2"),
   616 => (x"87",x"c5",x"c0",x"02"),
   617 => (x"c8",x"c8",x"48",x"c0"),
   618 => (x"19",x"a0",x"27",x"87"),
   619 => (x"bf",x"97",x"00",x"00"),
   620 => (x"b7",x"e9",x"c3",x"4a"),
   621 => (x"d5",x"c0",x"02",x"aa"),
   622 => (x"19",x"a0",x"27",x"87"),
   623 => (x"bf",x"97",x"00",x"00"),
   624 => (x"b7",x"eb",x"c3",x"4a"),
   625 => (x"c5",x"c0",x"02",x"aa"),
   626 => (x"c7",x"48",x"c0",x"87"),
   627 => (x"ab",x"27",x"87",x"e3"),
   628 => (x"97",x"00",x"00",x"19"),
   629 => (x"9a",x"72",x"4a",x"bf"),
   630 => (x"87",x"cf",x"c0",x"05"),
   631 => (x"00",x"19",x"ac",x"27"),
   632 => (x"4a",x"bf",x"97",x"00"),
   633 => (x"02",x"aa",x"b7",x"c2"),
   634 => (x"c0",x"87",x"c5",x"c0"),
   635 => (x"87",x"c1",x"c7",x"48"),
   636 => (x"00",x"19",x"ad",x"27"),
   637 => (x"48",x"bf",x"97",x"00"),
   638 => (x"00",x"1b",x"a4",x"27"),
   639 => (x"a0",x"27",x"58",x"00"),
   640 => (x"bf",x"00",x"00",x"1b"),
   641 => (x"c1",x"4b",x"72",x"4a"),
   642 => (x"1b",x"a4",x"27",x"8b"),
   643 => (x"73",x"49",x"00",x"00"),
   644 => (x"72",x"1e",x"73",x"79"),
   645 => (x"19",x"29",x"27",x"1e"),
   646 => (x"27",x"1e",x"00",x"00"),
   647 => (x"00",x"00",x"00",x"3f"),
   648 => (x"27",x"86",x"cc",x"0f"),
   649 => (x"00",x"00",x"19",x"ae"),
   650 => (x"74",x"4a",x"bf",x"97"),
   651 => (x"19",x"af",x"27",x"82"),
   652 => (x"bf",x"97",x"00",x"00"),
   653 => (x"73",x"33",x"c8",x"4b"),
   654 => (x"27",x"80",x"72",x"48"),
   655 => (x"00",x"00",x"1b",x"b8"),
   656 => (x"19",x"b0",x"27",x"58"),
   657 => (x"bf",x"97",x"00",x"00"),
   658 => (x"1b",x"cc",x"27",x"48"),
   659 => (x"27",x"58",x"00",x"00"),
   660 => (x"00",x"00",x"1b",x"a8"),
   661 => (x"df",x"c3",x"02",x"bf"),
   662 => (x"27",x"1e",x"c8",x"87"),
   663 => (x"00",x"00",x"18",x"ad"),
   664 => (x"19",x"f2",x"27",x"1e"),
   665 => (x"27",x"1e",x"00",x"00"),
   666 => (x"00",x"00",x"07",x"34"),
   667 => (x"70",x"86",x"cc",x"0f"),
   668 => (x"02",x"9a",x"72",x"4a"),
   669 => (x"c0",x"87",x"c5",x"c0"),
   670 => (x"87",x"f5",x"c4",x"48"),
   671 => (x"00",x"1b",x"a0",x"27"),
   672 => (x"73",x"4b",x"bf",x"00"),
   673 => (x"27",x"30",x"c4",x"48"),
   674 => (x"00",x"00",x"1b",x"d0"),
   675 => (x"1b",x"c4",x"27",x"58"),
   676 => (x"73",x"49",x"00",x"00"),
   677 => (x"19",x"c5",x"27",x"79"),
   678 => (x"bf",x"97",x"00",x"00"),
   679 => (x"27",x"32",x"c8",x"4a"),
   680 => (x"00",x"00",x"19",x"c4"),
   681 => (x"72",x"4c",x"bf",x"97"),
   682 => (x"27",x"82",x"74",x"4a"),
   683 => (x"00",x"00",x"19",x"c6"),
   684 => (x"d0",x"4c",x"bf",x"97"),
   685 => (x"74",x"4a",x"72",x"34"),
   686 => (x"19",x"c7",x"27",x"82"),
   687 => (x"bf",x"97",x"00",x"00"),
   688 => (x"72",x"34",x"d8",x"4c"),
   689 => (x"27",x"82",x"74",x"4a"),
   690 => (x"00",x"00",x"1b",x"d0"),
   691 => (x"72",x"79",x"72",x"49"),
   692 => (x"1b",x"c8",x"27",x"4a"),
   693 => (x"92",x"bf",x"00",x"00"),
   694 => (x"b4",x"27",x"4a",x"72"),
   695 => (x"bf",x"00",x"00",x"1b"),
   696 => (x"1b",x"b8",x"27",x"82"),
   697 => (x"72",x"49",x"00",x"00"),
   698 => (x"19",x"cd",x"27",x"79"),
   699 => (x"bf",x"97",x"00",x"00"),
   700 => (x"27",x"34",x"c8",x"4c"),
   701 => (x"00",x"00",x"19",x"cc"),
   702 => (x"74",x"4d",x"bf",x"97"),
   703 => (x"27",x"84",x"75",x"4c"),
   704 => (x"00",x"00",x"19",x"ce"),
   705 => (x"d0",x"4d",x"bf",x"97"),
   706 => (x"75",x"4c",x"74",x"35"),
   707 => (x"19",x"cf",x"27",x"84"),
   708 => (x"bf",x"97",x"00",x"00"),
   709 => (x"d8",x"9d",x"cf",x"4d"),
   710 => (x"75",x"4c",x"74",x"35"),
   711 => (x"1b",x"bc",x"27",x"84"),
   712 => (x"74",x"49",x"00",x"00"),
   713 => (x"73",x"8c",x"c2",x"79"),
   714 => (x"73",x"93",x"74",x"4b"),
   715 => (x"27",x"80",x"72",x"48"),
   716 => (x"00",x"00",x"1b",x"c4"),
   717 => (x"87",x"f7",x"c1",x"58"),
   718 => (x"00",x"19",x"b2",x"27"),
   719 => (x"4a",x"bf",x"97",x"00"),
   720 => (x"b1",x"27",x"32",x"c8"),
   721 => (x"97",x"00",x"00",x"19"),
   722 => (x"4a",x"72",x"4b",x"bf"),
   723 => (x"cc",x"27",x"82",x"73"),
   724 => (x"49",x"00",x"00",x"1b"),
   725 => (x"32",x"c5",x"79",x"72"),
   726 => (x"c9",x"82",x"ff",x"c7"),
   727 => (x"1b",x"c4",x"27",x"2a"),
   728 => (x"72",x"49",x"00",x"00"),
   729 => (x"19",x"b7",x"27",x"79"),
   730 => (x"bf",x"97",x"00",x"00"),
   731 => (x"27",x"33",x"c8",x"4b"),
   732 => (x"00",x"00",x"19",x"b6"),
   733 => (x"73",x"4c",x"bf",x"97"),
   734 => (x"27",x"83",x"74",x"4b"),
   735 => (x"00",x"00",x"1b",x"d0"),
   736 => (x"73",x"79",x"73",x"49"),
   737 => (x"1b",x"c8",x"27",x"4b"),
   738 => (x"93",x"bf",x"00",x"00"),
   739 => (x"b4",x"27",x"4b",x"73"),
   740 => (x"bf",x"00",x"00",x"1b"),
   741 => (x"1b",x"c0",x"27",x"83"),
   742 => (x"73",x"49",x"00",x"00"),
   743 => (x"1b",x"bc",x"27",x"79"),
   744 => (x"c0",x"49",x"00",x"00"),
   745 => (x"72",x"48",x"73",x"79"),
   746 => (x"1b",x"bc",x"27",x"80"),
   747 => (x"c1",x"58",x"00",x"00"),
   748 => (x"26",x"4d",x"26",x"48"),
   749 => (x"26",x"4b",x"26",x"4c"),
   750 => (x"0e",x"4f",x"26",x"4a"),
   751 => (x"5c",x"5b",x"5a",x"5e"),
   752 => (x"a8",x"27",x"0e",x"5d"),
   753 => (x"bf",x"00",x"00",x"1b"),
   754 => (x"87",x"cf",x"c0",x"02"),
   755 => (x"c7",x"4c",x"66",x"d4"),
   756 => (x"66",x"d4",x"2c",x"b7"),
   757 => (x"9b",x"ff",x"c1",x"4b"),
   758 => (x"d4",x"87",x"cc",x"c0"),
   759 => (x"b7",x"c8",x"4c",x"66"),
   760 => (x"4b",x"66",x"d4",x"2c"),
   761 => (x"27",x"9b",x"ff",x"c3"),
   762 => (x"00",x"00",x"19",x"a0"),
   763 => (x"1b",x"b4",x"27",x"1e"),
   764 => (x"4a",x"bf",x"00",x"00"),
   765 => (x"1e",x"72",x"82",x"74"),
   766 => (x"00",x"15",x"e4",x"27"),
   767 => (x"86",x"c8",x"0f",x"00"),
   768 => (x"9a",x"72",x"4a",x"70"),
   769 => (x"87",x"c5",x"c0",x"05"),
   770 => (x"f2",x"c0",x"48",x"c0"),
   771 => (x"1b",x"a8",x"27",x"87"),
   772 => (x"02",x"bf",x"00",x"00"),
   773 => (x"73",x"87",x"d7",x"c0"),
   774 => (x"72",x"92",x"c4",x"4a"),
   775 => (x"19",x"a0",x"27",x"4a"),
   776 => (x"6a",x"82",x"00",x"00"),
   777 => (x"ff",x"ff",x"cf",x"4d"),
   778 => (x"c0",x"9d",x"ff",x"ff"),
   779 => (x"4a",x"73",x"87",x"cf"),
   780 => (x"4a",x"72",x"92",x"c2"),
   781 => (x"00",x"19",x"a0",x"27"),
   782 => (x"6a",x"9f",x"82",x"00"),
   783 => (x"26",x"48",x"75",x"4d"),
   784 => (x"26",x"4c",x"26",x"4d"),
   785 => (x"26",x"4a",x"26",x"4b"),
   786 => (x"5a",x"5e",x"0e",x"4f"),
   787 => (x"0e",x"5d",x"5c",x"5b"),
   788 => (x"ff",x"cf",x"8e",x"cc"),
   789 => (x"4d",x"f8",x"ff",x"ff"),
   790 => (x"49",x"76",x"4c",x"c0"),
   791 => (x"00",x"1b",x"bc",x"27"),
   792 => (x"c4",x"79",x"bf",x"00"),
   793 => (x"c0",x"27",x"49",x"a6"),
   794 => (x"bf",x"00",x"00",x"1b"),
   795 => (x"1b",x"a8",x"27",x"79"),
   796 => (x"02",x"bf",x"00",x"00"),
   797 => (x"27",x"87",x"cc",x"c0"),
   798 => (x"00",x"00",x"1b",x"a0"),
   799 => (x"32",x"c4",x"4a",x"bf"),
   800 => (x"27",x"87",x"c9",x"c0"),
   801 => (x"00",x"00",x"1b",x"c4"),
   802 => (x"32",x"c4",x"4a",x"bf"),
   803 => (x"72",x"49",x"a6",x"c8"),
   804 => (x"c8",x"4b",x"c0",x"79"),
   805 => (x"a9",x"c0",x"49",x"66"),
   806 => (x"87",x"d0",x"c3",x"06"),
   807 => (x"9a",x"cf",x"4a",x"73"),
   808 => (x"c0",x"05",x"9a",x"72"),
   809 => (x"a0",x"27",x"87",x"e4"),
   810 => (x"1e",x"00",x"00",x"19"),
   811 => (x"c8",x"4a",x"66",x"c8"),
   812 => (x"80",x"c1",x"48",x"66"),
   813 => (x"72",x"58",x"a6",x"cc"),
   814 => (x"15",x"e4",x"27",x"1e"),
   815 => (x"c8",x"0f",x"00",x"00"),
   816 => (x"19",x"a0",x"27",x"86"),
   817 => (x"c0",x"4c",x"00",x"00"),
   818 => (x"e0",x"c0",x"87",x"c3"),
   819 => (x"4a",x"6c",x"97",x"84"),
   820 => (x"c2",x"02",x"9a",x"72"),
   821 => (x"6c",x"97",x"87",x"cd"),
   822 => (x"b7",x"e5",x"c3",x"4a"),
   823 => (x"c2",x"c2",x"02",x"aa"),
   824 => (x"cb",x"4a",x"74",x"87"),
   825 => (x"4a",x"6a",x"97",x"82"),
   826 => (x"9a",x"72",x"9a",x"d8"),
   827 => (x"87",x"f3",x"c1",x"05"),
   828 => (x"0f",x"27",x"1e",x"74"),
   829 => (x"0f",x"00",x"00",x"17"),
   830 => (x"1e",x"cb",x"86",x"c4"),
   831 => (x"1e",x"66",x"e8",x"c0"),
   832 => (x"34",x"27",x"1e",x"74"),
   833 => (x"0f",x"00",x"00",x"07"),
   834 => (x"4a",x"70",x"86",x"cc"),
   835 => (x"c1",x"05",x"9a",x"72"),
   836 => (x"4b",x"74",x"87",x"d1"),
   837 => (x"e0",x"c0",x"83",x"dc"),
   838 => (x"82",x"c4",x"4a",x"66"),
   839 => (x"4b",x"74",x"7a",x"6b"),
   840 => (x"e0",x"c0",x"83",x"da"),
   841 => (x"82",x"c8",x"4a",x"66"),
   842 => (x"70",x"48",x"6b",x"9f"),
   843 => (x"27",x"4d",x"72",x"7a"),
   844 => (x"00",x"00",x"1b",x"a8"),
   845 => (x"d5",x"c0",x"02",x"bf"),
   846 => (x"d4",x"4a",x"74",x"87"),
   847 => (x"4a",x"6a",x"9f",x"82"),
   848 => (x"9a",x"ff",x"ff",x"c0"),
   849 => (x"30",x"d0",x"48",x"72"),
   850 => (x"c0",x"58",x"a6",x"c4"),
   851 => (x"49",x"76",x"87",x"c4"),
   852 => (x"48",x"6e",x"79",x"c0"),
   853 => (x"7d",x"70",x"80",x"6d"),
   854 => (x"49",x"66",x"e0",x"c0"),
   855 => (x"48",x"c1",x"79",x"c0"),
   856 => (x"c1",x"87",x"ce",x"c1"),
   857 => (x"ab",x"66",x"c8",x"83"),
   858 => (x"87",x"f0",x"fc",x"04"),
   859 => (x"ff",x"ff",x"ff",x"cf"),
   860 => (x"a8",x"27",x"4d",x"f8"),
   861 => (x"bf",x"00",x"00",x"1b"),
   862 => (x"87",x"f3",x"c0",x"02"),
   863 => (x"bb",x"27",x"1e",x"6e"),
   864 => (x"0f",x"00",x"00",x"0b"),
   865 => (x"a6",x"c4",x"86",x"c4"),
   866 => (x"75",x"4a",x"6e",x"58"),
   867 => (x"02",x"aa",x"75",x"9a"),
   868 => (x"6e",x"87",x"dc",x"c0"),
   869 => (x"72",x"8a",x"c2",x"4a"),
   870 => (x"1b",x"a0",x"27",x"4a"),
   871 => (x"92",x"bf",x"00",x"00"),
   872 => (x"00",x"1b",x"b8",x"27"),
   873 => (x"72",x"48",x"bf",x"00"),
   874 => (x"58",x"a6",x"c8",x"80"),
   875 => (x"c0",x"87",x"e2",x"fb"),
   876 => (x"ff",x"ff",x"cf",x"48"),
   877 => (x"cc",x"4d",x"f8",x"ff"),
   878 => (x"26",x"4d",x"26",x"86"),
   879 => (x"26",x"4b",x"26",x"4c"),
   880 => (x"0e",x"4f",x"26",x"4a"),
   881 => (x"0e",x"5b",x"5a",x"5e"),
   882 => (x"4a",x"bf",x"66",x"cc"),
   883 => (x"66",x"cc",x"82",x"c1"),
   884 => (x"72",x"79",x"72",x"49"),
   885 => (x"1b",x"a4",x"27",x"4a"),
   886 => (x"9a",x"bf",x"00",x"00"),
   887 => (x"c0",x"05",x"9a",x"72"),
   888 => (x"66",x"cc",x"87",x"d3"),
   889 => (x"6a",x"82",x"c8",x"4a"),
   890 => (x"0b",x"bb",x"27",x"1e"),
   891 => (x"c4",x"0f",x"00",x"00"),
   892 => (x"73",x"4b",x"70",x"86"),
   893 => (x"26",x"48",x"c1",x"7a"),
   894 => (x"26",x"4a",x"26",x"4b"),
   895 => (x"5a",x"5e",x"0e",x"4f"),
   896 => (x"b8",x"27",x"0e",x"5b"),
   897 => (x"bf",x"00",x"00",x"1b"),
   898 => (x"4b",x"66",x"cc",x"4a"),
   899 => (x"4b",x"6b",x"83",x"c8"),
   900 => (x"4b",x"73",x"8b",x"c2"),
   901 => (x"00",x"1b",x"a0",x"27"),
   902 => (x"72",x"93",x"bf",x"00"),
   903 => (x"27",x"82",x"73",x"4a"),
   904 => (x"00",x"00",x"1b",x"a4"),
   905 => (x"66",x"cc",x"4b",x"bf"),
   906 => (x"4a",x"72",x"9b",x"bf"),
   907 => (x"66",x"d0",x"82",x"73"),
   908 => (x"27",x"1e",x"72",x"1e"),
   909 => (x"00",x"00",x"15",x"e4"),
   910 => (x"70",x"86",x"c8",x"0f"),
   911 => (x"05",x"9a",x"72",x"4a"),
   912 => (x"c0",x"87",x"c5",x"c0"),
   913 => (x"87",x"c2",x"c0",x"48"),
   914 => (x"4b",x"26",x"48",x"c1"),
   915 => (x"4f",x"26",x"4a",x"26"),
   916 => (x"5b",x"5a",x"5e",x"0e"),
   917 => (x"d8",x"0e",x"5d",x"5c"),
   918 => (x"66",x"d4",x"4c",x"66"),
   919 => (x"1b",x"d8",x"27",x"1e"),
   920 => (x"27",x"1e",x"00",x"00"),
   921 => (x"00",x"00",x"0c",x"49"),
   922 => (x"70",x"86",x"c8",x"0f"),
   923 => (x"02",x"9a",x"72",x"4a"),
   924 => (x"27",x"87",x"df",x"c1"),
   925 => (x"00",x"00",x"1b",x"dc"),
   926 => (x"ff",x"c7",x"4a",x"bf"),
   927 => (x"72",x"2a",x"c9",x"82"),
   928 => (x"27",x"4b",x"c0",x"4d"),
   929 => (x"00",x"00",x"0e",x"f4"),
   930 => (x"17",x"0f",x"27",x"1e"),
   931 => (x"c4",x"0f",x"00",x"00"),
   932 => (x"ad",x"b7",x"c0",x"86"),
   933 => (x"87",x"d0",x"c1",x"06"),
   934 => (x"d8",x"27",x"1e",x"74"),
   935 => (x"1e",x"00",x"00",x"1b"),
   936 => (x"00",x"0d",x"fd",x"27"),
   937 => (x"86",x"c8",x"0f",x"00"),
   938 => (x"9a",x"72",x"4a",x"70"),
   939 => (x"87",x"c5",x"c0",x"05"),
   940 => (x"f5",x"c0",x"48",x"c0"),
   941 => (x"1b",x"d8",x"27",x"87"),
   942 => (x"27",x"1e",x"00",x"00"),
   943 => (x"00",x"00",x"0d",x"c3"),
   944 => (x"c8",x"86",x"c4",x"0f"),
   945 => (x"83",x"c1",x"84",x"c0"),
   946 => (x"04",x"ab",x"b7",x"75"),
   947 => (x"c0",x"87",x"c9",x"ff"),
   948 => (x"66",x"d4",x"87",x"d6"),
   949 => (x"0f",x"0d",x"27",x"1e"),
   950 => (x"27",x"1e",x"00",x"00"),
   951 => (x"00",x"00",x"00",x"3f"),
   952 => (x"c0",x"86",x"c8",x"0f"),
   953 => (x"87",x"c2",x"c0",x"48"),
   954 => (x"4d",x"26",x"48",x"c1"),
   955 => (x"4b",x"26",x"4c",x"26"),
   956 => (x"4f",x"26",x"4a",x"26"),
   957 => (x"6e",x"65",x"70",x"4f"),
   958 => (x"66",x"20",x"64",x"65"),
   959 => (x"2c",x"65",x"6c",x"69"),
   960 => (x"61",x"6f",x"6c",x"20"),
   961 => (x"67",x"6e",x"69",x"64"),
   962 => (x"0a",x"2e",x"2e",x"2e"),
   963 => (x"6e",x"61",x"43",x"00"),
   964 => (x"6f",x"20",x"74",x"27"),
   965 => (x"20",x"6e",x"65",x"70"),
   966 => (x"00",x"0a",x"73",x"25"),
   967 => (x"c8",x"1e",x"72",x"1e"),
   968 => (x"d1",x"c0",x"02",x"66"),
   969 => (x"1b",x"e4",x"27",x"87"),
   970 => (x"c8",x"49",x"00",x"00"),
   971 => (x"ec",x"27",x"79",x"66"),
   972 => (x"49",x"00",x"00",x"1b"),
   973 => (x"ec",x"27",x"79",x"c0"),
   974 => (x"05",x"00",x"00",x"1b"),
   975 => (x"27",x"87",x"db",x"c0"),
   976 => (x"00",x"00",x"1b",x"e4"),
   977 => (x"c4",x"48",x"72",x"4a"),
   978 => (x"1b",x"e8",x"27",x"80"),
   979 => (x"27",x"58",x"00",x"00"),
   980 => (x"00",x"00",x"1b",x"e8"),
   981 => (x"c0",x"79",x"6a",x"49"),
   982 => (x"e8",x"27",x"87",x"ce"),
   983 => (x"48",x"00",x"00",x"1b"),
   984 => (x"ec",x"27",x"30",x"c8"),
   985 => (x"58",x"00",x"00",x"1b"),
   986 => (x"00",x"1b",x"ec",x"27"),
   987 => (x"82",x"c1",x"4a",x"00"),
   988 => (x"98",x"c3",x"48",x"72"),
   989 => (x"00",x"1b",x"f0",x"27"),
   990 => (x"e8",x"27",x"58",x"00"),
   991 => (x"4a",x"00",x"00",x"1b"),
   992 => (x"72",x"2a",x"b7",x"d8"),
   993 => (x"26",x"4a",x"26",x"48"),
   994 => (x"5a",x"5e",x"0e",x"4f"),
   995 => (x"66",x"cc",x"0e",x"5b"),
   996 => (x"87",x"c8",x"fe",x"1e"),
   997 => (x"4b",x"70",x"86",x"c4"),
   998 => (x"9b",x"73",x"4a",x"c0"),
   999 => (x"87",x"ce",x"c0",x"02"),
  1000 => (x"1e",x"c0",x"82",x"c1"),
  1001 => (x"c4",x"87",x"f5",x"fd"),
  1002 => (x"ff",x"4b",x"70",x"86"),
  1003 => (x"48",x"72",x"87",x"ec"),
  1004 => (x"4a",x"26",x"4b",x"26"),
  1005 => (x"5e",x"0e",x"4f",x"26"),
  1006 => (x"5d",x"5c",x"5b",x"5a"),
  1007 => (x"c0",x"8e",x"c8",x"0e"),
  1008 => (x"c4",x"c0",x"e4",x"f6"),
  1009 => (x"e4",x"f6",x"c0",x"4c"),
  1010 => (x"dc",x"4b",x"c0",x"c0"),
  1011 => (x"f8",x"fe",x"1e",x"66"),
  1012 => (x"70",x"86",x"c4",x"87"),
  1013 => (x"c2",x"4d",x"72",x"4a"),
  1014 => (x"c1",x"49",x"76",x"85"),
  1015 => (x"7c",x"9f",x"d0",x"79"),
  1016 => (x"9f",x"c1",x"c0",x"c1"),
  1017 => (x"4a",x"6b",x"9f",x"7b"),
  1018 => (x"c0",x"7b",x"9f",x"c0"),
  1019 => (x"6b",x"9f",x"7b",x"9f"),
  1020 => (x"58",x"a6",x"c8",x"48"),
  1021 => (x"72",x"9a",x"c0",x"c4"),
  1022 => (x"fd",x"c1",x"02",x"9a"),
  1023 => (x"c0",x"02",x"6e",x"87"),
  1024 => (x"66",x"c4",x"87",x"e6"),
  1025 => (x"c6",x"c0",x"c8",x"49"),
  1026 => (x"ed",x"c1",x"05",x"a9"),
  1027 => (x"c0",x"49",x"76",x"87"),
  1028 => (x"ca",x"eb",x"fa",x"79"),
  1029 => (x"9f",x"c1",x"7b",x"9f"),
  1030 => (x"7b",x"9f",x"c0",x"7b"),
  1031 => (x"c0",x"7b",x"9f",x"75"),
  1032 => (x"9f",x"c0",x"7b",x"9f"),
  1033 => (x"87",x"d2",x"c1",x"7b"),
  1034 => (x"2a",x"c1",x"4a",x"75"),
  1035 => (x"b2",x"c0",x"c0",x"c8"),
  1036 => (x"72",x"49",x"66",x"c4"),
  1037 => (x"c1",x"c1",x"05",x"a9"),
  1038 => (x"1e",x"66",x"dc",x"87"),
  1039 => (x"c4",x"87",x"dd",x"fb"),
  1040 => (x"58",x"a6",x"c4",x"86"),
  1041 => (x"8d",x"c1",x"4a",x"75"),
  1042 => (x"c0",x"02",x"9a",x"72"),
  1043 => (x"4c",x"6e",x"87",x"de"),
  1044 => (x"74",x"7b",x"97",x"74"),
  1045 => (x"c9",x"c0",x"02",x"9c"),
  1046 => (x"fa",x"1e",x"c0",x"87"),
  1047 => (x"86",x"c4",x"87",x"fe"),
  1048 => (x"4a",x"75",x"4c",x"70"),
  1049 => (x"9a",x"72",x"8d",x"c1"),
  1050 => (x"87",x"e4",x"ff",x"05"),
  1051 => (x"c0",x"e4",x"f6",x"c0"),
  1052 => (x"9f",x"d1",x"4c",x"c4"),
  1053 => (x"c0",x"48",x"c1",x"7c"),
  1054 => (x"9f",x"d1",x"87",x"c6"),
  1055 => (x"87",x"dd",x"fd",x"7c"),
  1056 => (x"4d",x"26",x"86",x"c8"),
  1057 => (x"4b",x"26",x"4c",x"26"),
  1058 => (x"4f",x"26",x"4a",x"26"),
  1059 => (x"5b",x"5a",x"5e",x"0e"),
  1060 => (x"e4",x"c0",x"0e",x"5c"),
  1061 => (x"4c",x"ff",x"c3",x"8e"),
  1062 => (x"c0",x"e4",x"f6",x"c0"),
  1063 => (x"7b",x"74",x"4b",x"c0"),
  1064 => (x"9a",x"74",x"4a",x"6b"),
  1065 => (x"48",x"6b",x"7b",x"74"),
  1066 => (x"a6",x"c4",x"98",x"74"),
  1067 => (x"c8",x"48",x"6e",x"58"),
  1068 => (x"58",x"a6",x"c8",x"30"),
  1069 => (x"72",x"49",x"a6",x"c8"),
  1070 => (x"c4",x"4a",x"72",x"79"),
  1071 => (x"7b",x"74",x"b2",x"66"),
  1072 => (x"98",x"74",x"48",x"6b"),
  1073 => (x"cc",x"58",x"a6",x"d0"),
  1074 => (x"30",x"d0",x"48",x"66"),
  1075 => (x"d4",x"58",x"a6",x"d4"),
  1076 => (x"79",x"72",x"49",x"a6"),
  1077 => (x"66",x"d0",x"4a",x"72"),
  1078 => (x"6b",x"7b",x"74",x"b2"),
  1079 => (x"dc",x"98",x"74",x"48"),
  1080 => (x"66",x"d8",x"58",x"a6"),
  1081 => (x"c0",x"30",x"d8",x"48"),
  1082 => (x"c0",x"58",x"a6",x"e0"),
  1083 => (x"72",x"49",x"a6",x"e0"),
  1084 => (x"dc",x"4a",x"72",x"79"),
  1085 => (x"48",x"72",x"b2",x"66"),
  1086 => (x"26",x"86",x"e4",x"c0"),
  1087 => (x"26",x"4b",x"26",x"4c"),
  1088 => (x"0e",x"4f",x"26",x"4a"),
  1089 => (x"5c",x"5b",x"5a",x"5e"),
  1090 => (x"c3",x"8e",x"d8",x"0e"),
  1091 => (x"f6",x"c0",x"4c",x"ff"),
  1092 => (x"4b",x"c0",x"c0",x"e4"),
  1093 => (x"4a",x"6b",x"7b",x"74"),
  1094 => (x"7b",x"74",x"9a",x"74"),
  1095 => (x"48",x"6b",x"32",x"c8"),
  1096 => (x"a6",x"c4",x"98",x"74"),
  1097 => (x"49",x"a6",x"c4",x"58"),
  1098 => (x"4a",x"72",x"79",x"72"),
  1099 => (x"7b",x"74",x"b2",x"6e"),
  1100 => (x"48",x"6b",x"32",x"c8"),
  1101 => (x"a6",x"cc",x"98",x"74"),
  1102 => (x"49",x"a6",x"cc",x"58"),
  1103 => (x"4a",x"72",x"79",x"72"),
  1104 => (x"74",x"b2",x"66",x"c8"),
  1105 => (x"6b",x"32",x"c8",x"7b"),
  1106 => (x"d4",x"98",x"74",x"48"),
  1107 => (x"a6",x"d4",x"58",x"a6"),
  1108 => (x"72",x"79",x"72",x"49"),
  1109 => (x"b2",x"66",x"d0",x"4a"),
  1110 => (x"86",x"d8",x"48",x"72"),
  1111 => (x"4b",x"26",x"4c",x"26"),
  1112 => (x"4f",x"26",x"4a",x"26"),
  1113 => (x"5b",x"5a",x"5e",x"0e"),
  1114 => (x"c0",x"0e",x"5d",x"5c"),
  1115 => (x"c0",x"c0",x"e4",x"f6"),
  1116 => (x"48",x"66",x"d4",x"4b"),
  1117 => (x"70",x"98",x"ff",x"c3"),
  1118 => (x"1b",x"f0",x"27",x"7b"),
  1119 => (x"05",x"bf",x"00",x"00"),
  1120 => (x"d8",x"87",x"c8",x"c0"),
  1121 => (x"30",x"c9",x"48",x"66"),
  1122 => (x"d8",x"58",x"a6",x"dc"),
  1123 => (x"2a",x"d8",x"4a",x"66"),
  1124 => (x"ff",x"c3",x"48",x"72"),
  1125 => (x"d8",x"7b",x"70",x"98"),
  1126 => (x"2a",x"d0",x"4a",x"66"),
  1127 => (x"ff",x"c3",x"48",x"72"),
  1128 => (x"d8",x"7b",x"70",x"98"),
  1129 => (x"2a",x"c8",x"4a",x"66"),
  1130 => (x"ff",x"c3",x"48",x"72"),
  1131 => (x"d8",x"7b",x"70",x"98"),
  1132 => (x"ff",x"c3",x"48",x"66"),
  1133 => (x"d4",x"7b",x"70",x"98"),
  1134 => (x"2a",x"d0",x"4a",x"66"),
  1135 => (x"ff",x"c3",x"48",x"72"),
  1136 => (x"6b",x"7b",x"70",x"98"),
  1137 => (x"9d",x"ff",x"c3",x"4d"),
  1138 => (x"4c",x"ff",x"f0",x"c9"),
  1139 => (x"ad",x"b7",x"ff",x"c3"),
  1140 => (x"87",x"d8",x"c0",x"05"),
  1141 => (x"72",x"4a",x"ff",x"c3"),
  1142 => (x"72",x"4d",x"6b",x"7b"),
  1143 => (x"74",x"8c",x"c1",x"9d"),
  1144 => (x"c7",x"c0",x"02",x"9c"),
  1145 => (x"ad",x"b7",x"72",x"87"),
  1146 => (x"87",x"eb",x"ff",x"02"),
  1147 => (x"4d",x"27",x"1e",x"75"),
  1148 => (x"1e",x"00",x"00",x"19"),
  1149 => (x"00",x"00",x"3f",x"27"),
  1150 => (x"86",x"c8",x"0f",x"00"),
  1151 => (x"4d",x"26",x"48",x"75"),
  1152 => (x"4b",x"26",x"4c",x"26"),
  1153 => (x"4f",x"26",x"4a",x"26"),
  1154 => (x"5b",x"5a",x"5e",x"0e"),
  1155 => (x"e4",x"f6",x"c0",x"0e"),
  1156 => (x"c0",x"4b",x"c0",x"c0"),
  1157 => (x"7b",x"ff",x"c3",x"4a"),
  1158 => (x"c8",x"c3",x"82",x"c1"),
  1159 => (x"ff",x"04",x"aa",x"b7"),
  1160 => (x"4b",x"26",x"87",x"f3"),
  1161 => (x"4f",x"26",x"4a",x"26"),
  1162 => (x"5b",x"5a",x"5e",x"0e"),
  1163 => (x"c1",x"0e",x"5d",x"5c"),
  1164 => (x"c0",x"c0",x"c0",x"c0"),
  1165 => (x"f6",x"c0",x"4c",x"c0"),
  1166 => (x"4b",x"c0",x"c0",x"e4"),
  1167 => (x"00",x"12",x"08",x"27"),
  1168 => (x"f8",x"c4",x"0f",x"00"),
  1169 => (x"1e",x"c0",x"4d",x"df"),
  1170 => (x"c1",x"f0",x"ff",x"c0"),
  1171 => (x"64",x"27",x"1e",x"f7"),
  1172 => (x"0f",x"00",x"00",x"11"),
  1173 => (x"4a",x"70",x"86",x"c8"),
  1174 => (x"05",x"aa",x"b7",x"c1"),
  1175 => (x"72",x"87",x"dc",x"c1"),
  1176 => (x"12",x"e9",x"27",x"1e"),
  1177 => (x"27",x"1e",x"00",x"00"),
  1178 => (x"00",x"00",x"00",x"3f"),
  1179 => (x"c3",x"86",x"c8",x"0f"),
  1180 => (x"1e",x"74",x"7b",x"ff"),
  1181 => (x"c1",x"f0",x"e1",x"c0"),
  1182 => (x"64",x"27",x"1e",x"e9"),
  1183 => (x"0f",x"00",x"00",x"11"),
  1184 => (x"4a",x"70",x"86",x"c8"),
  1185 => (x"c0",x"05",x"9a",x"72"),
  1186 => (x"1e",x"72",x"87",x"d8"),
  1187 => (x"00",x"12",x"df",x"27"),
  1188 => (x"3f",x"27",x"1e",x"00"),
  1189 => (x"0f",x"00",x"00",x"00"),
  1190 => (x"ff",x"c3",x"86",x"c8"),
  1191 => (x"c0",x"48",x"c1",x"7b"),
  1192 => (x"1e",x"72",x"87",x"f3"),
  1193 => (x"00",x"12",x"f3",x"27"),
  1194 => (x"3f",x"27",x"1e",x"00"),
  1195 => (x"0f",x"00",x"00",x"00"),
  1196 => (x"08",x"27",x"86",x"c8"),
  1197 => (x"0f",x"00",x"00",x"12"),
  1198 => (x"72",x"87",x"d0",x"c0"),
  1199 => (x"12",x"fd",x"27",x"1e"),
  1200 => (x"27",x"1e",x"00",x"00"),
  1201 => (x"00",x"00",x"00",x"3f"),
  1202 => (x"c1",x"86",x"c8",x"0f"),
  1203 => (x"05",x"9d",x"75",x"8d"),
  1204 => (x"c0",x"87",x"f3",x"fd"),
  1205 => (x"26",x"4d",x"26",x"48"),
  1206 => (x"26",x"4b",x"26",x"4c"),
  1207 => (x"43",x"4f",x"26",x"4a"),
  1208 => (x"31",x"34",x"44",x"4d"),
  1209 => (x"0a",x"64",x"25",x"20"),
  1210 => (x"44",x"4d",x"43",x"00"),
  1211 => (x"25",x"20",x"35",x"35"),
  1212 => (x"43",x"00",x"0a",x"64"),
  1213 => (x"31",x"34",x"44",x"4d"),
  1214 => (x"0a",x"64",x"25",x"20"),
  1215 => (x"44",x"4d",x"43",x"00"),
  1216 => (x"25",x"20",x"35",x"35"),
  1217 => (x"0e",x"00",x"0a",x"64"),
  1218 => (x"5c",x"5b",x"5a",x"5e"),
  1219 => (x"ff",x"c0",x"0e",x"5d"),
  1220 => (x"4d",x"c1",x"c1",x"f0"),
  1221 => (x"c0",x"e4",x"f6",x"c0"),
  1222 => (x"ff",x"c3",x"4b",x"c0"),
  1223 => (x"13",x"99",x"27",x"7b"),
  1224 => (x"27",x"1e",x"00",x"00"),
  1225 => (x"00",x"00",x"17",x"0f"),
  1226 => (x"d3",x"86",x"c4",x"0f"),
  1227 => (x"75",x"1e",x"c0",x"4c"),
  1228 => (x"11",x"64",x"27",x"1e"),
  1229 => (x"c8",x"0f",x"00",x"00"),
  1230 => (x"72",x"4a",x"70",x"86"),
  1231 => (x"d8",x"c0",x"05",x"9a"),
  1232 => (x"27",x"1e",x"72",x"87"),
  1233 => (x"00",x"00",x"13",x"83"),
  1234 => (x"00",x"3f",x"27",x"1e"),
  1235 => (x"c8",x"0f",x"00",x"00"),
  1236 => (x"7b",x"ff",x"c3",x"86"),
  1237 => (x"e0",x"c0",x"48",x"c1"),
  1238 => (x"27",x"1e",x"72",x"87"),
  1239 => (x"00",x"00",x"13",x"8e"),
  1240 => (x"00",x"3f",x"27",x"1e"),
  1241 => (x"c8",x"0f",x"00",x"00"),
  1242 => (x"12",x"08",x"27",x"86"),
  1243 => (x"c1",x"0f",x"00",x"00"),
  1244 => (x"05",x"9c",x"74",x"8c"),
  1245 => (x"c0",x"87",x"f6",x"fe"),
  1246 => (x"26",x"4d",x"26",x"48"),
  1247 => (x"26",x"4b",x"26",x"4c"),
  1248 => (x"69",x"4f",x"26",x"4a"),
  1249 => (x"20",x"74",x"69",x"6e"),
  1250 => (x"20",x"0a",x"64",x"25"),
  1251 => (x"6e",x"69",x"00",x"20"),
  1252 => (x"25",x"20",x"74",x"69"),
  1253 => (x"20",x"20",x"0a",x"64"),
  1254 => (x"64",x"6d",x"43",x"00"),
  1255 => (x"69",x"6e",x"69",x"5f"),
  1256 => (x"0e",x"00",x"0a",x"74"),
  1257 => (x"5c",x"5b",x"5a",x"5e"),
  1258 => (x"c3",x"1e",x"0e",x"5d"),
  1259 => (x"f6",x"c0",x"4d",x"ff"),
  1260 => (x"4b",x"c0",x"c0",x"e4"),
  1261 => (x"00",x"12",x"08",x"27"),
  1262 => (x"ea",x"c6",x"0f",x"00"),
  1263 => (x"f0",x"e1",x"c0",x"1e"),
  1264 => (x"27",x"1e",x"c8",x"c1"),
  1265 => (x"00",x"00",x"11",x"64"),
  1266 => (x"70",x"86",x"c8",x"0f"),
  1267 => (x"27",x"1e",x"72",x"4a"),
  1268 => (x"00",x"00",x"15",x"2c"),
  1269 => (x"00",x"3f",x"27",x"1e"),
  1270 => (x"c8",x"0f",x"00",x"00"),
  1271 => (x"aa",x"b7",x"c1",x"86"),
  1272 => (x"87",x"cb",x"c0",x"02"),
  1273 => (x"00",x"13",x"07",x"27"),
  1274 => (x"48",x"c0",x"0f",x"00"),
  1275 => (x"27",x"87",x"db",x"c3"),
  1276 => (x"00",x"00",x"11",x"03"),
  1277 => (x"74",x"4c",x"70",x"0f"),
  1278 => (x"ff",x"ff",x"cf",x"4a"),
  1279 => (x"b7",x"ea",x"c6",x"9a"),
  1280 => (x"db",x"c0",x"02",x"aa"),
  1281 => (x"27",x"1e",x"74",x"87"),
  1282 => (x"00",x"00",x"14",x"d5"),
  1283 => (x"00",x"3f",x"27",x"1e"),
  1284 => (x"c8",x"0f",x"00",x"00"),
  1285 => (x"13",x"07",x"27",x"86"),
  1286 => (x"c0",x"0f",x"00",x"00"),
  1287 => (x"87",x"ea",x"c2",x"48"),
  1288 => (x"49",x"76",x"7b",x"75"),
  1289 => (x"27",x"79",x"f1",x"c0"),
  1290 => (x"00",x"00",x"12",x"28"),
  1291 => (x"72",x"4a",x"70",x"0f"),
  1292 => (x"eb",x"c1",x"02",x"9a"),
  1293 => (x"c0",x"1e",x"c0",x"87"),
  1294 => (x"fa",x"c1",x"f0",x"ff"),
  1295 => (x"11",x"64",x"27",x"1e"),
  1296 => (x"c8",x"0f",x"00",x"00"),
  1297 => (x"74",x"4c",x"70",x"86"),
  1298 => (x"c3",x"c1",x"05",x"9c"),
  1299 => (x"27",x"1e",x"74",x"87"),
  1300 => (x"00",x"00",x"14",x"ea"),
  1301 => (x"00",x"3f",x"27",x"1e"),
  1302 => (x"c8",x"0f",x"00",x"00"),
  1303 => (x"6b",x"7b",x"75",x"86"),
  1304 => (x"74",x"9c",x"75",x"4c"),
  1305 => (x"14",x"f6",x"27",x"1e"),
  1306 => (x"27",x"1e",x"00",x"00"),
  1307 => (x"00",x"00",x"00",x"3f"),
  1308 => (x"75",x"86",x"c8",x"0f"),
  1309 => (x"75",x"7b",x"75",x"7b"),
  1310 => (x"74",x"7b",x"75",x"7b"),
  1311 => (x"9a",x"c0",x"c1",x"4a"),
  1312 => (x"c0",x"02",x"9a",x"72"),
  1313 => (x"48",x"c1",x"87",x"c5"),
  1314 => (x"c0",x"87",x"ff",x"c0"),
  1315 => (x"87",x"fa",x"c0",x"48"),
  1316 => (x"04",x"27",x"1e",x"74"),
  1317 => (x"1e",x"00",x"00",x"15"),
  1318 => (x"00",x"00",x"3f",x"27"),
  1319 => (x"86",x"c8",x"0f",x"00"),
  1320 => (x"b7",x"c2",x"49",x"6e"),
  1321 => (x"d3",x"c0",x"05",x"a9"),
  1322 => (x"15",x"10",x"27",x"87"),
  1323 => (x"27",x"1e",x"00",x"00"),
  1324 => (x"00",x"00",x"00",x"3f"),
  1325 => (x"c0",x"86",x"c4",x"0f"),
  1326 => (x"87",x"ce",x"c0",x"48"),
  1327 => (x"88",x"c1",x"48",x"6e"),
  1328 => (x"6e",x"58",x"a6",x"c4"),
  1329 => (x"87",x"df",x"fd",x"05"),
  1330 => (x"26",x"26",x"48",x"c0"),
  1331 => (x"26",x"4c",x"26",x"4d"),
  1332 => (x"26",x"4a",x"26",x"4b"),
  1333 => (x"44",x"4d",x"43",x"4f"),
  1334 => (x"20",x"34",x"5f",x"38"),
  1335 => (x"70",x"73",x"65",x"72"),
  1336 => (x"65",x"73",x"6e",x"6f"),
  1337 => (x"64",x"25",x"20",x"3a"),
  1338 => (x"4d",x"43",x"00",x"0a"),
  1339 => (x"20",x"38",x"35",x"44"),
  1340 => (x"20",x"0a",x"64",x"25"),
  1341 => (x"4d",x"43",x"00",x"20"),
  1342 => (x"5f",x"38",x"35",x"44"),
  1343 => (x"64",x"25",x"20",x"32"),
  1344 => (x"00",x"20",x"20",x"0a"),
  1345 => (x"35",x"44",x"4d",x"43"),
  1346 => (x"64",x"25",x"20",x"38"),
  1347 => (x"00",x"20",x"20",x"0a"),
  1348 => (x"43",x"48",x"44",x"53"),
  1349 => (x"69",x"6e",x"49",x"20"),
  1350 => (x"6c",x"61",x"69",x"74"),
  1351 => (x"74",x"61",x"7a",x"69"),
  1352 => (x"20",x"6e",x"6f",x"69"),
  1353 => (x"6f",x"72",x"72",x"65"),
  1354 => (x"00",x"0a",x"21",x"72"),
  1355 => (x"5f",x"64",x"6d",x"63"),
  1356 => (x"38",x"44",x"4d",x"43"),
  1357 => (x"73",x"65",x"72",x"20"),
  1358 => (x"73",x"6e",x"6f",x"70"),
  1359 => (x"25",x"20",x"3a",x"65"),
  1360 => (x"0e",x"00",x"0a",x"64"),
  1361 => (x"5c",x"5b",x"5a",x"5e"),
  1362 => (x"f6",x"c0",x"0e",x"5d"),
  1363 => (x"4d",x"c0",x"c0",x"e4"),
  1364 => (x"c0",x"e4",x"f6",x"c0"),
  1365 => (x"f0",x"27",x"4b",x"c4"),
  1366 => (x"49",x"00",x"00",x"1b"),
  1367 => (x"f6",x"c0",x"79",x"c1"),
  1368 => (x"49",x"c8",x"c0",x"e4"),
  1369 => (x"c7",x"79",x"e0",x"c0"),
  1370 => (x"27",x"7b",x"c3",x"4c"),
  1371 => (x"00",x"00",x"12",x"08"),
  1372 => (x"c3",x"7b",x"c2",x"0f"),
  1373 => (x"1e",x"c0",x"7d",x"ff"),
  1374 => (x"c1",x"d0",x"e5",x"c0"),
  1375 => (x"64",x"27",x"1e",x"c0"),
  1376 => (x"0f",x"00",x"00",x"11"),
  1377 => (x"4a",x"70",x"86",x"c8"),
  1378 => (x"05",x"aa",x"b7",x"c1"),
  1379 => (x"c1",x"87",x"c2",x"c0"),
  1380 => (x"ac",x"b7",x"c2",x"4c"),
  1381 => (x"87",x"c5",x"c0",x"05"),
  1382 => (x"f8",x"c0",x"48",x"c0"),
  1383 => (x"74",x"8c",x"c1",x"87"),
  1384 => (x"c4",x"ff",x"05",x"9c"),
  1385 => (x"13",x"a3",x"27",x"87"),
  1386 => (x"27",x"0f",x"00",x"00"),
  1387 => (x"00",x"00",x"1b",x"f4"),
  1388 => (x"1b",x"f0",x"27",x"58"),
  1389 => (x"05",x"bf",x"00",x"00"),
  1390 => (x"c1",x"87",x"d0",x"c0"),
  1391 => (x"f0",x"ff",x"c0",x"1e"),
  1392 => (x"27",x"1e",x"d0",x"c1"),
  1393 => (x"00",x"00",x"11",x"64"),
  1394 => (x"c3",x"86",x"c8",x"0f"),
  1395 => (x"7b",x"c3",x"7d",x"ff"),
  1396 => (x"c1",x"7d",x"ff",x"c3"),
  1397 => (x"26",x"4d",x"26",x"48"),
  1398 => (x"26",x"4b",x"26",x"4c"),
  1399 => (x"1e",x"4f",x"26",x"4a"),
  1400 => (x"4f",x"26",x"48",x"c0"),
  1401 => (x"5b",x"5a",x"5e",x"0e"),
  1402 => (x"c8",x"0e",x"5d",x"5c"),
  1403 => (x"66",x"e0",x"c0",x"8e"),
  1404 => (x"e4",x"f6",x"c0",x"4d"),
  1405 => (x"76",x"4b",x"c0",x"c0"),
  1406 => (x"75",x"79",x"c0",x"49"),
  1407 => (x"66",x"e0",x"c0",x"1e"),
  1408 => (x"16",x"c9",x"27",x"1e"),
  1409 => (x"27",x"1e",x"00",x"00"),
  1410 => (x"00",x"00",x"00",x"3f"),
  1411 => (x"c3",x"86",x"cc",x"0f"),
  1412 => (x"f6",x"c0",x"7b",x"ff"),
  1413 => (x"49",x"c4",x"c0",x"e4"),
  1414 => (x"f6",x"c0",x"79",x"c2"),
  1415 => (x"49",x"c8",x"c0",x"e4"),
  1416 => (x"ff",x"c3",x"79",x"c1"),
  1417 => (x"1e",x"66",x"dc",x"7b"),
  1418 => (x"c1",x"f0",x"ff",x"c0"),
  1419 => (x"64",x"27",x"1e",x"d1"),
  1420 => (x"0f",x"00",x"00",x"11"),
  1421 => (x"a6",x"c8",x"86",x"c8"),
  1422 => (x"02",x"66",x"c4",x"58"),
  1423 => (x"c4",x"87",x"d8",x"c0"),
  1424 => (x"e0",x"c0",x"1e",x"66"),
  1425 => (x"a9",x"27",x"1e",x"66"),
  1426 => (x"1e",x"00",x"00",x"16"),
  1427 => (x"00",x"00",x"3f",x"27"),
  1428 => (x"86",x"cc",x"0f",x"00"),
  1429 => (x"c5",x"87",x"c4",x"c1"),
  1430 => (x"4c",x"df",x"cd",x"ee"),
  1431 => (x"6b",x"7b",x"ff",x"c3"),
  1432 => (x"9a",x"ff",x"c3",x"4a"),
  1433 => (x"aa",x"b7",x"fe",x"c3"),
  1434 => (x"87",x"dc",x"c0",x"05"),
  1435 => (x"8c",x"27",x"4a",x"c0"),
  1436 => (x"0f",x"00",x"00",x"10"),
  1437 => (x"85",x"c4",x"7d",x"70"),
  1438 => (x"c0",x"c2",x"82",x"c1"),
  1439 => (x"ff",x"04",x"aa",x"b7"),
  1440 => (x"4c",x"c1",x"87",x"ec"),
  1441 => (x"79",x"c1",x"49",x"76"),
  1442 => (x"9c",x"74",x"8c",x"c1"),
  1443 => (x"87",x"cc",x"ff",x"05"),
  1444 => (x"c0",x"7b",x"ff",x"c3"),
  1445 => (x"c4",x"c0",x"e4",x"f6"),
  1446 => (x"6e",x"79",x"c3",x"49"),
  1447 => (x"26",x"86",x"c8",x"48"),
  1448 => (x"26",x"4c",x"26",x"4d"),
  1449 => (x"26",x"4a",x"26",x"4b"),
  1450 => (x"61",x"65",x"52",x"4f"),
  1451 => (x"6f",x"63",x"20",x"64"),
  1452 => (x"6e",x"61",x"6d",x"6d"),
  1453 => (x"61",x"66",x"20",x"64"),
  1454 => (x"64",x"65",x"6c",x"69"),
  1455 => (x"20",x"74",x"61",x"20"),
  1456 => (x"28",x"20",x"64",x"25"),
  1457 => (x"0a",x"29",x"64",x"25"),
  1458 => (x"5f",x"64",x"73",x"00"),
  1459 => (x"64",x"61",x"65",x"72"),
  1460 => (x"63",x"65",x"73",x"5f"),
  1461 => (x"20",x"72",x"6f",x"74"),
  1462 => (x"20",x"2c",x"64",x"25"),
  1463 => (x"00",x"0a",x"64",x"25"),
  1464 => (x"1e",x"1e",x"72",x"1e"),
  1465 => (x"c0",x"e8",x"f6",x"c0"),
  1466 => (x"48",x"6a",x"4a",x"c0"),
  1467 => (x"c4",x"98",x"c0",x"c4"),
  1468 => (x"05",x"6e",x"58",x"a6"),
  1469 => (x"6a",x"87",x"cd",x"c0"),
  1470 => (x"98",x"c0",x"c4",x"48"),
  1471 => (x"6e",x"58",x"a6",x"c4"),
  1472 => (x"87",x"f3",x"ff",x"02"),
  1473 => (x"cc",x"7a",x"66",x"cc"),
  1474 => (x"26",x"26",x"48",x"66"),
  1475 => (x"0e",x"4f",x"26",x"4a"),
  1476 => (x"5c",x"5b",x"5a",x"5e"),
  1477 => (x"4b",x"66",x"d0",x"0e"),
  1478 => (x"4a",x"13",x"4c",x"c0"),
  1479 => (x"c0",x"c0",x"c0",x"c1"),
  1480 => (x"c0",x"c4",x"92",x"c0"),
  1481 => (x"72",x"4a",x"92",x"b7"),
  1482 => (x"16",x"e0",x"27",x"1e"),
  1483 => (x"c4",x"0f",x"00",x"00"),
  1484 => (x"72",x"84",x"c1",x"86"),
  1485 => (x"e1",x"ff",x"05",x"9a"),
  1486 => (x"26",x"48",x"74",x"87"),
  1487 => (x"26",x"4b",x"26",x"4c"),
  1488 => (x"0e",x"4f",x"26",x"4a"),
  1489 => (x"5c",x"5b",x"5a",x"5e"),
  1490 => (x"8e",x"c8",x"0e",x"5d"),
  1491 => (x"4c",x"66",x"e0",x"c0"),
  1492 => (x"76",x"4a",x"66",x"dc"),
  1493 => (x"c0",x"79",x"c0",x"49"),
  1494 => (x"c1",x"06",x"ac",x"b7"),
  1495 => (x"4b",x"12",x"87",x"e2"),
  1496 => (x"8c",x"c1",x"33",x"c8"),
  1497 => (x"06",x"ac",x"b7",x"c0"),
  1498 => (x"12",x"87",x"c8",x"c0"),
  1499 => (x"58",x"a6",x"c8",x"48"),
  1500 => (x"c4",x"87",x"c5",x"c0"),
  1501 => (x"79",x"c0",x"49",x"a6"),
  1502 => (x"66",x"c4",x"4b",x"73"),
  1503 => (x"c1",x"33",x"c8",x"b3"),
  1504 => (x"ac",x"b7",x"c0",x"8c"),
  1505 => (x"87",x"c5",x"c0",x"06"),
  1506 => (x"c2",x"c0",x"4d",x"12"),
  1507 => (x"73",x"4d",x"c0",x"87"),
  1508 => (x"c8",x"b3",x"75",x"4b"),
  1509 => (x"c0",x"8c",x"c1",x"33"),
  1510 => (x"c0",x"06",x"ac",x"b7"),
  1511 => (x"48",x"12",x"87",x"c8"),
  1512 => (x"c0",x"58",x"a6",x"c8"),
  1513 => (x"a6",x"c4",x"87",x"c5"),
  1514 => (x"73",x"79",x"c0",x"49"),
  1515 => (x"b3",x"66",x"c4",x"4b"),
  1516 => (x"80",x"6e",x"48",x"73"),
  1517 => (x"c1",x"58",x"a6",x"c4"),
  1518 => (x"ac",x"b7",x"c0",x"8c"),
  1519 => (x"87",x"de",x"fe",x"01"),
  1520 => (x"86",x"c8",x"48",x"6e"),
  1521 => (x"4c",x"26",x"4d",x"26"),
  1522 => (x"4a",x"26",x"4b",x"26"),
  1523 => (x"68",x"43",x"4f",x"26"),
  1524 => (x"73",x"6b",x"63",x"65"),
  1525 => (x"74",x"20",x"6d",x"75"),
  1526 => (x"64",x"25",x"20",x"6f"),
  1527 => (x"64",x"25",x"20",x"3a"),
  1528 => (x"65",x"52",x"00",x"0a"),
  1529 => (x"6f",x"20",x"64",x"61"),
  1530 => (x"42",x"4d",x"20",x"66"),
  1531 => (x"61",x"66",x"20",x"52"),
  1532 => (x"64",x"65",x"6c",x"69"),
  1533 => (x"6f",x"4e",x"00",x"0a"),
  1534 => (x"72",x"61",x"70",x"20"),
  1535 => (x"69",x"74",x"69",x"74"),
  1536 => (x"73",x"20",x"6e",x"6f"),
  1537 => (x"61",x"6e",x"67",x"69"),
  1538 => (x"65",x"72",x"75",x"74"),
  1539 => (x"75",x"6f",x"66",x"20"),
  1540 => (x"00",x"0a",x"64",x"6e"),
  1541 => (x"73",x"52",x"42",x"4d"),
  1542 => (x"3a",x"65",x"7a",x"69"),
  1543 => (x"2c",x"64",x"25",x"20"),
  1544 => (x"72",x"61",x"70",x"20"),
  1545 => (x"69",x"74",x"69",x"74"),
  1546 => (x"69",x"73",x"6e",x"6f"),
  1547 => (x"20",x"3a",x"65",x"7a"),
  1548 => (x"20",x"2c",x"64",x"25"),
  1549 => (x"73",x"66",x"66",x"6f"),
  1550 => (x"6f",x"20",x"74",x"65"),
  1551 => (x"69",x"73",x"20",x"66"),
  1552 => (x"25",x"20",x"3a",x"67"),
  1553 => (x"73",x"20",x"2c",x"64"),
  1554 => (x"30",x"20",x"67",x"69"),
  1555 => (x"0a",x"78",x"25",x"78"),
  1556 => (x"61",x"65",x"52",x"00"),
  1557 => (x"67",x"6e",x"69",x"64"),
  1558 => (x"6f",x"6f",x"62",x"20"),
  1559 => (x"65",x"73",x"20",x"74"),
  1560 => (x"72",x"6f",x"74",x"63"),
  1561 => (x"0a",x"64",x"25",x"20"),
  1562 => (x"61",x"65",x"52",x"00"),
  1563 => (x"6f",x"62",x"20",x"64"),
  1564 => (x"73",x"20",x"74",x"6f"),
  1565 => (x"6f",x"74",x"63",x"65"),
  1566 => (x"72",x"66",x"20",x"72"),
  1567 => (x"66",x"20",x"6d",x"6f"),
  1568 => (x"74",x"73",x"72",x"69"),
  1569 => (x"72",x"61",x"70",x"20"),
  1570 => (x"69",x"74",x"69",x"74"),
  1571 => (x"00",x"0a",x"6e",x"6f"),
  1572 => (x"75",x"73",x"6e",x"55"),
  1573 => (x"72",x"6f",x"70",x"70"),
  1574 => (x"20",x"64",x"65",x"74"),
  1575 => (x"74",x"72",x"61",x"70"),
  1576 => (x"6f",x"69",x"74",x"69"),
  1577 => (x"79",x"74",x"20",x"6e"),
  1578 => (x"0d",x"21",x"65",x"70"),
  1579 => (x"54",x"41",x"46",x"00"),
  1580 => (x"20",x"20",x"32",x"33"),
  1581 => (x"65",x"52",x"00",x"20"),
  1582 => (x"6e",x"69",x"64",x"61"),
  1583 => (x"42",x"4d",x"20",x"67"),
  1584 => (x"4d",x"00",x"0a",x"52"),
  1585 => (x"73",x"20",x"52",x"42"),
  1586 => (x"65",x"63",x"63",x"75"),
  1587 => (x"75",x"66",x"73",x"73"),
  1588 => (x"20",x"79",x"6c",x"6c"),
  1589 => (x"64",x"61",x"65",x"72"),
  1590 => (x"41",x"46",x"00",x"0a"),
  1591 => (x"20",x"36",x"31",x"54"),
  1592 => (x"46",x"00",x"20",x"20"),
  1593 => (x"32",x"33",x"54",x"41"),
  1594 => (x"00",x"20",x"20",x"20"),
  1595 => (x"74",x"72",x"61",x"50"),
  1596 => (x"6f",x"69",x"74",x"69"),
  1597 => (x"75",x"6f",x"63",x"6e"),
  1598 => (x"25",x"20",x"74",x"6e"),
  1599 => (x"48",x"00",x"0a",x"64"),
  1600 => (x"69",x"74",x"6e",x"75"),
  1601 => (x"66",x"20",x"67",x"6e"),
  1602 => (x"66",x"20",x"72",x"6f"),
  1603 => (x"73",x"65",x"6c",x"69"),
  1604 => (x"65",x"74",x"73",x"79"),
  1605 => (x"46",x"00",x"0a",x"6d"),
  1606 => (x"32",x"33",x"54",x"41"),
  1607 => (x"00",x"20",x"20",x"20"),
  1608 => (x"31",x"54",x"41",x"46"),
  1609 => (x"20",x"20",x"20",x"36"),
  1610 => (x"75",x"6c",x"43",x"00"),
  1611 => (x"72",x"65",x"74",x"73"),
  1612 => (x"7a",x"69",x"73",x"20"),
  1613 => (x"25",x"20",x"3a",x"65"),
  1614 => (x"43",x"20",x"2c",x"64"),
  1615 => (x"74",x"73",x"75",x"6c"),
  1616 => (x"6d",x"20",x"72",x"65"),
  1617 => (x"2c",x"6b",x"73",x"61"),
  1618 => (x"0a",x"64",x"25",x"20"),
  1619 => (x"74",x"6f",x"47",x"00"),
  1620 => (x"73",x"65",x"72",x"20"),
  1621 => (x"20",x"74",x"6c",x"75"),
  1622 => (x"0a",x"20",x"64",x"25"),
  1623 => (x"0a",x"20",x"64",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
