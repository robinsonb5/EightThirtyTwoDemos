
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of OSDBoot_832_ROM is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"d7",x"01"),
     1 => (x"58",x"0e",x"87",x"da"),
     2 => (x"27",x"0e",x"59",x"5e"),
     3 => (x"00",x"00",x"00",x"41"),
     4 => (x"26",x"49",x"26",x"0f"),
     5 => (x"26",x"80",x"ff",x"48"),
     6 => (x"26",x"27",x"4f",x"08"),
     7 => (x"4f",x"00",x"00",x"00"),
     8 => (x"00",x"00",x"33",x"27"),
     9 => (x"c0",x"c2",x"4f",x"00"),
    10 => (x"9f",x"27",x"4e",x"c0"),
    11 => (x"0f",x"00",x"00",x"05"),
    12 => (x"c1",x"87",x"fd",x"00"),
    13 => (x"27",x"4e",x"c0",x"f0"),
    14 => (x"00",x"00",x"00",x"40"),
    15 => (x"87",x"fd",x"00",x"0f"),
    16 => (x"5e",x"0e",x"4f",x"4f"),
    17 => (x"5d",x"5c",x"5b",x"5a"),
    18 => (x"c0",x"8e",x"d0",x"0e"),
    19 => (x"49",x"a6",x"c4",x"4c"),
    20 => (x"e8",x"c0",x"79",x"c0"),
    21 => (x"e4",x"c0",x"4b",x"a6"),
    22 => (x"e4",x"c0",x"4a",x"66"),
    23 => (x"80",x"c1",x"48",x"66"),
    24 => (x"58",x"a6",x"e8",x"c0"),
    25 => (x"c0",x"c1",x"48",x"12"),
    26 => (x"90",x"c0",x"c0",x"c0"),
    27 => (x"90",x"b7",x"c0",x"c4"),
    28 => (x"58",x"a6",x"c4",x"48"),
    29 => (x"c2",x"c5",x"02",x"6e"),
    30 => (x"02",x"66",x"c4",x"87"),
    31 => (x"c4",x"87",x"fe",x"c3"),
    32 => (x"79",x"c0",x"49",x"a6"),
    33 => (x"49",x"6e",x"4a",x"6e"),
    34 => (x"02",x"a9",x"f0",x"c0"),
    35 => (x"c1",x"87",x"c4",x"c3"),
    36 => (x"c3",x"02",x"aa",x"e3"),
    37 => (x"e4",x"c1",x"87",x"c5"),
    38 => (x"e3",x"c0",x"02",x"aa"),
    39 => (x"aa",x"ec",x"c1",x"87"),
    40 => (x"87",x"ef",x"c2",x"02"),
    41 => (x"02",x"aa",x"f0",x"c1"),
    42 => (x"c1",x"87",x"d5",x"c0"),
    43 => (x"c2",x"02",x"aa",x"f3"),
    44 => (x"f5",x"c1",x"87",x"c8"),
    45 => (x"c7",x"c0",x"02",x"aa"),
    46 => (x"aa",x"f8",x"c1",x"87"),
    47 => (x"87",x"f0",x"c2",x"05"),
    48 => (x"4a",x"73",x"83",x"c4"),
    49 => (x"49",x"76",x"8a",x"c4"),
    50 => (x"02",x"6e",x"79",x"6a"),
    51 => (x"c8",x"87",x"db",x"c1"),
    52 => (x"79",x"c0",x"49",x"a6"),
    53 => (x"c0",x"49",x"a6",x"cc"),
    54 => (x"dc",x"4a",x"6e",x"79"),
    55 => (x"4d",x"72",x"2a",x"b7"),
    56 => (x"48",x"6e",x"9d",x"cf"),
    57 => (x"a6",x"c4",x"30",x"c4"),
    58 => (x"02",x"9d",x"75",x"58"),
    59 => (x"c8",x"87",x"c5",x"c0"),
    60 => (x"79",x"c1",x"49",x"a6"),
    61 => (x"c0",x"06",x"ad",x"c9"),
    62 => (x"f7",x"c0",x"87",x"c6"),
    63 => (x"87",x"c3",x"c0",x"85"),
    64 => (x"c8",x"85",x"f0",x"c0"),
    65 => (x"cc",x"c0",x"02",x"66"),
    66 => (x"27",x"1e",x"75",x"87"),
    67 => (x"00",x"00",x"17",x"f6"),
    68 => (x"c1",x"86",x"c4",x"0f"),
    69 => (x"48",x"66",x"cc",x"84"),
    70 => (x"a6",x"d0",x"80",x"c1"),
    71 => (x"49",x"66",x"cc",x"58"),
    72 => (x"04",x"a9",x"b7",x"c8"),
    73 => (x"c1",x"87",x"f2",x"fe"),
    74 => (x"f0",x"c0",x"87",x"ee"),
    75 => (x"17",x"f6",x"27",x"1e"),
    76 => (x"c4",x"0f",x"00",x"00"),
    77 => (x"c1",x"84",x"c1",x"86"),
    78 => (x"83",x"c4",x"87",x"de"),
    79 => (x"8a",x"c4",x"4a",x"73"),
    80 => (x"25",x"27",x"1e",x"6a"),
    81 => (x"0f",x"00",x"00",x"18"),
    82 => (x"4a",x"70",x"86",x"c4"),
    83 => (x"84",x"72",x"4c",x"74"),
    84 => (x"c4",x"87",x"c5",x"c1"),
    85 => (x"79",x"c1",x"49",x"a6"),
    86 => (x"c4",x"87",x"fd",x"c0"),
    87 => (x"c4",x"4a",x"73",x"83"),
    88 => (x"27",x"1e",x"6a",x"8a"),
    89 => (x"00",x"00",x"17",x"f6"),
    90 => (x"c1",x"86",x"c4",x"0f"),
    91 => (x"87",x"e8",x"c0",x"84"),
    92 => (x"f6",x"27",x"1e",x"6e"),
    93 => (x"0f",x"00",x"00",x"17"),
    94 => (x"db",x"c0",x"86",x"c4"),
    95 => (x"c0",x"49",x"6e",x"87"),
    96 => (x"c0",x"05",x"a9",x"e5"),
    97 => (x"a6",x"c4",x"87",x"c8"),
    98 => (x"c0",x"79",x"c1",x"49"),
    99 => (x"1e",x"6e",x"87",x"ca"),
   100 => (x"00",x"17",x"f6",x"27"),
   101 => (x"86",x"c4",x"0f",x"00"),
   102 => (x"4a",x"66",x"e4",x"c0"),
   103 => (x"48",x"66",x"e4",x"c0"),
   104 => (x"e8",x"c0",x"80",x"c1"),
   105 => (x"48",x"12",x"58",x"a6"),
   106 => (x"c0",x"c0",x"c0",x"c1"),
   107 => (x"c0",x"c4",x"90",x"c0"),
   108 => (x"c4",x"48",x"90",x"b7"),
   109 => (x"05",x"6e",x"58",x"a6"),
   110 => (x"74",x"87",x"fe",x"fa"),
   111 => (x"26",x"86",x"d0",x"48"),
   112 => (x"26",x"4c",x"26",x"4d"),
   113 => (x"26",x"4a",x"26",x"4b"),
   114 => (x"5a",x"5e",x"0e",x"4f"),
   115 => (x"66",x"cc",x"0e",x"5b"),
   116 => (x"c3",x"2a",x"d8",x"4a"),
   117 => (x"66",x"cc",x"9a",x"ff"),
   118 => (x"cf",x"2b",x"c8",x"4b"),
   119 => (x"72",x"9b",x"c0",x"fc"),
   120 => (x"cc",x"b2",x"73",x"4a"),
   121 => (x"33",x"c8",x"4b",x"66"),
   122 => (x"c0",x"f0",x"ff",x"c0"),
   123 => (x"4a",x"72",x"9b",x"c0"),
   124 => (x"66",x"cc",x"b2",x"73"),
   125 => (x"cf",x"33",x"d8",x"4b"),
   126 => (x"c0",x"c0",x"c0",x"fc"),
   127 => (x"73",x"4a",x"72",x"9b"),
   128 => (x"26",x"48",x"72",x"b2"),
   129 => (x"26",x"4a",x"26",x"4b"),
   130 => (x"5a",x"5e",x"0e",x"4f"),
   131 => (x"66",x"cc",x"0e",x"5b"),
   132 => (x"c3",x"2a",x"c8",x"4a"),
   133 => (x"66",x"cc",x"9a",x"ff"),
   134 => (x"cf",x"33",x"c8",x"4b"),
   135 => (x"72",x"9b",x"c0",x"fc"),
   136 => (x"72",x"b2",x"73",x"4a"),
   137 => (x"26",x"4b",x"26",x"48"),
   138 => (x"0e",x"4f",x"26",x"4a"),
   139 => (x"0e",x"5b",x"5a",x"5e"),
   140 => (x"d0",x"4a",x"66",x"cc"),
   141 => (x"ff",x"ff",x"cf",x"2a"),
   142 => (x"4b",x"66",x"cc",x"9a"),
   143 => (x"c0",x"f0",x"33",x"d0"),
   144 => (x"4a",x"72",x"9b",x"c0"),
   145 => (x"48",x"72",x"b2",x"73"),
   146 => (x"4a",x"26",x"4b",x"26"),
   147 => (x"27",x"1e",x"4f",x"26"),
   148 => (x"10",x"00",x"00",x"00"),
   149 => (x"87",x"fd",x"ff",x"0f"),
   150 => (x"72",x"1e",x"4f",x"26"),
   151 => (x"4a",x"66",x"cc",x"1e"),
   152 => (x"c0",x"9a",x"df",x"c3"),
   153 => (x"b7",x"c0",x"8a",x"f7"),
   154 => (x"c3",x"c0",x"03",x"aa"),
   155 => (x"82",x"e7",x"c0",x"87"),
   156 => (x"c4",x"48",x"66",x"c8"),
   157 => (x"58",x"a6",x"cc",x"30"),
   158 => (x"72",x"48",x"66",x"c8"),
   159 => (x"58",x"a6",x"cc",x"b0"),
   160 => (x"26",x"48",x"66",x"c8"),
   161 => (x"0e",x"4f",x"26",x"4a"),
   162 => (x"5c",x"5b",x"5a",x"5e"),
   163 => (x"f6",x"c0",x"0e",x"5d"),
   164 => (x"4b",x"c0",x"c0",x"e8"),
   165 => (x"00",x"1a",x"a0",x"27"),
   166 => (x"c1",x"48",x"bf",x"00"),
   167 => (x"1a",x"a4",x"27",x"80"),
   168 => (x"97",x"58",x"00",x"00"),
   169 => (x"c1",x"4a",x"66",x"d4"),
   170 => (x"c0",x"c0",x"c0",x"c0"),
   171 => (x"b7",x"c0",x"c4",x"92"),
   172 => (x"d3",x"c1",x"4a",x"92"),
   173 => (x"c0",x"05",x"aa",x"b7"),
   174 => (x"a0",x"27",x"87",x"e6"),
   175 => (x"49",x"00",x"00",x"1a"),
   176 => (x"a4",x"27",x"79",x"c0"),
   177 => (x"49",x"00",x"00",x"1a"),
   178 => (x"ac",x"27",x"79",x"c0"),
   179 => (x"49",x"00",x"00",x"1a"),
   180 => (x"b0",x"27",x"79",x"c0"),
   181 => (x"49",x"00",x"00",x"1a"),
   182 => (x"d3",x"c1",x"79",x"c0"),
   183 => (x"87",x"ef",x"c9",x"7b"),
   184 => (x"00",x"1a",x"a0",x"27"),
   185 => (x"c1",x"49",x"bf",x"00"),
   186 => (x"c1",x"05",x"a9",x"b7"),
   187 => (x"f4",x"c1",x"87",x"d5"),
   188 => (x"66",x"d4",x"97",x"7b"),
   189 => (x"c0",x"c0",x"c1",x"4a"),
   190 => (x"c4",x"92",x"c0",x"c0"),
   191 => (x"4a",x"92",x"b7",x"c0"),
   192 => (x"b0",x"27",x"1e",x"72"),
   193 => (x"bf",x"00",x"00",x"1a"),
   194 => (x"02",x"5a",x"27",x"1e"),
   195 => (x"c8",x"0f",x"00",x"00"),
   196 => (x"1a",x"b4",x"27",x"86"),
   197 => (x"27",x"58",x"00",x"00"),
   198 => (x"00",x"00",x"1a",x"b0"),
   199 => (x"b7",x"c3",x"4d",x"bf"),
   200 => (x"c6",x"c0",x"06",x"ad"),
   201 => (x"75",x"48",x"ca",x"87"),
   202 => (x"75",x"4d",x"70",x"88"),
   203 => (x"72",x"82",x"c1",x"4a"),
   204 => (x"27",x"30",x"c1",x"48"),
   205 => (x"00",x"00",x"1a",x"ac"),
   206 => (x"c0",x"48",x"75",x"58"),
   207 => (x"7b",x"70",x"80",x"f0"),
   208 => (x"27",x"87",x"cc",x"c8"),
   209 => (x"00",x"00",x"1a",x"b0"),
   210 => (x"b7",x"c9",x"49",x"bf"),
   211 => (x"fe",x"c7",x"01",x"a9"),
   212 => (x"1a",x"b0",x"27",x"87"),
   213 => (x"49",x"bf",x"00",x"00"),
   214 => (x"06",x"a9",x"b7",x"c0"),
   215 => (x"27",x"87",x"f0",x"c7"),
   216 => (x"00",x"00",x"1a",x"b0"),
   217 => (x"f0",x"c0",x"48",x"bf"),
   218 => (x"27",x"7b",x"70",x"80"),
   219 => (x"00",x"00",x"1a",x"a0"),
   220 => (x"b7",x"c3",x"49",x"bf"),
   221 => (x"e9",x"c0",x"01",x"a9"),
   222 => (x"66",x"d4",x"97",x"87"),
   223 => (x"c0",x"c0",x"c1",x"4a"),
   224 => (x"c4",x"92",x"c0",x"c0"),
   225 => (x"4a",x"92",x"b7",x"c0"),
   226 => (x"ac",x"27",x"1e",x"72"),
   227 => (x"bf",x"00",x"00",x"1a"),
   228 => (x"02",x"5a",x"27",x"1e"),
   229 => (x"c8",x"0f",x"00",x"00"),
   230 => (x"1a",x"b0",x"27",x"86"),
   231 => (x"c6",x"58",x"00",x"00"),
   232 => (x"a8",x"27",x"87",x"ed"),
   233 => (x"bf",x"00",x"00",x"1a"),
   234 => (x"27",x"82",x"c3",x"4a"),
   235 => (x"00",x"00",x"1a",x"a0"),
   236 => (x"b7",x"72",x"49",x"bf"),
   237 => (x"f1",x"c0",x"01",x"a9"),
   238 => (x"66",x"d4",x"97",x"87"),
   239 => (x"c0",x"c0",x"c1",x"4a"),
   240 => (x"c4",x"92",x"c0",x"c0"),
   241 => (x"4a",x"92",x"b7",x"c0"),
   242 => (x"a4",x"27",x"1e",x"72"),
   243 => (x"bf",x"00",x"00",x"1a"),
   244 => (x"02",x"5a",x"27",x"1e"),
   245 => (x"c8",x"0f",x"00",x"00"),
   246 => (x"1a",x"a8",x"27",x"86"),
   247 => (x"27",x"58",x"00",x"00"),
   248 => (x"00",x"00",x"1a",x"b4"),
   249 => (x"c5",x"79",x"c1",x"49"),
   250 => (x"b0",x"27",x"87",x"e5"),
   251 => (x"bf",x"00",x"00",x"1a"),
   252 => (x"a9",x"b7",x"c0",x"49"),
   253 => (x"87",x"d0",x"c3",x"06"),
   254 => (x"00",x"1a",x"b0",x"27"),
   255 => (x"c3",x"49",x"bf",x"00"),
   256 => (x"c3",x"01",x"a9",x"b7"),
   257 => (x"ac",x"27",x"87",x"c2"),
   258 => (x"bf",x"00",x"00",x"1a"),
   259 => (x"c1",x"32",x"c1",x"4a"),
   260 => (x"1a",x"a0",x"27",x"82"),
   261 => (x"49",x"bf",x"00",x"00"),
   262 => (x"01",x"a9",x"b7",x"72"),
   263 => (x"97",x"87",x"c2",x"c2"),
   264 => (x"c1",x"4a",x"66",x"d4"),
   265 => (x"c0",x"c0",x"c0",x"c0"),
   266 => (x"b7",x"c0",x"c4",x"92"),
   267 => (x"1e",x"72",x"4a",x"92"),
   268 => (x"00",x"1a",x"b8",x"27"),
   269 => (x"27",x"1e",x"bf",x"00"),
   270 => (x"00",x"00",x"02",x"5a"),
   271 => (x"27",x"86",x"c8",x"0f"),
   272 => (x"00",x"00",x"1a",x"bc"),
   273 => (x"1a",x"b4",x"27",x"58"),
   274 => (x"4a",x"bf",x"00",x"00"),
   275 => (x"b4",x"27",x"8a",x"c1"),
   276 => (x"49",x"00",x"00",x"1a"),
   277 => (x"b7",x"c0",x"79",x"72"),
   278 => (x"f2",x"c3",x"03",x"aa"),
   279 => (x"1a",x"a4",x"27",x"87"),
   280 => (x"4a",x"bf",x"00",x"00"),
   281 => (x"00",x"1a",x"b8",x"27"),
   282 => (x"52",x"bf",x"97",x"00"),
   283 => (x"00",x"1a",x"a4",x"27"),
   284 => (x"c1",x"4a",x"bf",x"00"),
   285 => (x"1a",x"a4",x"27",x"82"),
   286 => (x"72",x"49",x"00",x"00"),
   287 => (x"1a",x"bc",x"27",x"79"),
   288 => (x"b7",x"bf",x"00",x"00"),
   289 => (x"cd",x"c0",x"06",x"aa"),
   290 => (x"1a",x"bc",x"27",x"87"),
   291 => (x"27",x"49",x"00",x"00"),
   292 => (x"00",x"00",x"1a",x"a4"),
   293 => (x"b4",x"27",x"79",x"bf"),
   294 => (x"49",x"00",x"00",x"1a"),
   295 => (x"ee",x"c2",x"79",x"c1"),
   296 => (x"1a",x"b4",x"27",x"87"),
   297 => (x"05",x"bf",x"00",x"00"),
   298 => (x"27",x"87",x"e4",x"c2"),
   299 => (x"00",x"00",x"1a",x"b8"),
   300 => (x"32",x"c4",x"4a",x"bf"),
   301 => (x"00",x"1a",x"b8",x"27"),
   302 => (x"79",x"72",x"49",x"00"),
   303 => (x"00",x"1a",x"a4",x"27"),
   304 => (x"72",x"49",x"bf",x"00"),
   305 => (x"87",x"c7",x"c2",x"51"),
   306 => (x"00",x"1a",x"b0",x"27"),
   307 => (x"c7",x"49",x"bf",x"00"),
   308 => (x"c1",x"04",x"a9",x"b7"),
   309 => (x"4c",x"c0",x"87",x"ed"),
   310 => (x"c1",x"49",x"f4",x"fe"),
   311 => (x"1a",x"a4",x"27",x"79"),
   312 => (x"27",x"49",x"00",x"00"),
   313 => (x"10",x"00",x"00",x"00"),
   314 => (x"00",x"00",x"27",x"79"),
   315 => (x"27",x"49",x"10",x"00"),
   316 => (x"00",x"00",x"1a",x"bc"),
   317 => (x"03",x"a9",x"b7",x"bf"),
   318 => (x"27",x"87",x"e5",x"c0"),
   319 => (x"00",x"00",x"1a",x"a4"),
   320 => (x"27",x"84",x"bf",x"bf"),
   321 => (x"00",x"00",x"1a",x"a4"),
   322 => (x"82",x"c4",x"4a",x"bf"),
   323 => (x"00",x"1a",x"a4",x"27"),
   324 => (x"79",x"72",x"49",x"00"),
   325 => (x"00",x"1a",x"bc",x"27"),
   326 => (x"aa",x"b7",x"bf",x"00"),
   327 => (x"87",x"db",x"ff",x"04"),
   328 => (x"bc",x"27",x"1e",x"74"),
   329 => (x"bf",x"00",x"00",x"1a"),
   330 => (x"18",x"f0",x"27",x"1e"),
   331 => (x"27",x"1e",x"00",x"00"),
   332 => (x"00",x"00",x"00",x"42"),
   333 => (x"c1",x"86",x"cc",x"0f"),
   334 => (x"00",x"27",x"7b",x"c2"),
   335 => (x"0f",x"10",x"00",x"00"),
   336 => (x"27",x"87",x"cc",x"c0"),
   337 => (x"00",x"00",x"1a",x"b0"),
   338 => (x"f0",x"c0",x"48",x"bf"),
   339 => (x"26",x"7b",x"70",x"80"),
   340 => (x"26",x"4c",x"26",x"4d"),
   341 => (x"26",x"4a",x"26",x"4b"),
   342 => (x"5a",x"5e",x"0e",x"4f"),
   343 => (x"0e",x"5d",x"5c",x"5b"),
   344 => (x"c0",x"4d",x"66",x"d8"),
   345 => (x"4a",x"66",x"d4",x"4c"),
   346 => (x"72",x"2a",x"b7",x"dc"),
   347 => (x"d4",x"9b",x"cf",x"4b"),
   348 => (x"30",x"c4",x"48",x"66"),
   349 => (x"c9",x"58",x"a6",x"d8"),
   350 => (x"c0",x"06",x"ab",x"b7"),
   351 => (x"f7",x"c0",x"87",x"c6"),
   352 => (x"87",x"c3",x"c0",x"83"),
   353 => (x"73",x"83",x"f0",x"c0"),
   354 => (x"85",x"c1",x"7d",x"97"),
   355 => (x"b7",x"c8",x"84",x"c1"),
   356 => (x"d0",x"ff",x"04",x"ac"),
   357 => (x"26",x"4d",x"26",x"87"),
   358 => (x"26",x"4b",x"26",x"4c"),
   359 => (x"0e",x"4f",x"26",x"4a"),
   360 => (x"5c",x"5b",x"5a",x"5e"),
   361 => (x"8e",x"d0",x"0e",x"5d"),
   362 => (x"00",x"07",x"b0",x"27"),
   363 => (x"25",x"27",x"1e",x"00"),
   364 => (x"0f",x"00",x"00",x"18"),
   365 => (x"59",x"27",x"86",x"c4"),
   366 => (x"0f",x"00",x"00",x"16"),
   367 => (x"9a",x"72",x"4a",x"70"),
   368 => (x"87",x"fb",x"c4",x"02"),
   369 => (x"00",x"07",x"99",x"27"),
   370 => (x"25",x"27",x"1e",x"00"),
   371 => (x"0f",x"00",x"00",x"18"),
   372 => (x"37",x"27",x"86",x"c4"),
   373 => (x"0f",x"00",x"00",x"08"),
   374 => (x"9a",x"72",x"4a",x"70"),
   375 => (x"87",x"d1",x"c4",x"02"),
   376 => (x"00",x"00",x"00",x"27"),
   377 => (x"71",x"27",x"1e",x"10"),
   378 => (x"1e",x"00",x"00",x"07"),
   379 => (x"00",x"0f",x"59",x"27"),
   380 => (x"86",x"c8",x"0f",x"00"),
   381 => (x"9b",x"73",x"4b",x"70"),
   382 => (x"87",x"c3",x"c4",x"02"),
   383 => (x"c0",x"49",x"a6",x"c8"),
   384 => (x"49",x"a6",x"c4",x"79"),
   385 => (x"00",x"00",x"00",x"27"),
   386 => (x"a6",x"cc",x"79",x"10"),
   387 => (x"c3",x"79",x"c0",x"49"),
   388 => (x"27",x"9b",x"fc",x"83"),
   389 => (x"10",x"00",x"00",x"00"),
   390 => (x"75",x"85",x"73",x"4d"),
   391 => (x"07",x"65",x"27",x"1e"),
   392 => (x"27",x"1e",x"00",x"00"),
   393 => (x"00",x"00",x"0f",x"59"),
   394 => (x"70",x"86",x"c8",x"0f"),
   395 => (x"02",x"9a",x"72",x"4a"),
   396 => (x"c7",x"87",x"e0",x"c2"),
   397 => (x"06",x"ab",x"b7",x"ff"),
   398 => (x"c8",x"87",x"d8",x"c2"),
   399 => (x"66",x"c8",x"1e",x"c0"),
   400 => (x"82",x"66",x"d0",x"4a"),
   401 => (x"59",x"27",x"1e",x"72"),
   402 => (x"0f",x"00",x"00",x"18"),
   403 => (x"4a",x"70",x"86",x"c8"),
   404 => (x"49",x"76",x"4c",x"72"),
   405 => (x"66",x"cc",x"79",x"25"),
   406 => (x"80",x"c0",x"c8",x"48"),
   407 => (x"c8",x"58",x"a6",x"d0"),
   408 => (x"b7",x"6e",x"8b",x"c0"),
   409 => (x"e2",x"c1",x"02",x"ac"),
   410 => (x"48",x"66",x"c8",x"87"),
   411 => (x"a6",x"cc",x"80",x"c1"),
   412 => (x"1a",x"80",x"27",x"58"),
   413 => (x"d0",x"1e",x"00",x"00"),
   414 => (x"59",x"27",x"1e",x"66"),
   415 => (x"0f",x"00",x"00",x"05"),
   416 => (x"88",x"27",x"86",x"c8"),
   417 => (x"49",x"00",x"00",x"1a"),
   418 => (x"27",x"51",x"e0",x"c0"),
   419 => (x"00",x"00",x"1a",x"89"),
   420 => (x"27",x"1e",x"74",x"1e"),
   421 => (x"00",x"00",x"05",x"59"),
   422 => (x"27",x"86",x"c8",x"0f"),
   423 => (x"00",x"00",x"1a",x"91"),
   424 => (x"51",x"e0",x"c0",x"49"),
   425 => (x"00",x"1a",x"92",x"27"),
   426 => (x"66",x"c4",x"1e",x"00"),
   427 => (x"05",x"59",x"27",x"1e"),
   428 => (x"c8",x"0f",x"00",x"00"),
   429 => (x"1a",x"9a",x"27",x"86"),
   430 => (x"c0",x"49",x"00",x"00"),
   431 => (x"1a",x"80",x"27",x"51"),
   432 => (x"27",x"1e",x"00",x"00"),
   433 => (x"00",x"00",x"10",x"c4"),
   434 => (x"c7",x"86",x"c4",x"0f"),
   435 => (x"01",x"ab",x"b7",x"ff"),
   436 => (x"c8",x"87",x"e8",x"fd"),
   437 => (x"e6",x"c0",x"05",x"66"),
   438 => (x"00",x"00",x"27",x"87"),
   439 => (x"bf",x"97",x"10",x"00"),
   440 => (x"c0",x"c0",x"c1",x"4a"),
   441 => (x"c4",x"92",x"c0",x"c0"),
   442 => (x"4a",x"92",x"b7",x"c0"),
   443 => (x"ce",x"c0",x"0f",x"72"),
   444 => (x"07",x"7d",x"27",x"87"),
   445 => (x"27",x"1e",x"00",x"00"),
   446 => (x"00",x"00",x"18",x"25"),
   447 => (x"27",x"86",x"c4",x"0f"),
   448 => (x"00",x"00",x"07",x"c6"),
   449 => (x"18",x"25",x"27",x"1e"),
   450 => (x"c4",x"0f",x"00",x"00"),
   451 => (x"1a",x"bc",x"27",x"86"),
   452 => (x"c0",x"49",x"00",x"00"),
   453 => (x"e8",x"f6",x"c0",x"79"),
   454 => (x"c0",x"4d",x"c0",x"c0"),
   455 => (x"f6",x"27",x"1e",x"ee"),
   456 => (x"0f",x"00",x"00",x"17"),
   457 => (x"f4",x"c3",x"86",x"c4"),
   458 => (x"6d",x"4b",x"ff",x"c8"),
   459 => (x"c8",x"4a",x"74",x"4c"),
   460 => (x"9a",x"72",x"9a",x"c0"),
   461 => (x"87",x"d4",x"c0",x"02"),
   462 => (x"ff",x"c3",x"4a",x"74"),
   463 => (x"27",x"1e",x"72",x"9a"),
   464 => (x"00",x"00",x"02",x"87"),
   465 => (x"c3",x"86",x"c4",x"0f"),
   466 => (x"4b",x"c0",x"c9",x"f4"),
   467 => (x"8b",x"c1",x"4a",x"73"),
   468 => (x"ff",x"05",x"9a",x"72"),
   469 => (x"c2",x"ff",x"87",x"d5"),
   470 => (x"26",x"86",x"d0",x"87"),
   471 => (x"26",x"4c",x"26",x"4d"),
   472 => (x"26",x"4a",x"26",x"4b"),
   473 => (x"45",x"48",x"43",x"4f"),
   474 => (x"55",x"53",x"4b",x"43"),
   475 => (x"4e",x"49",x"42",x"4d"),
   476 => (x"44",x"53",x"4f",x"00"),
   477 => (x"30",x"32",x"33",x"38"),
   478 => (x"53",x"59",x"53",x"31"),
   479 => (x"61",x"6e",x"55",x"00"),
   480 => (x"20",x"65",x"6c",x"62"),
   481 => (x"6c",x"20",x"6f",x"74"),
   482 => (x"74",x"61",x"63",x"6f"),
   483 => (x"61",x"70",x"20",x"65"),
   484 => (x"74",x"69",x"74",x"72"),
   485 => (x"0a",x"6e",x"6f",x"69"),
   486 => (x"6e",x"75",x"48",x"00"),
   487 => (x"67",x"6e",x"69",x"74"),
   488 => (x"72",x"6f",x"66",x"20"),
   489 => (x"72",x"61",x"70",x"20"),
   490 => (x"69",x"74",x"69",x"74"),
   491 => (x"00",x"0a",x"6e",x"6f"),
   492 => (x"74",x"69",x"6e",x"49"),
   493 => (x"69",x"6c",x"61",x"69"),
   494 => (x"67",x"6e",x"69",x"7a"),
   495 => (x"20",x"44",x"53",x"20"),
   496 => (x"64",x"72",x"61",x"63"),
   497 => (x"6f",x"42",x"00",x"0a"),
   498 => (x"6e",x"69",x"74",x"6f"),
   499 => (x"72",x"66",x"20",x"67"),
   500 => (x"52",x"20",x"6d",x"6f"),
   501 => (x"32",x"33",x"32",x"53"),
   502 => (x"5e",x"0e",x"00",x"2e"),
   503 => (x"5d",x"5c",x"5b",x"5a"),
   504 => (x"4d",x"66",x"d4",x"0e"),
   505 => (x"66",x"dc",x"4c",x"c0"),
   506 => (x"a9",x"b7",x"c0",x"49"),
   507 => (x"87",x"fb",x"c0",x"06"),
   508 => (x"c0",x"c1",x"4b",x"15"),
   509 => (x"93",x"c0",x"c0",x"c0"),
   510 => (x"93",x"b7",x"c0",x"c4"),
   511 => (x"97",x"66",x"d8",x"4b"),
   512 => (x"c0",x"c1",x"4a",x"bf"),
   513 => (x"92",x"c0",x"c0",x"c0"),
   514 => (x"92",x"b7",x"c0",x"c4"),
   515 => (x"48",x"66",x"d8",x"4a"),
   516 => (x"a6",x"dc",x"80",x"c1"),
   517 => (x"ab",x"b7",x"72",x"58"),
   518 => (x"87",x"c5",x"c0",x"02"),
   519 => (x"cc",x"c0",x"48",x"c1"),
   520 => (x"dc",x"84",x"c1",x"87"),
   521 => (x"04",x"ac",x"b7",x"66"),
   522 => (x"c0",x"87",x"c5",x"ff"),
   523 => (x"26",x"4d",x"26",x"48"),
   524 => (x"26",x"4b",x"26",x"4c"),
   525 => (x"0e",x"4f",x"26",x"4a"),
   526 => (x"5c",x"5b",x"5a",x"5e"),
   527 => (x"c8",x"27",x"0e",x"5d"),
   528 => (x"49",x"00",x"00",x"1c"),
   529 => (x"d8",x"27",x"79",x"c0"),
   530 => (x"1e",x"00",x"00",x"19"),
   531 => (x"00",x"18",x"25",x"27"),
   532 => (x"86",x"c4",x"0f",x"00"),
   533 => (x"00",x"1a",x"c0",x"27"),
   534 => (x"1e",x"c0",x"1e",x"00"),
   535 => (x"00",x"16",x"fa",x"27"),
   536 => (x"86",x"c8",x"0f",x"00"),
   537 => (x"9a",x"72",x"4a",x"70"),
   538 => (x"87",x"d3",x"c0",x"05"),
   539 => (x"00",x"19",x"04",x"27"),
   540 => (x"25",x"27",x"1e",x"00"),
   541 => (x"0f",x"00",x"00",x"18"),
   542 => (x"48",x"c0",x"86",x"c4"),
   543 => (x"27",x"87",x"e6",x"d0"),
   544 => (x"00",x"00",x"19",x"e5"),
   545 => (x"18",x"25",x"27",x"1e"),
   546 => (x"c4",x"0f",x"00",x"00"),
   547 => (x"27",x"4c",x"c0",x"86"),
   548 => (x"00",x"00",x"1c",x"f4"),
   549 => (x"c8",x"79",x"c1",x"49"),
   550 => (x"19",x"fc",x"27",x"1e"),
   551 => (x"27",x"1e",x"00",x"00"),
   552 => (x"00",x"00",x"1a",x"f6"),
   553 => (x"07",x"da",x"27",x"1e"),
   554 => (x"cc",x"0f",x"00",x"00"),
   555 => (x"72",x"4a",x"70",x"86"),
   556 => (x"c8",x"c0",x"05",x"9a"),
   557 => (x"1c",x"f4",x"27",x"87"),
   558 => (x"c0",x"49",x"00",x"00"),
   559 => (x"27",x"1e",x"c8",x"79"),
   560 => (x"00",x"00",x"1a",x"05"),
   561 => (x"1b",x"12",x"27",x"1e"),
   562 => (x"27",x"1e",x"00",x"00"),
   563 => (x"00",x"00",x"07",x"da"),
   564 => (x"70",x"86",x"cc",x"0f"),
   565 => (x"05",x"9a",x"72",x"4a"),
   566 => (x"27",x"87",x"c8",x"c0"),
   567 => (x"00",x"00",x"1c",x"f4"),
   568 => (x"27",x"79",x"c0",x"49"),
   569 => (x"00",x"00",x"1c",x"f4"),
   570 => (x"0e",x"27",x"1e",x"bf"),
   571 => (x"1e",x"00",x"00",x"1a"),
   572 => (x"00",x"00",x"42",x"27"),
   573 => (x"86",x"c8",x"0f",x"00"),
   574 => (x"00",x"1c",x"f4",x"27"),
   575 => (x"c3",x"02",x"bf",x"00"),
   576 => (x"c0",x"27",x"87",x"cc"),
   577 => (x"4d",x"00",x"00",x"1a"),
   578 => (x"00",x"1c",x"7e",x"27"),
   579 => (x"be",x"27",x"4b",x"00"),
   580 => (x"9f",x"00",x"00",x"1c"),
   581 => (x"ff",x"cf",x"4a",x"bf"),
   582 => (x"1e",x"72",x"9a",x"ff"),
   583 => (x"00",x"1c",x"be",x"27"),
   584 => (x"c0",x"27",x"4a",x"00"),
   585 => (x"8a",x"00",x"00",x"1a"),
   586 => (x"1e",x"d0",x"1e",x"72"),
   587 => (x"27",x"1e",x"c0",x"c8"),
   588 => (x"00",x"00",x"19",x"36"),
   589 => (x"00",x"42",x"27",x"1e"),
   590 => (x"d4",x"0f",x"00",x"00"),
   591 => (x"c8",x"4a",x"73",x"86"),
   592 => (x"27",x"4c",x"6a",x"82"),
   593 => (x"00",x"00",x"1c",x"be"),
   594 => (x"cf",x"4a",x"bf",x"9f"),
   595 => (x"c5",x"9a",x"ff",x"ff"),
   596 => (x"aa",x"b7",x"ea",x"d6"),
   597 => (x"87",x"d3",x"c0",x"05"),
   598 => (x"82",x"c8",x"4a",x"73"),
   599 => (x"c9",x"27",x"1e",x"6a"),
   600 => (x"0f",x"00",x"00",x"01"),
   601 => (x"4c",x"70",x"86",x"c4"),
   602 => (x"75",x"87",x"e8",x"c0"),
   603 => (x"82",x"fe",x"c7",x"4a"),
   604 => (x"cf",x"4a",x"6a",x"9f"),
   605 => (x"ca",x"9a",x"ff",x"ff"),
   606 => (x"aa",x"b7",x"d5",x"e9"),
   607 => (x"87",x"d3",x"c0",x"02"),
   608 => (x"00",x"19",x"18",x"27"),
   609 => (x"25",x"27",x"1e",x"00"),
   610 => (x"0f",x"00",x"00",x"18"),
   611 => (x"48",x"c0",x"86",x"c4"),
   612 => (x"74",x"87",x"d2",x"cc"),
   613 => (x"19",x"73",x"27",x"1e"),
   614 => (x"27",x"1e",x"00",x"00"),
   615 => (x"00",x"00",x"00",x"42"),
   616 => (x"27",x"86",x"c8",x"0f"),
   617 => (x"00",x"00",x"1a",x"c0"),
   618 => (x"27",x"1e",x"74",x"1e"),
   619 => (x"00",x"00",x"16",x"fa"),
   620 => (x"70",x"86",x"c8",x"0f"),
   621 => (x"05",x"9a",x"72",x"4a"),
   622 => (x"c0",x"87",x"c5",x"c0"),
   623 => (x"87",x"e5",x"cb",x"48"),
   624 => (x"00",x"19",x"8b",x"27"),
   625 => (x"25",x"27",x"1e",x"00"),
   626 => (x"0f",x"00",x"00",x"18"),
   627 => (x"21",x"27",x"86",x"c4"),
   628 => (x"1e",x"00",x"00",x"1a"),
   629 => (x"00",x"00",x"42",x"27"),
   630 => (x"86",x"c4",x"0f",x"00"),
   631 => (x"39",x"27",x"1e",x"c8"),
   632 => (x"1e",x"00",x"00",x"1a"),
   633 => (x"00",x"1b",x"12",x"27"),
   634 => (x"da",x"27",x"1e",x"00"),
   635 => (x"0f",x"00",x"00",x"07"),
   636 => (x"4a",x"70",x"86",x"cc"),
   637 => (x"c0",x"05",x"9a",x"72"),
   638 => (x"c8",x"27",x"87",x"cb"),
   639 => (x"49",x"00",x"00",x"1c"),
   640 => (x"f1",x"c0",x"79",x"c1"),
   641 => (x"27",x"1e",x"c8",x"87"),
   642 => (x"00",x"00",x"1a",x"42"),
   643 => (x"1a",x"f6",x"27",x"1e"),
   644 => (x"27",x"1e",x"00",x"00"),
   645 => (x"00",x"00",x"07",x"da"),
   646 => (x"70",x"86",x"cc",x"0f"),
   647 => (x"02",x"9a",x"72",x"4a"),
   648 => (x"27",x"87",x"d3",x"c0"),
   649 => (x"00",x"00",x"19",x"b2"),
   650 => (x"00",x"42",x"27",x"1e"),
   651 => (x"c4",x"0f",x"00",x"00"),
   652 => (x"c9",x"48",x"c0",x"86"),
   653 => (x"be",x"27",x"87",x"ef"),
   654 => (x"97",x"00",x"00",x"1c"),
   655 => (x"ff",x"c3",x"4a",x"bf"),
   656 => (x"b7",x"d5",x"c1",x"9a"),
   657 => (x"d3",x"c0",x"05",x"aa"),
   658 => (x"1c",x"bf",x"27",x"87"),
   659 => (x"bf",x"97",x"00",x"00"),
   660 => (x"9a",x"ff",x"c3",x"4a"),
   661 => (x"aa",x"b7",x"ea",x"c2"),
   662 => (x"87",x"c5",x"c0",x"02"),
   663 => (x"c4",x"c9",x"48",x"c0"),
   664 => (x"1a",x"c0",x"27",x"87"),
   665 => (x"bf",x"97",x"00",x"00"),
   666 => (x"9a",x"ff",x"c3",x"4a"),
   667 => (x"aa",x"b7",x"e9",x"c3"),
   668 => (x"87",x"d8",x"c0",x"02"),
   669 => (x"00",x"1a",x"c0",x"27"),
   670 => (x"4a",x"bf",x"97",x"00"),
   671 => (x"c3",x"9a",x"ff",x"c3"),
   672 => (x"02",x"aa",x"b7",x"eb"),
   673 => (x"c0",x"87",x"c5",x"c0"),
   674 => (x"87",x"d9",x"c8",x"48"),
   675 => (x"00",x"1a",x"cb",x"27"),
   676 => (x"4a",x"bf",x"97",x"00"),
   677 => (x"72",x"9a",x"ff",x"c3"),
   678 => (x"d2",x"c0",x"05",x"9a"),
   679 => (x"1a",x"cc",x"27",x"87"),
   680 => (x"bf",x"97",x"00",x"00"),
   681 => (x"9a",x"ff",x"c3",x"4a"),
   682 => (x"02",x"aa",x"b7",x"c2"),
   683 => (x"c0",x"87",x"c5",x"c0"),
   684 => (x"87",x"f1",x"c7",x"48"),
   685 => (x"00",x"1a",x"cd",x"27"),
   686 => (x"48",x"bf",x"97",x"00"),
   687 => (x"27",x"98",x"ff",x"c3"),
   688 => (x"00",x"00",x"1c",x"c4"),
   689 => (x"1c",x"c0",x"27",x"58"),
   690 => (x"4a",x"bf",x"00",x"00"),
   691 => (x"8b",x"c1",x"4b",x"72"),
   692 => (x"00",x"1c",x"c4",x"27"),
   693 => (x"79",x"73",x"49",x"00"),
   694 => (x"1e",x"72",x"1e",x"73"),
   695 => (x"00",x"1a",x"4b",x"27"),
   696 => (x"42",x"27",x"1e",x"00"),
   697 => (x"0f",x"00",x"00",x"00"),
   698 => (x"ce",x"27",x"86",x"cc"),
   699 => (x"97",x"00",x"00",x"1a"),
   700 => (x"ff",x"c3",x"4a",x"bf"),
   701 => (x"27",x"82",x"74",x"9a"),
   702 => (x"00",x"00",x"1a",x"cf"),
   703 => (x"c3",x"4b",x"bf",x"97"),
   704 => (x"33",x"c8",x"9b",x"ff"),
   705 => (x"80",x"72",x"48",x"73"),
   706 => (x"00",x"1c",x"d8",x"27"),
   707 => (x"d0",x"27",x"58",x"00"),
   708 => (x"97",x"00",x"00",x"1a"),
   709 => (x"ff",x"c3",x"48",x"bf"),
   710 => (x"1c",x"ec",x"27",x"98"),
   711 => (x"27",x"58",x"00",x"00"),
   712 => (x"00",x"00",x"1c",x"c8"),
   713 => (x"f7",x"c3",x"02",x"bf"),
   714 => (x"27",x"1e",x"c8",x"87"),
   715 => (x"00",x"00",x"19",x"cf"),
   716 => (x"1b",x"12",x"27",x"1e"),
   717 => (x"27",x"1e",x"00",x"00"),
   718 => (x"00",x"00",x"07",x"da"),
   719 => (x"70",x"86",x"cc",x"0f"),
   720 => (x"02",x"9a",x"72",x"4a"),
   721 => (x"c0",x"87",x"c5",x"c0"),
   722 => (x"87",x"d9",x"c5",x"48"),
   723 => (x"00",x"1c",x"c0",x"27"),
   724 => (x"73",x"4b",x"bf",x"00"),
   725 => (x"27",x"30",x"c4",x"48"),
   726 => (x"00",x"00",x"1c",x"f0"),
   727 => (x"1c",x"e4",x"27",x"58"),
   728 => (x"73",x"49",x"00",x"00"),
   729 => (x"1a",x"e5",x"27",x"79"),
   730 => (x"bf",x"97",x"00",x"00"),
   731 => (x"9a",x"ff",x"c3",x"4a"),
   732 => (x"e4",x"27",x"32",x"c8"),
   733 => (x"97",x"00",x"00",x"1a"),
   734 => (x"ff",x"c3",x"4c",x"bf"),
   735 => (x"74",x"4a",x"72",x"9c"),
   736 => (x"1a",x"e6",x"27",x"82"),
   737 => (x"bf",x"97",x"00",x"00"),
   738 => (x"9c",x"ff",x"c3",x"4c"),
   739 => (x"4a",x"72",x"34",x"d0"),
   740 => (x"e7",x"27",x"82",x"74"),
   741 => (x"97",x"00",x"00",x"1a"),
   742 => (x"ff",x"c3",x"4c",x"bf"),
   743 => (x"72",x"34",x"d8",x"9c"),
   744 => (x"27",x"82",x"74",x"4a"),
   745 => (x"00",x"00",x"1c",x"f0"),
   746 => (x"72",x"79",x"72",x"49"),
   747 => (x"1c",x"e8",x"27",x"4a"),
   748 => (x"92",x"bf",x"00",x"00"),
   749 => (x"d4",x"27",x"4a",x"72"),
   750 => (x"bf",x"00",x"00",x"1c"),
   751 => (x"1c",x"d8",x"27",x"82"),
   752 => (x"72",x"49",x"00",x"00"),
   753 => (x"1a",x"ed",x"27",x"79"),
   754 => (x"bf",x"97",x"00",x"00"),
   755 => (x"9c",x"ff",x"c3",x"4c"),
   756 => (x"ec",x"27",x"34",x"c8"),
   757 => (x"97",x"00",x"00",x"1a"),
   758 => (x"ff",x"c3",x"4d",x"bf"),
   759 => (x"75",x"4c",x"74",x"9d"),
   760 => (x"1a",x"ee",x"27",x"84"),
   761 => (x"bf",x"97",x"00",x"00"),
   762 => (x"9d",x"ff",x"c3",x"4d"),
   763 => (x"4c",x"74",x"35",x"d0"),
   764 => (x"ef",x"27",x"84",x"75"),
   765 => (x"97",x"00",x"00",x"1a"),
   766 => (x"ff",x"c3",x"4d",x"bf"),
   767 => (x"d8",x"9d",x"cf",x"9d"),
   768 => (x"75",x"4c",x"74",x"35"),
   769 => (x"1c",x"dc",x"27",x"84"),
   770 => (x"74",x"49",x"00",x"00"),
   771 => (x"73",x"8c",x"c2",x"79"),
   772 => (x"73",x"93",x"74",x"4b"),
   773 => (x"27",x"80",x"72",x"48"),
   774 => (x"00",x"00",x"1c",x"e4"),
   775 => (x"87",x"c3",x"c2",x"58"),
   776 => (x"00",x"1a",x"d2",x"27"),
   777 => (x"4a",x"bf",x"97",x"00"),
   778 => (x"c8",x"9a",x"ff",x"c3"),
   779 => (x"1a",x"d1",x"27",x"32"),
   780 => (x"bf",x"97",x"00",x"00"),
   781 => (x"9b",x"ff",x"c3",x"4b"),
   782 => (x"82",x"73",x"4a",x"72"),
   783 => (x"00",x"1c",x"ec",x"27"),
   784 => (x"79",x"72",x"49",x"00"),
   785 => (x"ff",x"c7",x"32",x"c5"),
   786 => (x"27",x"2a",x"c9",x"82"),
   787 => (x"00",x"00",x"1c",x"e4"),
   788 => (x"27",x"79",x"72",x"49"),
   789 => (x"00",x"00",x"1a",x"d7"),
   790 => (x"c3",x"4b",x"bf",x"97"),
   791 => (x"33",x"c8",x"9b",x"ff"),
   792 => (x"00",x"1a",x"d6",x"27"),
   793 => (x"4c",x"bf",x"97",x"00"),
   794 => (x"73",x"9c",x"ff",x"c3"),
   795 => (x"27",x"83",x"74",x"4b"),
   796 => (x"00",x"00",x"1c",x"f0"),
   797 => (x"73",x"79",x"73",x"49"),
   798 => (x"1c",x"e8",x"27",x"4b"),
   799 => (x"93",x"bf",x"00",x"00"),
   800 => (x"d4",x"27",x"4b",x"73"),
   801 => (x"bf",x"00",x"00",x"1c"),
   802 => (x"1c",x"e0",x"27",x"83"),
   803 => (x"73",x"49",x"00",x"00"),
   804 => (x"1c",x"dc",x"27",x"79"),
   805 => (x"c0",x"49",x"00",x"00"),
   806 => (x"72",x"48",x"73",x"79"),
   807 => (x"1c",x"dc",x"27",x"80"),
   808 => (x"c1",x"58",x"00",x"00"),
   809 => (x"26",x"4d",x"26",x"48"),
   810 => (x"26",x"4b",x"26",x"4c"),
   811 => (x"0e",x"4f",x"26",x"4a"),
   812 => (x"5c",x"5b",x"5a",x"5e"),
   813 => (x"c8",x"27",x"0e",x"5d"),
   814 => (x"bf",x"00",x"00",x"1c"),
   815 => (x"87",x"cf",x"c0",x"02"),
   816 => (x"c7",x"4d",x"66",x"d4"),
   817 => (x"66",x"d4",x"2d",x"b7"),
   818 => (x"9b",x"ff",x"c1",x"4b"),
   819 => (x"d4",x"87",x"cc",x"c0"),
   820 => (x"b7",x"c8",x"4d",x"66"),
   821 => (x"4b",x"66",x"d4",x"2d"),
   822 => (x"27",x"9b",x"ff",x"c3"),
   823 => (x"00",x"00",x"1a",x"c0"),
   824 => (x"1c",x"d4",x"27",x"1e"),
   825 => (x"4a",x"bf",x"00",x"00"),
   826 => (x"1e",x"72",x"82",x"75"),
   827 => (x"00",x"16",x"fa",x"27"),
   828 => (x"86",x"c8",x"0f",x"00"),
   829 => (x"9a",x"72",x"4a",x"70"),
   830 => (x"87",x"c5",x"c0",x"05"),
   831 => (x"f6",x"c0",x"48",x"c0"),
   832 => (x"1c",x"c8",x"27",x"87"),
   833 => (x"02",x"bf",x"00",x"00"),
   834 => (x"73",x"87",x"d7",x"c0"),
   835 => (x"72",x"92",x"c4",x"4a"),
   836 => (x"1a",x"c0",x"27",x"4a"),
   837 => (x"6a",x"82",x"00",x"00"),
   838 => (x"ff",x"ff",x"cf",x"4c"),
   839 => (x"c0",x"9c",x"ff",x"ff"),
   840 => (x"4a",x"73",x"87",x"d3"),
   841 => (x"4a",x"72",x"92",x"c2"),
   842 => (x"00",x"1a",x"c0",x"27"),
   843 => (x"6a",x"9f",x"82",x"00"),
   844 => (x"ff",x"ff",x"cf",x"4c"),
   845 => (x"26",x"48",x"74",x"9c"),
   846 => (x"26",x"4c",x"26",x"4d"),
   847 => (x"26",x"4a",x"26",x"4b"),
   848 => (x"5a",x"5e",x"0e",x"4f"),
   849 => (x"0e",x"5d",x"5c",x"5b"),
   850 => (x"ff",x"cf",x"8e",x"cc"),
   851 => (x"4d",x"f8",x"ff",x"ff"),
   852 => (x"49",x"76",x"4c",x"c0"),
   853 => (x"00",x"1c",x"dc",x"27"),
   854 => (x"c4",x"79",x"bf",x"00"),
   855 => (x"e0",x"27",x"49",x"a6"),
   856 => (x"bf",x"00",x"00",x"1c"),
   857 => (x"1c",x"c8",x"27",x"79"),
   858 => (x"02",x"bf",x"00",x"00"),
   859 => (x"27",x"87",x"cc",x"c0"),
   860 => (x"00",x"00",x"1c",x"c0"),
   861 => (x"32",x"c4",x"4a",x"bf"),
   862 => (x"27",x"87",x"c9",x"c0"),
   863 => (x"00",x"00",x"1c",x"e4"),
   864 => (x"32",x"c4",x"4a",x"bf"),
   865 => (x"72",x"49",x"a6",x"c8"),
   866 => (x"c8",x"4b",x"c0",x"79"),
   867 => (x"a9",x"c0",x"49",x"66"),
   868 => (x"87",x"e1",x"c3",x"06"),
   869 => (x"9a",x"cf",x"4a",x"73"),
   870 => (x"c0",x"05",x"9a",x"72"),
   871 => (x"c0",x"27",x"87",x"e4"),
   872 => (x"1e",x"00",x"00",x"1a"),
   873 => (x"c8",x"4a",x"66",x"c8"),
   874 => (x"80",x"c1",x"48",x"66"),
   875 => (x"72",x"58",x"a6",x"cc"),
   876 => (x"16",x"fa",x"27",x"1e"),
   877 => (x"c8",x"0f",x"00",x"00"),
   878 => (x"1a",x"c0",x"27",x"86"),
   879 => (x"c0",x"4c",x"00",x"00"),
   880 => (x"e0",x"c0",x"87",x"c3"),
   881 => (x"4a",x"6c",x"97",x"84"),
   882 => (x"72",x"9a",x"ff",x"c3"),
   883 => (x"db",x"c2",x"02",x"9a"),
   884 => (x"4a",x"6c",x"97",x"87"),
   885 => (x"c3",x"9a",x"ff",x"c3"),
   886 => (x"02",x"aa",x"b7",x"e5"),
   887 => (x"74",x"87",x"cd",x"c2"),
   888 => (x"97",x"82",x"cb",x"4a"),
   889 => (x"ff",x"c3",x"4a",x"6a"),
   890 => (x"72",x"9a",x"d8",x"9a"),
   891 => (x"fb",x"c1",x"05",x"9a"),
   892 => (x"27",x"1e",x"74",x"87"),
   893 => (x"00",x"00",x"18",x"25"),
   894 => (x"cb",x"86",x"c4",x"0f"),
   895 => (x"66",x"e8",x"c0",x"1e"),
   896 => (x"27",x"1e",x"74",x"1e"),
   897 => (x"00",x"00",x"07",x"da"),
   898 => (x"70",x"86",x"cc",x"0f"),
   899 => (x"05",x"9a",x"72",x"4a"),
   900 => (x"74",x"87",x"d9",x"c1"),
   901 => (x"c0",x"83",x"dc",x"4b"),
   902 => (x"c4",x"4a",x"66",x"e0"),
   903 => (x"74",x"7a",x"6b",x"82"),
   904 => (x"c0",x"83",x"da",x"4b"),
   905 => (x"c8",x"4a",x"66",x"e0"),
   906 => (x"48",x"6b",x"9f",x"82"),
   907 => (x"98",x"ff",x"ff",x"cf"),
   908 => (x"4d",x"72",x"7a",x"70"),
   909 => (x"00",x"1c",x"c8",x"27"),
   910 => (x"c0",x"02",x"bf",x"00"),
   911 => (x"4a",x"74",x"87",x"d9"),
   912 => (x"6a",x"9f",x"82",x"d4"),
   913 => (x"ff",x"ff",x"cf",x"4a"),
   914 => (x"ff",x"ff",x"c0",x"9a"),
   915 => (x"d0",x"48",x"72",x"9a"),
   916 => (x"58",x"a6",x"c4",x"30"),
   917 => (x"76",x"87",x"c4",x"c0"),
   918 => (x"6e",x"79",x"c0",x"49"),
   919 => (x"70",x"80",x"6d",x"48"),
   920 => (x"66",x"e0",x"c0",x"7d"),
   921 => (x"c1",x"79",x"c0",x"49"),
   922 => (x"87",x"ce",x"c1",x"48"),
   923 => (x"66",x"c8",x"83",x"c1"),
   924 => (x"df",x"fc",x"04",x"ab"),
   925 => (x"ff",x"ff",x"cf",x"87"),
   926 => (x"27",x"4d",x"f8",x"ff"),
   927 => (x"00",x"00",x"1c",x"c8"),
   928 => (x"f3",x"c0",x"02",x"bf"),
   929 => (x"27",x"1e",x"6e",x"87"),
   930 => (x"00",x"00",x"0c",x"af"),
   931 => (x"c4",x"86",x"c4",x"0f"),
   932 => (x"4a",x"6e",x"58",x"a6"),
   933 => (x"aa",x"75",x"9a",x"75"),
   934 => (x"87",x"dc",x"c0",x"02"),
   935 => (x"8a",x"c2",x"4a",x"6e"),
   936 => (x"c0",x"27",x"4a",x"72"),
   937 => (x"bf",x"00",x"00",x"1c"),
   938 => (x"1c",x"d8",x"27",x"92"),
   939 => (x"48",x"bf",x"00",x"00"),
   940 => (x"a6",x"c8",x"80",x"72"),
   941 => (x"87",x"d1",x"fb",x"58"),
   942 => (x"ff",x"cf",x"48",x"c0"),
   943 => (x"4d",x"f8",x"ff",x"ff"),
   944 => (x"4d",x"26",x"86",x"cc"),
   945 => (x"4b",x"26",x"4c",x"26"),
   946 => (x"4f",x"26",x"4a",x"26"),
   947 => (x"5b",x"5a",x"5e",x"0e"),
   948 => (x"bf",x"66",x"cc",x"0e"),
   949 => (x"cc",x"82",x"c1",x"4a"),
   950 => (x"79",x"72",x"49",x"66"),
   951 => (x"c4",x"27",x"4a",x"72"),
   952 => (x"bf",x"00",x"00",x"1c"),
   953 => (x"05",x"9a",x"72",x"9a"),
   954 => (x"cc",x"87",x"d3",x"c0"),
   955 => (x"82",x"c8",x"4a",x"66"),
   956 => (x"af",x"27",x"1e",x"6a"),
   957 => (x"0f",x"00",x"00",x"0c"),
   958 => (x"4b",x"70",x"86",x"c4"),
   959 => (x"48",x"c1",x"7a",x"73"),
   960 => (x"4a",x"26",x"4b",x"26"),
   961 => (x"5e",x"0e",x"4f",x"26"),
   962 => (x"27",x"0e",x"5b",x"5a"),
   963 => (x"00",x"00",x"1c",x"d8"),
   964 => (x"66",x"cc",x"4a",x"bf"),
   965 => (x"6b",x"83",x"c8",x"4b"),
   966 => (x"73",x"8b",x"c2",x"4b"),
   967 => (x"1c",x"c0",x"27",x"4b"),
   968 => (x"93",x"bf",x"00",x"00"),
   969 => (x"82",x"73",x"4a",x"72"),
   970 => (x"00",x"1c",x"c4",x"27"),
   971 => (x"cc",x"4b",x"bf",x"00"),
   972 => (x"72",x"9b",x"bf",x"66"),
   973 => (x"d0",x"82",x"73",x"4a"),
   974 => (x"1e",x"72",x"1e",x"66"),
   975 => (x"00",x"16",x"fa",x"27"),
   976 => (x"86",x"c8",x"0f",x"00"),
   977 => (x"9a",x"72",x"4a",x"70"),
   978 => (x"87",x"c5",x"c0",x"05"),
   979 => (x"c2",x"c0",x"48",x"c0"),
   980 => (x"26",x"48",x"c1",x"87"),
   981 => (x"26",x"4a",x"26",x"4b"),
   982 => (x"5a",x"5e",x"0e",x"4f"),
   983 => (x"0e",x"5d",x"5c",x"5b"),
   984 => (x"d4",x"4c",x"66",x"d8"),
   985 => (x"f8",x"27",x"1e",x"66"),
   986 => (x"1e",x"00",x"00",x"1c"),
   987 => (x"00",x"0d",x"41",x"27"),
   988 => (x"86",x"c8",x"0f",x"00"),
   989 => (x"9a",x"72",x"4a",x"70"),
   990 => (x"87",x"df",x"c1",x"02"),
   991 => (x"00",x"1c",x"fc",x"27"),
   992 => (x"c7",x"4a",x"bf",x"00"),
   993 => (x"2a",x"c9",x"82",x"ff"),
   994 => (x"4b",x"c0",x"4d",x"72"),
   995 => (x"00",x"0f",x"fd",x"27"),
   996 => (x"25",x"27",x"1e",x"00"),
   997 => (x"0f",x"00",x"00",x"18"),
   998 => (x"b7",x"c0",x"86",x"c4"),
   999 => (x"d0",x"c1",x"06",x"ad"),
  1000 => (x"27",x"1e",x"74",x"87"),
  1001 => (x"00",x"00",x"1c",x"f8"),
  1002 => (x"0f",x"06",x"27",x"1e"),
  1003 => (x"c8",x"0f",x"00",x"00"),
  1004 => (x"72",x"4a",x"70",x"86"),
  1005 => (x"c5",x"c0",x"05",x"9a"),
  1006 => (x"c0",x"48",x"c0",x"87"),
  1007 => (x"f8",x"27",x"87",x"f5"),
  1008 => (x"1e",x"00",x"00",x"1c"),
  1009 => (x"00",x"0e",x"cc",x"27"),
  1010 => (x"86",x"c4",x"0f",x"00"),
  1011 => (x"c1",x"84",x"c0",x"c8"),
  1012 => (x"ab",x"b7",x"75",x"83"),
  1013 => (x"87",x"c9",x"ff",x"04"),
  1014 => (x"d4",x"87",x"d6",x"c0"),
  1015 => (x"16",x"27",x"1e",x"66"),
  1016 => (x"1e",x"00",x"00",x"10"),
  1017 => (x"00",x"00",x"42",x"27"),
  1018 => (x"86",x"c8",x"0f",x"00"),
  1019 => (x"c2",x"c0",x"48",x"c0"),
  1020 => (x"26",x"48",x"c1",x"87"),
  1021 => (x"26",x"4c",x"26",x"4d"),
  1022 => (x"26",x"4a",x"26",x"4b"),
  1023 => (x"65",x"70",x"4f",x"4f"),
  1024 => (x"20",x"64",x"65",x"6e"),
  1025 => (x"65",x"6c",x"69",x"66"),
  1026 => (x"6f",x"6c",x"20",x"2c"),
  1027 => (x"6e",x"69",x"64",x"61"),
  1028 => (x"2e",x"2e",x"2e",x"67"),
  1029 => (x"61",x"43",x"00",x"0a"),
  1030 => (x"20",x"74",x"27",x"6e"),
  1031 => (x"6e",x"65",x"70",x"6f"),
  1032 => (x"0a",x"73",x"25",x"20"),
  1033 => (x"1e",x"72",x"1e",x"00"),
  1034 => (x"c0",x"02",x"66",x"c8"),
  1035 => (x"04",x"27",x"87",x"d1"),
  1036 => (x"49",x"00",x"00",x"1d"),
  1037 => (x"27",x"79",x"66",x"c8"),
  1038 => (x"00",x"00",x"1d",x"0c"),
  1039 => (x"27",x"79",x"c0",x"49"),
  1040 => (x"00",x"00",x"1d",x"0c"),
  1041 => (x"dc",x"c0",x"05",x"bf"),
  1042 => (x"1d",x"04",x"27",x"87"),
  1043 => (x"4a",x"bf",x"00",x"00"),
  1044 => (x"80",x"c4",x"48",x"72"),
  1045 => (x"00",x"1d",x"08",x"27"),
  1046 => (x"08",x"27",x"58",x"00"),
  1047 => (x"49",x"00",x"00",x"1d"),
  1048 => (x"cf",x"c0",x"79",x"6a"),
  1049 => (x"1d",x"08",x"27",x"87"),
  1050 => (x"48",x"bf",x"00",x"00"),
  1051 => (x"0c",x"27",x"30",x"c8"),
  1052 => (x"58",x"00",x"00",x"1d"),
  1053 => (x"00",x"1d",x"0c",x"27"),
  1054 => (x"c1",x"4a",x"bf",x"00"),
  1055 => (x"c3",x"48",x"72",x"82"),
  1056 => (x"1d",x"10",x"27",x"98"),
  1057 => (x"27",x"58",x"00",x"00"),
  1058 => (x"00",x"00",x"1d",x"08"),
  1059 => (x"b7",x"d8",x"4a",x"bf"),
  1060 => (x"26",x"48",x"72",x"2a"),
  1061 => (x"0e",x"4f",x"26",x"4a"),
  1062 => (x"0e",x"5b",x"5a",x"5e"),
  1063 => (x"fe",x"1e",x"66",x"cc"),
  1064 => (x"86",x"c4",x"87",x"c3"),
  1065 => (x"4a",x"c0",x"4b",x"70"),
  1066 => (x"c0",x"02",x"9b",x"73"),
  1067 => (x"82",x"c1",x"87",x"ce"),
  1068 => (x"f0",x"fd",x"1e",x"c0"),
  1069 => (x"70",x"86",x"c4",x"87"),
  1070 => (x"87",x"ec",x"ff",x"4b"),
  1071 => (x"4b",x"26",x"48",x"72"),
  1072 => (x"4f",x"26",x"4a",x"26"),
  1073 => (x"5b",x"5a",x"5e",x"0e"),
  1074 => (x"c8",x"0e",x"5d",x"5c"),
  1075 => (x"e4",x"f6",x"c0",x"8e"),
  1076 => (x"c0",x"4c",x"c4",x"c0"),
  1077 => (x"c0",x"c0",x"e4",x"f6"),
  1078 => (x"1e",x"66",x"dc",x"4b"),
  1079 => (x"c4",x"87",x"f8",x"fe"),
  1080 => (x"72",x"4a",x"70",x"86"),
  1081 => (x"76",x"85",x"c2",x"4d"),
  1082 => (x"d0",x"79",x"c1",x"49"),
  1083 => (x"c0",x"c1",x"7c",x"9f"),
  1084 => (x"9f",x"7b",x"9f",x"c1"),
  1085 => (x"ff",x"cf",x"4a",x"6b"),
  1086 => (x"9f",x"c0",x"9a",x"ff"),
  1087 => (x"7b",x"9f",x"c0",x"7b"),
  1088 => (x"cf",x"48",x"6b",x"9f"),
  1089 => (x"c8",x"98",x"ff",x"ff"),
  1090 => (x"c0",x"c4",x"58",x"a6"),
  1091 => (x"02",x"9a",x"72",x"9a"),
  1092 => (x"6e",x"87",x"fd",x"c1"),
  1093 => (x"87",x"e6",x"c0",x"02"),
  1094 => (x"c8",x"49",x"66",x"c4"),
  1095 => (x"05",x"a9",x"c6",x"c0"),
  1096 => (x"76",x"87",x"ed",x"c1"),
  1097 => (x"fa",x"79",x"c0",x"49"),
  1098 => (x"7b",x"9f",x"ca",x"eb"),
  1099 => (x"c0",x"7b",x"9f",x"c1"),
  1100 => (x"9f",x"75",x"7b",x"9f"),
  1101 => (x"7b",x"9f",x"c0",x"7b"),
  1102 => (x"c1",x"7b",x"9f",x"c0"),
  1103 => (x"4a",x"75",x"87",x"d2"),
  1104 => (x"c0",x"c8",x"2a",x"c1"),
  1105 => (x"66",x"c4",x"b2",x"c0"),
  1106 => (x"05",x"a9",x"72",x"49"),
  1107 => (x"dc",x"87",x"c1",x"c1"),
  1108 => (x"d0",x"fb",x"1e",x"66"),
  1109 => (x"c4",x"86",x"c4",x"87"),
  1110 => (x"4a",x"75",x"58",x"a6"),
  1111 => (x"9a",x"72",x"8d",x"c1"),
  1112 => (x"87",x"de",x"c0",x"02"),
  1113 => (x"97",x"74",x"4c",x"6e"),
  1114 => (x"02",x"9c",x"74",x"7b"),
  1115 => (x"c0",x"87",x"c9",x"c0"),
  1116 => (x"87",x"f1",x"fa",x"1e"),
  1117 => (x"4c",x"70",x"86",x"c4"),
  1118 => (x"8d",x"c1",x"4a",x"75"),
  1119 => (x"ff",x"05",x"9a",x"72"),
  1120 => (x"f6",x"c0",x"87",x"e4"),
  1121 => (x"4c",x"c4",x"c0",x"e4"),
  1122 => (x"c1",x"7c",x"9f",x"d1"),
  1123 => (x"87",x"c6",x"c0",x"48"),
  1124 => (x"fd",x"7c",x"9f",x"d1"),
  1125 => (x"86",x"c8",x"87",x"d5"),
  1126 => (x"4c",x"26",x"4d",x"26"),
  1127 => (x"4a",x"26",x"4b",x"26"),
  1128 => (x"5e",x"0e",x"4f",x"26"),
  1129 => (x"0e",x"5c",x"5b",x"5a"),
  1130 => (x"c3",x"8e",x"e4",x"c0"),
  1131 => (x"f6",x"c0",x"4c",x"ff"),
  1132 => (x"4b",x"c0",x"c0",x"e4"),
  1133 => (x"4a",x"6b",x"7b",x"74"),
  1134 => (x"7b",x"74",x"9a",x"74"),
  1135 => (x"98",x"74",x"48",x"6b"),
  1136 => (x"6e",x"58",x"a6",x"c4"),
  1137 => (x"c8",x"30",x"c8",x"48"),
  1138 => (x"a6",x"c8",x"58",x"a6"),
  1139 => (x"72",x"79",x"72",x"49"),
  1140 => (x"b2",x"66",x"c4",x"4a"),
  1141 => (x"48",x"6b",x"7b",x"74"),
  1142 => (x"a6",x"d0",x"98",x"74"),
  1143 => (x"48",x"66",x"cc",x"58"),
  1144 => (x"a6",x"d4",x"30",x"d0"),
  1145 => (x"49",x"a6",x"d4",x"58"),
  1146 => (x"4a",x"72",x"79",x"72"),
  1147 => (x"74",x"b2",x"66",x"d0"),
  1148 => (x"74",x"48",x"6b",x"7b"),
  1149 => (x"58",x"a6",x"dc",x"98"),
  1150 => (x"d8",x"48",x"66",x"d8"),
  1151 => (x"a6",x"e0",x"c0",x"30"),
  1152 => (x"a6",x"e0",x"c0",x"58"),
  1153 => (x"72",x"79",x"72",x"49"),
  1154 => (x"b2",x"66",x"dc",x"4a"),
  1155 => (x"e4",x"c0",x"48",x"72"),
  1156 => (x"26",x"4c",x"26",x"86"),
  1157 => (x"26",x"4a",x"26",x"4b"),
  1158 => (x"5a",x"5e",x"0e",x"4f"),
  1159 => (x"d8",x"0e",x"5c",x"5b"),
  1160 => (x"4c",x"ff",x"c3",x"8e"),
  1161 => (x"c0",x"e4",x"f6",x"c0"),
  1162 => (x"7b",x"74",x"4b",x"c0"),
  1163 => (x"9a",x"74",x"4a",x"6b"),
  1164 => (x"32",x"c8",x"7b",x"74"),
  1165 => (x"98",x"74",x"48",x"6b"),
  1166 => (x"c4",x"58",x"a6",x"c4"),
  1167 => (x"79",x"72",x"49",x"a6"),
  1168 => (x"b2",x"6e",x"4a",x"72"),
  1169 => (x"32",x"c8",x"7b",x"74"),
  1170 => (x"98",x"74",x"48",x"6b"),
  1171 => (x"cc",x"58",x"a6",x"cc"),
  1172 => (x"79",x"72",x"49",x"a6"),
  1173 => (x"66",x"c8",x"4a",x"72"),
  1174 => (x"c8",x"7b",x"74",x"b2"),
  1175 => (x"74",x"48",x"6b",x"32"),
  1176 => (x"58",x"a6",x"d4",x"98"),
  1177 => (x"72",x"49",x"a6",x"d4"),
  1178 => (x"d0",x"4a",x"72",x"79"),
  1179 => (x"48",x"72",x"b2",x"66"),
  1180 => (x"4c",x"26",x"86",x"d8"),
  1181 => (x"4a",x"26",x"4b",x"26"),
  1182 => (x"5e",x"0e",x"4f",x"26"),
  1183 => (x"5d",x"5c",x"5b",x"5a"),
  1184 => (x"e4",x"f6",x"c0",x"0e"),
  1185 => (x"d4",x"4b",x"c0",x"c0"),
  1186 => (x"ff",x"c3",x"48",x"66"),
  1187 => (x"27",x"7b",x"70",x"98"),
  1188 => (x"00",x"00",x"1d",x"10"),
  1189 => (x"c8",x"c0",x"05",x"bf"),
  1190 => (x"48",x"66",x"d8",x"87"),
  1191 => (x"a6",x"dc",x"30",x"c9"),
  1192 => (x"4a",x"66",x"d8",x"58"),
  1193 => (x"48",x"72",x"2a",x"d8"),
  1194 => (x"70",x"98",x"ff",x"c3"),
  1195 => (x"4a",x"66",x"d8",x"7b"),
  1196 => (x"48",x"72",x"2a",x"d0"),
  1197 => (x"70",x"98",x"ff",x"c3"),
  1198 => (x"4a",x"66",x"d8",x"7b"),
  1199 => (x"48",x"72",x"2a",x"c8"),
  1200 => (x"70",x"98",x"ff",x"c3"),
  1201 => (x"48",x"66",x"d8",x"7b"),
  1202 => (x"70",x"98",x"ff",x"c3"),
  1203 => (x"4a",x"66",x"d4",x"7b"),
  1204 => (x"48",x"72",x"2a",x"d0"),
  1205 => (x"70",x"98",x"ff",x"c3"),
  1206 => (x"c3",x"4d",x"6b",x"7b"),
  1207 => (x"f0",x"c9",x"9d",x"ff"),
  1208 => (x"ff",x"c3",x"4c",x"ff"),
  1209 => (x"c0",x"05",x"ad",x"b7"),
  1210 => (x"ff",x"c3",x"87",x"d8"),
  1211 => (x"6b",x"7b",x"72",x"4a"),
  1212 => (x"c1",x"9d",x"72",x"4d"),
  1213 => (x"02",x"9c",x"74",x"8c"),
  1214 => (x"72",x"87",x"c7",x"c0"),
  1215 => (x"ff",x"02",x"ad",x"b7"),
  1216 => (x"1e",x"75",x"87",x"eb"),
  1217 => (x"00",x"1a",x"6f",x"27"),
  1218 => (x"42",x"27",x"1e",x"00"),
  1219 => (x"0f",x"00",x"00",x"00"),
  1220 => (x"48",x"75",x"86",x"c8"),
  1221 => (x"4c",x"26",x"4d",x"26"),
  1222 => (x"4a",x"26",x"4b",x"26"),
  1223 => (x"5e",x"0e",x"4f",x"26"),
  1224 => (x"c0",x"0e",x"5b",x"5a"),
  1225 => (x"c0",x"c0",x"e4",x"f6"),
  1226 => (x"c3",x"4a",x"c0",x"4b"),
  1227 => (x"82",x"c1",x"7b",x"ff"),
  1228 => (x"aa",x"b7",x"c8",x"c3"),
  1229 => (x"87",x"f3",x"ff",x"04"),
  1230 => (x"4a",x"26",x"4b",x"26"),
  1231 => (x"5e",x"0e",x"4f",x"26"),
  1232 => (x"5d",x"5c",x"5b",x"5a"),
  1233 => (x"c0",x"c0",x"c1",x"0e"),
  1234 => (x"4c",x"c0",x"c0",x"c0"),
  1235 => (x"c0",x"e4",x"f6",x"c0"),
  1236 => (x"1e",x"27",x"4b",x"c0"),
  1237 => (x"0f",x"00",x"00",x"13"),
  1238 => (x"4d",x"df",x"f8",x"c4"),
  1239 => (x"ff",x"c0",x"1e",x"c0"),
  1240 => (x"1e",x"f7",x"c1",x"f0"),
  1241 => (x"00",x"12",x"7a",x"27"),
  1242 => (x"86",x"c8",x"0f",x"00"),
  1243 => (x"b7",x"c1",x"4a",x"70"),
  1244 => (x"dc",x"c1",x"05",x"aa"),
  1245 => (x"27",x"1e",x"72",x"87"),
  1246 => (x"00",x"00",x"13",x"ff"),
  1247 => (x"00",x"42",x"27",x"1e"),
  1248 => (x"c8",x"0f",x"00",x"00"),
  1249 => (x"7b",x"ff",x"c3",x"86"),
  1250 => (x"e1",x"c0",x"1e",x"74"),
  1251 => (x"1e",x"e9",x"c1",x"f0"),
  1252 => (x"00",x"12",x"7a",x"27"),
  1253 => (x"86",x"c8",x"0f",x"00"),
  1254 => (x"9a",x"72",x"4a",x"70"),
  1255 => (x"87",x"d8",x"c0",x"05"),
  1256 => (x"f5",x"27",x"1e",x"72"),
  1257 => (x"1e",x"00",x"00",x"13"),
  1258 => (x"00",x"00",x"42",x"27"),
  1259 => (x"86",x"c8",x"0f",x"00"),
  1260 => (x"c1",x"7b",x"ff",x"c3"),
  1261 => (x"87",x"f3",x"c0",x"48"),
  1262 => (x"09",x"27",x"1e",x"72"),
  1263 => (x"1e",x"00",x"00",x"14"),
  1264 => (x"00",x"00",x"42",x"27"),
  1265 => (x"86",x"c8",x"0f",x"00"),
  1266 => (x"00",x"13",x"1e",x"27"),
  1267 => (x"d0",x"c0",x"0f",x"00"),
  1268 => (x"27",x"1e",x"72",x"87"),
  1269 => (x"00",x"00",x"14",x"13"),
  1270 => (x"00",x"42",x"27",x"1e"),
  1271 => (x"c8",x"0f",x"00",x"00"),
  1272 => (x"75",x"8d",x"c1",x"86"),
  1273 => (x"f3",x"fd",x"05",x"9d"),
  1274 => (x"26",x"48",x"c0",x"87"),
  1275 => (x"26",x"4c",x"26",x"4d"),
  1276 => (x"26",x"4a",x"26",x"4b"),
  1277 => (x"44",x"4d",x"43",x"4f"),
  1278 => (x"25",x"20",x"31",x"34"),
  1279 => (x"43",x"00",x"0a",x"64"),
  1280 => (x"35",x"35",x"44",x"4d"),
  1281 => (x"0a",x"64",x"25",x"20"),
  1282 => (x"44",x"4d",x"43",x"00"),
  1283 => (x"25",x"20",x"31",x"34"),
  1284 => (x"43",x"00",x"0a",x"64"),
  1285 => (x"35",x"35",x"44",x"4d"),
  1286 => (x"0a",x"64",x"25",x"20"),
  1287 => (x"5a",x"5e",x"0e",x"00"),
  1288 => (x"0e",x"5d",x"5c",x"5b"),
  1289 => (x"c1",x"f0",x"ff",x"c0"),
  1290 => (x"f6",x"c0",x"4d",x"c1"),
  1291 => (x"4b",x"c0",x"c0",x"e4"),
  1292 => (x"27",x"7b",x"ff",x"c3"),
  1293 => (x"00",x"00",x"14",x"af"),
  1294 => (x"18",x"25",x"27",x"1e"),
  1295 => (x"c4",x"0f",x"00",x"00"),
  1296 => (x"c0",x"4c",x"d3",x"86"),
  1297 => (x"27",x"1e",x"75",x"1e"),
  1298 => (x"00",x"00",x"12",x"7a"),
  1299 => (x"70",x"86",x"c8",x"0f"),
  1300 => (x"05",x"9a",x"72",x"4a"),
  1301 => (x"72",x"87",x"d8",x"c0"),
  1302 => (x"14",x"99",x"27",x"1e"),
  1303 => (x"27",x"1e",x"00",x"00"),
  1304 => (x"00",x"00",x"00",x"42"),
  1305 => (x"c3",x"86",x"c8",x"0f"),
  1306 => (x"48",x"c1",x"7b",x"ff"),
  1307 => (x"72",x"87",x"e0",x"c0"),
  1308 => (x"14",x"a4",x"27",x"1e"),
  1309 => (x"27",x"1e",x"00",x"00"),
  1310 => (x"00",x"00",x"00",x"42"),
  1311 => (x"27",x"86",x"c8",x"0f"),
  1312 => (x"00",x"00",x"13",x"1e"),
  1313 => (x"74",x"8c",x"c1",x"0f"),
  1314 => (x"f6",x"fe",x"05",x"9c"),
  1315 => (x"26",x"48",x"c0",x"87"),
  1316 => (x"26",x"4c",x"26",x"4d"),
  1317 => (x"26",x"4a",x"26",x"4b"),
  1318 => (x"69",x"6e",x"69",x"4f"),
  1319 => (x"64",x"25",x"20",x"74"),
  1320 => (x"00",x"20",x"20",x"0a"),
  1321 => (x"74",x"69",x"6e",x"69"),
  1322 => (x"0a",x"64",x"25",x"20"),
  1323 => (x"43",x"00",x"20",x"20"),
  1324 => (x"69",x"5f",x"64",x"6d"),
  1325 => (x"0a",x"74",x"69",x"6e"),
  1326 => (x"5a",x"5e",x"0e",x"00"),
  1327 => (x"0e",x"5d",x"5c",x"5b"),
  1328 => (x"4d",x"ff",x"c3",x"1e"),
  1329 => (x"c0",x"e4",x"f6",x"c0"),
  1330 => (x"1e",x"27",x"4b",x"c0"),
  1331 => (x"0f",x"00",x"00",x"13"),
  1332 => (x"c0",x"1e",x"ea",x"c6"),
  1333 => (x"c8",x"c1",x"f0",x"e1"),
  1334 => (x"12",x"7a",x"27",x"1e"),
  1335 => (x"c8",x"0f",x"00",x"00"),
  1336 => (x"72",x"4a",x"70",x"86"),
  1337 => (x"16",x"42",x"27",x"1e"),
  1338 => (x"27",x"1e",x"00",x"00"),
  1339 => (x"00",x"00",x"00",x"42"),
  1340 => (x"c1",x"86",x"c8",x"0f"),
  1341 => (x"c0",x"02",x"aa",x"b7"),
  1342 => (x"1d",x"27",x"87",x"cb"),
  1343 => (x"0f",x"00",x"00",x"14"),
  1344 => (x"db",x"c3",x"48",x"c0"),
  1345 => (x"12",x"19",x"27",x"87"),
  1346 => (x"70",x"0f",x"00",x"00"),
  1347 => (x"cf",x"4a",x"74",x"4c"),
  1348 => (x"c6",x"9a",x"ff",x"ff"),
  1349 => (x"02",x"aa",x"b7",x"ea"),
  1350 => (x"74",x"87",x"db",x"c0"),
  1351 => (x"15",x"eb",x"27",x"1e"),
  1352 => (x"27",x"1e",x"00",x"00"),
  1353 => (x"00",x"00",x"00",x"42"),
  1354 => (x"27",x"86",x"c8",x"0f"),
  1355 => (x"00",x"00",x"14",x"1d"),
  1356 => (x"c2",x"48",x"c0",x"0f"),
  1357 => (x"7b",x"75",x"87",x"ea"),
  1358 => (x"f1",x"c0",x"49",x"76"),
  1359 => (x"13",x"3e",x"27",x"79"),
  1360 => (x"70",x"0f",x"00",x"00"),
  1361 => (x"02",x"9a",x"72",x"4a"),
  1362 => (x"c0",x"87",x"eb",x"c1"),
  1363 => (x"f0",x"ff",x"c0",x"1e"),
  1364 => (x"27",x"1e",x"fa",x"c1"),
  1365 => (x"00",x"00",x"12",x"7a"),
  1366 => (x"70",x"86",x"c8",x"0f"),
  1367 => (x"05",x"9c",x"74",x"4c"),
  1368 => (x"74",x"87",x"c3",x"c1"),
  1369 => (x"16",x"00",x"27",x"1e"),
  1370 => (x"27",x"1e",x"00",x"00"),
  1371 => (x"00",x"00",x"00",x"42"),
  1372 => (x"75",x"86",x"c8",x"0f"),
  1373 => (x"75",x"4c",x"6b",x"7b"),
  1374 => (x"27",x"1e",x"74",x"9c"),
  1375 => (x"00",x"00",x"16",x"0c"),
  1376 => (x"00",x"42",x"27",x"1e"),
  1377 => (x"c8",x"0f",x"00",x"00"),
  1378 => (x"75",x"7b",x"75",x"86"),
  1379 => (x"75",x"7b",x"75",x"7b"),
  1380 => (x"c1",x"4a",x"74",x"7b"),
  1381 => (x"9a",x"72",x"9a",x"c0"),
  1382 => (x"87",x"c5",x"c0",x"02"),
  1383 => (x"ff",x"c0",x"48",x"c1"),
  1384 => (x"c0",x"48",x"c0",x"87"),
  1385 => (x"1e",x"74",x"87",x"fa"),
  1386 => (x"00",x"16",x"1a",x"27"),
  1387 => (x"42",x"27",x"1e",x"00"),
  1388 => (x"0f",x"00",x"00",x"00"),
  1389 => (x"49",x"6e",x"86",x"c8"),
  1390 => (x"05",x"a9",x"b7",x"c2"),
  1391 => (x"27",x"87",x"d3",x"c0"),
  1392 => (x"00",x"00",x"16",x"26"),
  1393 => (x"00",x"42",x"27",x"1e"),
  1394 => (x"c4",x"0f",x"00",x"00"),
  1395 => (x"c0",x"48",x"c0",x"86"),
  1396 => (x"48",x"6e",x"87",x"ce"),
  1397 => (x"a6",x"c4",x"88",x"c1"),
  1398 => (x"fd",x"05",x"6e",x"58"),
  1399 => (x"48",x"c0",x"87",x"df"),
  1400 => (x"26",x"4d",x"26",x"26"),
  1401 => (x"26",x"4b",x"26",x"4c"),
  1402 => (x"43",x"4f",x"26",x"4a"),
  1403 => (x"5f",x"38",x"44",x"4d"),
  1404 => (x"65",x"72",x"20",x"34"),
  1405 => (x"6e",x"6f",x"70",x"73"),
  1406 => (x"20",x"3a",x"65",x"73"),
  1407 => (x"00",x"0a",x"64",x"25"),
  1408 => (x"35",x"44",x"4d",x"43"),
  1409 => (x"64",x"25",x"20",x"38"),
  1410 => (x"00",x"20",x"20",x"0a"),
  1411 => (x"35",x"44",x"4d",x"43"),
  1412 => (x"20",x"32",x"5f",x"38"),
  1413 => (x"20",x"0a",x"64",x"25"),
  1414 => (x"4d",x"43",x"00",x"20"),
  1415 => (x"20",x"38",x"35",x"44"),
  1416 => (x"20",x"0a",x"64",x"25"),
  1417 => (x"44",x"53",x"00",x"20"),
  1418 => (x"49",x"20",x"43",x"48"),
  1419 => (x"69",x"74",x"69",x"6e"),
  1420 => (x"7a",x"69",x"6c",x"61"),
  1421 => (x"6f",x"69",x"74",x"61"),
  1422 => (x"72",x"65",x"20",x"6e"),
  1423 => (x"21",x"72",x"6f",x"72"),
  1424 => (x"6d",x"63",x"00",x"0a"),
  1425 => (x"4d",x"43",x"5f",x"64"),
  1426 => (x"72",x"20",x"38",x"44"),
  1427 => (x"6f",x"70",x"73",x"65"),
  1428 => (x"3a",x"65",x"73",x"6e"),
  1429 => (x"0a",x"64",x"25",x"20"),
  1430 => (x"5a",x"5e",x"0e",x"00"),
  1431 => (x"0e",x"5d",x"5c",x"5b"),
  1432 => (x"c0",x"e4",x"f6",x"c0"),
  1433 => (x"f6",x"c0",x"4d",x"c0"),
  1434 => (x"4b",x"c4",x"c0",x"e4"),
  1435 => (x"00",x"1d",x"10",x"27"),
  1436 => (x"79",x"c1",x"49",x"00"),
  1437 => (x"c0",x"e4",x"f6",x"c0"),
  1438 => (x"e0",x"c0",x"49",x"c8"),
  1439 => (x"c3",x"4c",x"c7",x"79"),
  1440 => (x"13",x"1e",x"27",x"7b"),
  1441 => (x"c2",x"0f",x"00",x"00"),
  1442 => (x"7d",x"ff",x"c3",x"7b"),
  1443 => (x"e5",x"c0",x"1e",x"c0"),
  1444 => (x"1e",x"c0",x"c1",x"d0"),
  1445 => (x"00",x"12",x"7a",x"27"),
  1446 => (x"86",x"c8",x"0f",x"00"),
  1447 => (x"b7",x"c1",x"4a",x"70"),
  1448 => (x"c2",x"c0",x"05",x"aa"),
  1449 => (x"c2",x"4c",x"c1",x"87"),
  1450 => (x"c0",x"05",x"ac",x"b7"),
  1451 => (x"48",x"c0",x"87",x"c5"),
  1452 => (x"c1",x"87",x"f8",x"c0"),
  1453 => (x"05",x"9c",x"74",x"8c"),
  1454 => (x"27",x"87",x"c4",x"ff"),
  1455 => (x"00",x"00",x"14",x"b9"),
  1456 => (x"1d",x"14",x"27",x"0f"),
  1457 => (x"27",x"58",x"00",x"00"),
  1458 => (x"00",x"00",x"1d",x"10"),
  1459 => (x"d0",x"c0",x"05",x"bf"),
  1460 => (x"c0",x"1e",x"c1",x"87"),
  1461 => (x"d0",x"c1",x"f0",x"ff"),
  1462 => (x"12",x"7a",x"27",x"1e"),
  1463 => (x"c8",x"0f",x"00",x"00"),
  1464 => (x"7d",x"ff",x"c3",x"86"),
  1465 => (x"ff",x"c3",x"7b",x"c3"),
  1466 => (x"26",x"48",x"c1",x"7d"),
  1467 => (x"26",x"4c",x"26",x"4d"),
  1468 => (x"26",x"4a",x"26",x"4b"),
  1469 => (x"48",x"c0",x"1e",x"4f"),
  1470 => (x"5e",x"0e",x"4f",x"26"),
  1471 => (x"5d",x"5c",x"5b",x"5a"),
  1472 => (x"c0",x"8e",x"c8",x"0e"),
  1473 => (x"c0",x"4d",x"66",x"e0"),
  1474 => (x"c0",x"c0",x"e4",x"f6"),
  1475 => (x"c0",x"49",x"76",x"4b"),
  1476 => (x"c0",x"1e",x"75",x"79"),
  1477 => (x"27",x"1e",x"66",x"e0"),
  1478 => (x"00",x"00",x"17",x"df"),
  1479 => (x"00",x"42",x"27",x"1e"),
  1480 => (x"cc",x"0f",x"00",x"00"),
  1481 => (x"7b",x"ff",x"c3",x"86"),
  1482 => (x"c0",x"e4",x"f6",x"c0"),
  1483 => (x"79",x"c2",x"49",x"c4"),
  1484 => (x"c0",x"e4",x"f6",x"c0"),
  1485 => (x"79",x"c1",x"49",x"c8"),
  1486 => (x"dc",x"7b",x"ff",x"c3"),
  1487 => (x"ff",x"c0",x"1e",x"66"),
  1488 => (x"1e",x"d1",x"c1",x"f0"),
  1489 => (x"00",x"12",x"7a",x"27"),
  1490 => (x"86",x"c8",x"0f",x"00"),
  1491 => (x"c4",x"58",x"a6",x"c8"),
  1492 => (x"d8",x"c0",x"02",x"66"),
  1493 => (x"1e",x"66",x"c4",x"87"),
  1494 => (x"1e",x"66",x"e0",x"c0"),
  1495 => (x"00",x"17",x"bf",x"27"),
  1496 => (x"42",x"27",x"1e",x"00"),
  1497 => (x"0f",x"00",x"00",x"00"),
  1498 => (x"c4",x"c1",x"86",x"cc"),
  1499 => (x"cd",x"ee",x"c5",x"87"),
  1500 => (x"ff",x"c3",x"4c",x"df"),
  1501 => (x"c3",x"4a",x"6b",x"7b"),
  1502 => (x"fe",x"c3",x"9a",x"ff"),
  1503 => (x"c0",x"05",x"aa",x"b7"),
  1504 => (x"4a",x"c0",x"87",x"dc"),
  1505 => (x"00",x"11",x"a2",x"27"),
  1506 => (x"7d",x"70",x"0f",x"00"),
  1507 => (x"82",x"c1",x"85",x"c4"),
  1508 => (x"aa",x"b7",x"c0",x"c2"),
  1509 => (x"87",x"ec",x"ff",x"04"),
  1510 => (x"49",x"76",x"4c",x"c1"),
  1511 => (x"8c",x"c1",x"79",x"c1"),
  1512 => (x"ff",x"05",x"9c",x"74"),
  1513 => (x"ff",x"c3",x"87",x"cc"),
  1514 => (x"e4",x"f6",x"c0",x"7b"),
  1515 => (x"c3",x"49",x"c4",x"c0"),
  1516 => (x"c8",x"48",x"6e",x"79"),
  1517 => (x"26",x"4d",x"26",x"86"),
  1518 => (x"26",x"4b",x"26",x"4c"),
  1519 => (x"52",x"4f",x"26",x"4a"),
  1520 => (x"20",x"64",x"61",x"65"),
  1521 => (x"6d",x"6d",x"6f",x"63"),
  1522 => (x"20",x"64",x"6e",x"61"),
  1523 => (x"6c",x"69",x"61",x"66"),
  1524 => (x"61",x"20",x"64",x"65"),
  1525 => (x"64",x"25",x"20",x"74"),
  1526 => (x"64",x"25",x"28",x"20"),
  1527 => (x"73",x"00",x"0a",x"29"),
  1528 => (x"65",x"72",x"5f",x"64"),
  1529 => (x"73",x"5f",x"64",x"61"),
  1530 => (x"6f",x"74",x"63",x"65"),
  1531 => (x"64",x"25",x"20",x"72"),
  1532 => (x"64",x"25",x"20",x"2c"),
  1533 => (x"72",x"1e",x"00",x"0a"),
  1534 => (x"f6",x"c0",x"1e",x"1e"),
  1535 => (x"4a",x"c0",x"c0",x"e8"),
  1536 => (x"c0",x"c4",x"48",x"6a"),
  1537 => (x"58",x"a6",x"c4",x"98"),
  1538 => (x"cd",x"c0",x"05",x"6e"),
  1539 => (x"c4",x"48",x"6a",x"87"),
  1540 => (x"a6",x"c4",x"98",x"c0"),
  1541 => (x"ff",x"02",x"6e",x"58"),
  1542 => (x"66",x"cc",x"87",x"f3"),
  1543 => (x"48",x"66",x"cc",x"7a"),
  1544 => (x"26",x"4a",x"26",x"26"),
  1545 => (x"5a",x"5e",x"0e",x"4f"),
  1546 => (x"d0",x"0e",x"5c",x"5b"),
  1547 => (x"4c",x"c0",x"4b",x"66"),
  1548 => (x"c0",x"c1",x"4a",x"13"),
  1549 => (x"92",x"c0",x"c0",x"c0"),
  1550 => (x"92",x"b7",x"c0",x"c4"),
  1551 => (x"27",x"1e",x"72",x"4a"),
  1552 => (x"00",x"00",x"17",x"f6"),
  1553 => (x"c1",x"86",x"c4",x"0f"),
  1554 => (x"05",x"9a",x"72",x"84"),
  1555 => (x"74",x"87",x"e1",x"ff"),
  1556 => (x"26",x"4c",x"26",x"48"),
  1557 => (x"26",x"4a",x"26",x"4b"),
  1558 => (x"5a",x"5e",x"0e",x"4f"),
  1559 => (x"0e",x"5d",x"5c",x"5b"),
  1560 => (x"e0",x"c0",x"8e",x"c8"),
  1561 => (x"66",x"dc",x"4c",x"66"),
  1562 => (x"c0",x"49",x"76",x"4a"),
  1563 => (x"ac",x"b7",x"c0",x"79"),
  1564 => (x"87",x"ee",x"c1",x"06"),
  1565 => (x"ff",x"c3",x"4b",x"12"),
  1566 => (x"c1",x"33",x"c8",x"9b"),
  1567 => (x"ac",x"b7",x"c0",x"8c"),
  1568 => (x"87",x"cb",x"c0",x"06"),
  1569 => (x"ff",x"c3",x"48",x"12"),
  1570 => (x"58",x"a6",x"c8",x"98"),
  1571 => (x"c4",x"87",x"c5",x"c0"),
  1572 => (x"79",x"c0",x"49",x"a6"),
  1573 => (x"66",x"c4",x"4b",x"73"),
  1574 => (x"c1",x"33",x"c8",x"b3"),
  1575 => (x"ac",x"b7",x"c0",x"8c"),
  1576 => (x"87",x"c8",x"c0",x"06"),
  1577 => (x"ff",x"c3",x"4d",x"12"),
  1578 => (x"87",x"c2",x"c0",x"9d"),
  1579 => (x"4b",x"73",x"4d",x"c0"),
  1580 => (x"33",x"c8",x"b3",x"75"),
  1581 => (x"b7",x"c0",x"8c",x"c1"),
  1582 => (x"cb",x"c0",x"06",x"ac"),
  1583 => (x"c3",x"48",x"12",x"87"),
  1584 => (x"a6",x"c8",x"98",x"ff"),
  1585 => (x"87",x"c5",x"c0",x"58"),
  1586 => (x"c0",x"49",x"a6",x"c4"),
  1587 => (x"c4",x"4b",x"73",x"79"),
  1588 => (x"48",x"73",x"b3",x"66"),
  1589 => (x"a6",x"c4",x"80",x"6e"),
  1590 => (x"c0",x"8c",x"c1",x"58"),
  1591 => (x"fe",x"01",x"ac",x"b7"),
  1592 => (x"48",x"6e",x"87",x"d2"),
  1593 => (x"4d",x"26",x"86",x"c8"),
  1594 => (x"4b",x"26",x"4c",x"26"),
  1595 => (x"4f",x"26",x"4a",x"26"),
  1596 => (x"63",x"65",x"68",x"43"),
  1597 => (x"6d",x"75",x"73",x"6b"),
  1598 => (x"20",x"6f",x"74",x"20"),
  1599 => (x"20",x"3a",x"64",x"25"),
  1600 => (x"00",x"0a",x"64",x"25"),
  1601 => (x"64",x"61",x"65",x"52"),
  1602 => (x"20",x"66",x"6f",x"20"),
  1603 => (x"20",x"52",x"42",x"4d"),
  1604 => (x"6c",x"69",x"61",x"66"),
  1605 => (x"00",x"0a",x"64",x"65"),
  1606 => (x"70",x"20",x"6f",x"4e"),
  1607 => (x"69",x"74",x"72",x"61"),
  1608 => (x"6e",x"6f",x"69",x"74"),
  1609 => (x"67",x"69",x"73",x"20"),
  1610 => (x"75",x"74",x"61",x"6e"),
  1611 => (x"66",x"20",x"65",x"72"),
  1612 => (x"64",x"6e",x"75",x"6f"),
  1613 => (x"42",x"4d",x"00",x"0a"),
  1614 => (x"7a",x"69",x"73",x"52"),
  1615 => (x"25",x"20",x"3a",x"65"),
  1616 => (x"70",x"20",x"2c",x"64"),
  1617 => (x"69",x"74",x"72",x"61"),
  1618 => (x"6e",x"6f",x"69",x"74"),
  1619 => (x"65",x"7a",x"69",x"73"),
  1620 => (x"64",x"25",x"20",x"3a"),
  1621 => (x"66",x"6f",x"20",x"2c"),
  1622 => (x"74",x"65",x"73",x"66"),
  1623 => (x"20",x"66",x"6f",x"20"),
  1624 => (x"3a",x"67",x"69",x"73"),
  1625 => (x"2c",x"64",x"25",x"20"),
  1626 => (x"67",x"69",x"73",x"20"),
  1627 => (x"25",x"78",x"30",x"20"),
  1628 => (x"52",x"00",x"0a",x"78"),
  1629 => (x"69",x"64",x"61",x"65"),
  1630 => (x"62",x"20",x"67",x"6e"),
  1631 => (x"20",x"74",x"6f",x"6f"),
  1632 => (x"74",x"63",x"65",x"73"),
  1633 => (x"25",x"20",x"72",x"6f"),
  1634 => (x"52",x"00",x"0a",x"64"),
  1635 => (x"20",x"64",x"61",x"65"),
  1636 => (x"74",x"6f",x"6f",x"62"),
  1637 => (x"63",x"65",x"73",x"20"),
  1638 => (x"20",x"72",x"6f",x"74"),
  1639 => (x"6d",x"6f",x"72",x"66"),
  1640 => (x"72",x"69",x"66",x"20"),
  1641 => (x"70",x"20",x"74",x"73"),
  1642 => (x"69",x"74",x"72",x"61"),
  1643 => (x"6e",x"6f",x"69",x"74"),
  1644 => (x"6e",x"55",x"00",x"0a"),
  1645 => (x"70",x"70",x"75",x"73"),
  1646 => (x"65",x"74",x"72",x"6f"),
  1647 => (x"61",x"70",x"20",x"64"),
  1648 => (x"74",x"69",x"74",x"72"),
  1649 => (x"20",x"6e",x"6f",x"69"),
  1650 => (x"65",x"70",x"79",x"74"),
  1651 => (x"46",x"00",x"0d",x"21"),
  1652 => (x"32",x"33",x"54",x"41"),
  1653 => (x"00",x"20",x"20",x"20"),
  1654 => (x"64",x"61",x"65",x"52"),
  1655 => (x"20",x"67",x"6e",x"69"),
  1656 => (x"0a",x"52",x"42",x"4d"),
  1657 => (x"52",x"42",x"4d",x"00"),
  1658 => (x"63",x"75",x"73",x"20"),
  1659 => (x"73",x"73",x"65",x"63"),
  1660 => (x"6c",x"6c",x"75",x"66"),
  1661 => (x"65",x"72",x"20",x"79"),
  1662 => (x"00",x"0a",x"64",x"61"),
  1663 => (x"31",x"54",x"41",x"46"),
  1664 => (x"20",x"20",x"20",x"36"),
  1665 => (x"54",x"41",x"46",x"00"),
  1666 => (x"20",x"20",x"32",x"33"),
  1667 => (x"61",x"50",x"00",x"20"),
  1668 => (x"74",x"69",x"74",x"72"),
  1669 => (x"63",x"6e",x"6f",x"69"),
  1670 => (x"74",x"6e",x"75",x"6f"),
  1671 => (x"0a",x"64",x"25",x"20"),
  1672 => (x"6e",x"75",x"48",x"00"),
  1673 => (x"67",x"6e",x"69",x"74"),
  1674 => (x"72",x"6f",x"66",x"20"),
  1675 => (x"6c",x"69",x"66",x"20"),
  1676 => (x"73",x"79",x"73",x"65"),
  1677 => (x"0a",x"6d",x"65",x"74"),
  1678 => (x"54",x"41",x"46",x"00"),
  1679 => (x"20",x"20",x"32",x"33"),
  1680 => (x"41",x"46",x"00",x"20"),
  1681 => (x"20",x"36",x"31",x"54"),
  1682 => (x"43",x"00",x"20",x"20"),
  1683 => (x"74",x"73",x"75",x"6c"),
  1684 => (x"73",x"20",x"72",x"65"),
  1685 => (x"3a",x"65",x"7a",x"69"),
  1686 => (x"2c",x"64",x"25",x"20"),
  1687 => (x"75",x"6c",x"43",x"20"),
  1688 => (x"72",x"65",x"74",x"73"),
  1689 => (x"73",x"61",x"6d",x"20"),
  1690 => (x"25",x"20",x"2c",x"6b"),
  1691 => (x"47",x"00",x"0a",x"64"),
  1692 => (x"72",x"20",x"74",x"6f"),
  1693 => (x"6c",x"75",x"73",x"65"),
  1694 => (x"64",x"25",x"20",x"74"),
  1695 => (x"64",x"00",x"0a",x"20"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
