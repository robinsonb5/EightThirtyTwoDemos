
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"3b",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"38"),
    10 => (x"20",x"00",x"27",x"4f"),
    11 => (x"27",x"4e",x"00",x"00"),
    12 => (x"00",x"00",x"13",x"c6"),
    13 => (x"87",x"fd",x"00",x"0f"),
    14 => (x"4f",x"87",x"fd",x"00"),
    15 => (x"c0",x"ff",x"1e",x"1e"),
    16 => (x"c4",x"48",x"69",x"49"),
    17 => (x"a6",x"c4",x"98",x"c0"),
    18 => (x"f4",x"02",x"6e",x"58"),
    19 => (x"79",x"66",x"c8",x"87"),
    20 => (x"87",x"c6",x"26",x"48"),
    21 => (x"4c",x"26",x"4d",x"26"),
    22 => (x"4f",x"26",x"4b",x"26"),
    23 => (x"5c",x"5b",x"5e",x"0e"),
    24 => (x"4c",x"66",x"cc",x"0e"),
    25 => (x"4a",x"14",x"4b",x"c0"),
    26 => (x"72",x"9a",x"ff",x"c3"),
    27 => (x"87",x"d5",x"02",x"9a"),
    28 => (x"1e",x"71",x"49",x"72"),
    29 => (x"c4",x"87",x"c5",x"ff"),
    30 => (x"14",x"83",x"c1",x"86"),
    31 => (x"9a",x"ff",x"c3",x"4a"),
    32 => (x"eb",x"05",x"9a",x"72"),
    33 => (x"ff",x"48",x"73",x"87"),
    34 => (x"5e",x"0e",x"87",x"cc"),
    35 => (x"0e",x"5d",x"5c",x"5b"),
    36 => (x"4b",x"c0",x"86",x"f0"),
    37 => (x"c0",x"48",x"a6",x"c4"),
    38 => (x"a6",x"e4",x"c0",x"78"),
    39 => (x"66",x"e0",x"c0",x"4c"),
    40 => (x"80",x"c1",x"48",x"49"),
    41 => (x"58",x"a6",x"e4",x"c0"),
    42 => (x"c0",x"fe",x"4a",x"11"),
    43 => (x"9a",x"72",x"ba",x"82"),
    44 => (x"87",x"d3",x"c4",x"02"),
    45 => (x"c3",x"02",x"66",x"c4"),
    46 => (x"a6",x"c4",x"87",x"e2"),
    47 => (x"72",x"78",x"c0",x"48"),
    48 => (x"aa",x"f0",x"c0",x"49"),
    49 => (x"87",x"f2",x"c2",x"02"),
    50 => (x"02",x"a9",x"e3",x"c1"),
    51 => (x"c1",x"87",x"f3",x"c2"),
    52 => (x"c0",x"02",x"a9",x"e4"),
    53 => (x"ec",x"c1",x"87",x"e1"),
    54 => (x"dd",x"c2",x"02",x"a9"),
    55 => (x"a9",x"f0",x"c1",x"87"),
    56 => (x"c1",x"87",x"d4",x"02"),
    57 => (x"c1",x"02",x"a9",x"f3"),
    58 => (x"f5",x"c1",x"87",x"fc"),
    59 => (x"87",x"c7",x"02",x"a9"),
    60 => (x"05",x"a9",x"f8",x"c1"),
    61 => (x"c4",x"87",x"dc",x"c2"),
    62 => (x"c4",x"49",x"74",x"84"),
    63 => (x"69",x"48",x"76",x"89"),
    64 => (x"c1",x"02",x"6e",x"78"),
    65 => (x"80",x"c8",x"87",x"d3"),
    66 => (x"a6",x"cc",x"78",x"c0"),
    67 => (x"6e",x"78",x"c0",x"48"),
    68 => (x"29",x"b7",x"dc",x"49"),
    69 => (x"9a",x"cf",x"4a",x"71"),
    70 => (x"30",x"c4",x"48",x"6e"),
    71 => (x"72",x"58",x"a6",x"c4"),
    72 => (x"87",x"c5",x"02",x"9a"),
    73 => (x"c1",x"48",x"a6",x"c8"),
    74 => (x"06",x"aa",x"c9",x"78"),
    75 => (x"f7",x"c0",x"87",x"c5"),
    76 => (x"c0",x"87",x"c3",x"82"),
    77 => (x"66",x"c8",x"82",x"f0"),
    78 => (x"72",x"87",x"c9",x"02"),
    79 => (x"87",x"fc",x"fb",x"1e"),
    80 => (x"83",x"c1",x"86",x"c4"),
    81 => (x"c1",x"48",x"66",x"cc"),
    82 => (x"58",x"a6",x"d0",x"80"),
    83 => (x"c8",x"48",x"66",x"cc"),
    84 => (x"fe",x"04",x"a8",x"b7"),
    85 => (x"d7",x"c1",x"87",x"f9"),
    86 => (x"1e",x"f0",x"c0",x"87"),
    87 => (x"c4",x"87",x"dd",x"fb"),
    88 => (x"c1",x"83",x"c1",x"86"),
    89 => (x"84",x"c4",x"87",x"ca"),
    90 => (x"89",x"c4",x"49",x"74"),
    91 => (x"eb",x"fb",x"1e",x"69"),
    92 => (x"70",x"86",x"c4",x"87"),
    93 => (x"c0",x"83",x"71",x"49"),
    94 => (x"a6",x"c4",x"87",x"f6"),
    95 => (x"c0",x"78",x"c1",x"48"),
    96 => (x"84",x"c4",x"87",x"ee"),
    97 => (x"89",x"c4",x"49",x"74"),
    98 => (x"ef",x"fa",x"1e",x"69"),
    99 => (x"c1",x"86",x"c4",x"87"),
   100 => (x"72",x"87",x"dd",x"83"),
   101 => (x"87",x"e4",x"fa",x"1e"),
   102 => (x"87",x"d4",x"86",x"c4"),
   103 => (x"05",x"aa",x"e5",x"c0"),
   104 => (x"a6",x"c4",x"87",x"c7"),
   105 => (x"c7",x"78",x"c1",x"48"),
   106 => (x"fa",x"1e",x"72",x"87"),
   107 => (x"86",x"c4",x"87",x"ce"),
   108 => (x"49",x"66",x"e0",x"c0"),
   109 => (x"c0",x"80",x"c1",x"48"),
   110 => (x"11",x"58",x"a6",x"e4"),
   111 => (x"82",x"c0",x"fe",x"4a"),
   112 => (x"05",x"9a",x"72",x"ba"),
   113 => (x"73",x"87",x"ed",x"fb"),
   114 => (x"26",x"8e",x"f0",x"48"),
   115 => (x"26",x"4c",x"26",x"4d"),
   116 => (x"0e",x"4f",x"26",x"4b"),
   117 => (x"86",x"e8",x"0e",x"5e"),
   118 => (x"c3",x"4a",x"d4",x"ff"),
   119 => (x"49",x"6a",x"7a",x"ff"),
   120 => (x"6a",x"7a",x"ff",x"c3"),
   121 => (x"c4",x"30",x"c8",x"48"),
   122 => (x"a6",x"c8",x"58",x"a6"),
   123 => (x"c3",x"b1",x"6e",x"59"),
   124 => (x"48",x"6a",x"7a",x"ff"),
   125 => (x"a6",x"cc",x"30",x"d0"),
   126 => (x"59",x"a6",x"d0",x"58"),
   127 => (x"c3",x"b1",x"66",x"c8"),
   128 => (x"48",x"6a",x"7a",x"ff"),
   129 => (x"a6",x"d4",x"30",x"d8"),
   130 => (x"59",x"a6",x"d8",x"58"),
   131 => (x"71",x"b1",x"66",x"d0"),
   132 => (x"c6",x"8e",x"e8",x"48"),
   133 => (x"26",x"4d",x"26",x"87"),
   134 => (x"26",x"4b",x"26",x"4c"),
   135 => (x"0e",x"5e",x"0e",x"4f"),
   136 => (x"d4",x"ff",x"86",x"f4"),
   137 => (x"7a",x"ff",x"c3",x"4a"),
   138 => (x"ff",x"c3",x"49",x"6a"),
   139 => (x"c8",x"48",x"71",x"7a"),
   140 => (x"58",x"a6",x"c4",x"30"),
   141 => (x"b1",x"6e",x"49",x"6a"),
   142 => (x"71",x"7a",x"ff",x"c3"),
   143 => (x"c8",x"30",x"c8",x"48"),
   144 => (x"49",x"6a",x"58",x"a6"),
   145 => (x"c3",x"b1",x"66",x"c4"),
   146 => (x"48",x"71",x"7a",x"ff"),
   147 => (x"a6",x"cc",x"30",x"c8"),
   148 => (x"c8",x"49",x"6a",x"58"),
   149 => (x"48",x"71",x"b1",x"66"),
   150 => (x"fe",x"fe",x"8e",x"f4"),
   151 => (x"5b",x"5e",x"0e",x"87"),
   152 => (x"d4",x"ff",x"0e",x"5c"),
   153 => (x"48",x"66",x"cc",x"4c"),
   154 => (x"70",x"98",x"ff",x"c3"),
   155 => (x"cc",x"d4",x"c1",x"7c"),
   156 => (x"87",x"c8",x"05",x"bf"),
   157 => (x"c9",x"48",x"66",x"d0"),
   158 => (x"58",x"a6",x"d4",x"30"),
   159 => (x"d8",x"49",x"66",x"d0"),
   160 => (x"c3",x"48",x"71",x"29"),
   161 => (x"7c",x"70",x"98",x"ff"),
   162 => (x"d0",x"49",x"66",x"d0"),
   163 => (x"c3",x"48",x"71",x"29"),
   164 => (x"7c",x"70",x"98",x"ff"),
   165 => (x"c8",x"49",x"66",x"d0"),
   166 => (x"c3",x"48",x"71",x"29"),
   167 => (x"7c",x"70",x"98",x"ff"),
   168 => (x"c3",x"48",x"66",x"d0"),
   169 => (x"7c",x"70",x"98",x"ff"),
   170 => (x"d0",x"49",x"66",x"cc"),
   171 => (x"c3",x"48",x"71",x"29"),
   172 => (x"7c",x"70",x"98",x"ff"),
   173 => (x"f0",x"c9",x"4a",x"6c"),
   174 => (x"ff",x"c3",x"4b",x"ff"),
   175 => (x"87",x"d2",x"05",x"aa"),
   176 => (x"6c",x"7c",x"ff",x"c3"),
   177 => (x"73",x"8b",x"c1",x"4a"),
   178 => (x"87",x"c6",x"02",x"9b"),
   179 => (x"02",x"aa",x"ff",x"c3"),
   180 => (x"48",x"72",x"87",x"ee"),
   181 => (x"1e",x"87",x"c0",x"fd"),
   182 => (x"d4",x"ff",x"49",x"c0"),
   183 => (x"78",x"ff",x"c3",x"48"),
   184 => (x"c8",x"c3",x"81",x"c1"),
   185 => (x"f1",x"04",x"a9",x"b7"),
   186 => (x"87",x"ef",x"fc",x"87"),
   187 => (x"0e",x"5b",x"5e",x"0e"),
   188 => (x"f8",x"c4",x"87",x"e5"),
   189 => (x"1e",x"c0",x"4b",x"df"),
   190 => (x"c1",x"f0",x"ff",x"c0"),
   191 => (x"dc",x"fd",x"1e",x"f7"),
   192 => (x"c1",x"86",x"c8",x"87"),
   193 => (x"ea",x"c0",x"05",x"a8"),
   194 => (x"48",x"d4",x"ff",x"87"),
   195 => (x"c1",x"78",x"ff",x"c3"),
   196 => (x"c0",x"c0",x"c0",x"c0"),
   197 => (x"e1",x"c0",x"1e",x"c0"),
   198 => (x"1e",x"e9",x"c1",x"f0"),
   199 => (x"c8",x"87",x"fe",x"fc"),
   200 => (x"05",x"98",x"70",x"86"),
   201 => (x"d4",x"ff",x"87",x"ca"),
   202 => (x"78",x"ff",x"c3",x"48"),
   203 => (x"87",x"cd",x"48",x"c1"),
   204 => (x"c1",x"87",x"e4",x"fe"),
   205 => (x"05",x"9b",x"73",x"8b"),
   206 => (x"c0",x"87",x"fb",x"fe"),
   207 => (x"87",x"d9",x"fb",x"48"),
   208 => (x"0e",x"5b",x"5e",x"0e"),
   209 => (x"c3",x"48",x"d4",x"ff"),
   210 => (x"e5",x"c0",x"78",x"ff"),
   211 => (x"cb",x"f4",x"1e",x"cd"),
   212 => (x"d3",x"86",x"c4",x"87"),
   213 => (x"c0",x"1e",x"c0",x"4b"),
   214 => (x"c1",x"c1",x"f0",x"ff"),
   215 => (x"87",x"fd",x"fb",x"1e"),
   216 => (x"98",x"70",x"86",x"c8"),
   217 => (x"ff",x"87",x"ca",x"05"),
   218 => (x"ff",x"c3",x"48",x"d4"),
   219 => (x"cd",x"48",x"c1",x"78"),
   220 => (x"87",x"e3",x"fd",x"87"),
   221 => (x"9b",x"73",x"8b",x"c1"),
   222 => (x"87",x"d9",x"ff",x"05"),
   223 => (x"d8",x"fa",x"48",x"c0"),
   224 => (x"5b",x"5e",x"0e",x"87"),
   225 => (x"ff",x"0e",x"5d",x"5c"),
   226 => (x"ca",x"fd",x"4d",x"d4"),
   227 => (x"1e",x"ea",x"c6",x"87"),
   228 => (x"c1",x"f0",x"e1",x"c0"),
   229 => (x"c4",x"fb",x"1e",x"c8"),
   230 => (x"70",x"86",x"c8",x"87"),
   231 => (x"d2",x"1e",x"73",x"4b"),
   232 => (x"e5",x"f3",x"1e",x"cc"),
   233 => (x"c1",x"86",x"c8",x"87"),
   234 => (x"87",x"c8",x"02",x"ab"),
   235 => (x"c0",x"87",x"d1",x"fe"),
   236 => (x"87",x"d3",x"c2",x"48"),
   237 => (x"70",x"87",x"e6",x"f9"),
   238 => (x"ff",x"ff",x"cf",x"49"),
   239 => (x"a9",x"ea",x"c6",x"99"),
   240 => (x"fd",x"87",x"c8",x"02"),
   241 => (x"48",x"c0",x"87",x"fa"),
   242 => (x"c3",x"87",x"fc",x"c1"),
   243 => (x"f1",x"c0",x"7d",x"ff"),
   244 => (x"87",x"d8",x"fc",x"4c"),
   245 => (x"c1",x"02",x"98",x"70"),
   246 => (x"1e",x"c0",x"87",x"d2"),
   247 => (x"c1",x"f0",x"ff",x"c0"),
   248 => (x"f8",x"f9",x"1e",x"fa"),
   249 => (x"70",x"86",x"c8",x"87"),
   250 => (x"05",x"9b",x"73",x"4b"),
   251 => (x"73",x"87",x"f3",x"c0"),
   252 => (x"1e",x"ca",x"d1",x"1e"),
   253 => (x"c8",x"87",x"d3",x"f2"),
   254 => (x"7d",x"ff",x"c3",x"86"),
   255 => (x"1e",x"73",x"4b",x"6d"),
   256 => (x"f2",x"1e",x"d6",x"d1"),
   257 => (x"86",x"c8",x"87",x"c4"),
   258 => (x"7d",x"7d",x"ff",x"c3"),
   259 => (x"49",x"73",x"7d",x"7d"),
   260 => (x"71",x"99",x"c0",x"c1"),
   261 => (x"87",x"c5",x"02",x"99"),
   262 => (x"ea",x"c0",x"48",x"c1"),
   263 => (x"c0",x"48",x"c0",x"87"),
   264 => (x"1e",x"73",x"87",x"e5"),
   265 => (x"f1",x"1e",x"e4",x"d1"),
   266 => (x"86",x"c8",x"87",x"e0"),
   267 => (x"cc",x"05",x"ac",x"c2"),
   268 => (x"1e",x"f0",x"d1",x"87"),
   269 => (x"c4",x"87",x"d3",x"f1"),
   270 => (x"ca",x"48",x"c0",x"86"),
   271 => (x"74",x"8c",x"c1",x"87"),
   272 => (x"cc",x"fe",x"05",x"9c"),
   273 => (x"f7",x"48",x"c0",x"87"),
   274 => (x"4d",x"43",x"87",x"cb"),
   275 => (x"20",x"38",x"35",x"44"),
   276 => (x"20",x"0a",x"64",x"25"),
   277 => (x"4d",x"43",x"00",x"20"),
   278 => (x"5f",x"38",x"35",x"44"),
   279 => (x"64",x"25",x"20",x"32"),
   280 => (x"00",x"20",x"20",x"0a"),
   281 => (x"35",x"44",x"4d",x"43"),
   282 => (x"64",x"25",x"20",x"38"),
   283 => (x"00",x"20",x"20",x"0a"),
   284 => (x"43",x"48",x"44",x"53"),
   285 => (x"69",x"6e",x"49",x"20"),
   286 => (x"6c",x"61",x"69",x"74"),
   287 => (x"74",x"61",x"7a",x"69"),
   288 => (x"20",x"6e",x"6f",x"69"),
   289 => (x"6f",x"72",x"72",x"65"),
   290 => (x"00",x"0a",x"21",x"72"),
   291 => (x"5f",x"64",x"6d",x"63"),
   292 => (x"38",x"44",x"4d",x"43"),
   293 => (x"73",x"65",x"72",x"20"),
   294 => (x"73",x"6e",x"6f",x"70"),
   295 => (x"25",x"20",x"3a",x"65"),
   296 => (x"0e",x"00",x"0a",x"64"),
   297 => (x"5d",x"5c",x"5b",x"5e"),
   298 => (x"d0",x"ff",x"1e",x"0e"),
   299 => (x"c0",x"c0",x"c8",x"4d"),
   300 => (x"cc",x"d4",x"c1",x"4b"),
   301 => (x"d6",x"78",x"c1",x"48"),
   302 => (x"df",x"ee",x"1e",x"c9"),
   303 => (x"c7",x"86",x"c4",x"87"),
   304 => (x"73",x"48",x"6d",x"4c"),
   305 => (x"58",x"a6",x"c4",x"98"),
   306 => (x"cc",x"c0",x"02",x"6e"),
   307 => (x"73",x"48",x"6d",x"87"),
   308 => (x"58",x"a6",x"c4",x"98"),
   309 => (x"f4",x"ff",x"05",x"6e"),
   310 => (x"f7",x"7d",x"c0",x"87"),
   311 => (x"48",x"6d",x"87",x"f9"),
   312 => (x"a6",x"c4",x"98",x"73"),
   313 => (x"c0",x"02",x"6e",x"58"),
   314 => (x"48",x"6d",x"87",x"cc"),
   315 => (x"a6",x"c4",x"98",x"73"),
   316 => (x"ff",x"05",x"6e",x"58"),
   317 => (x"7d",x"c1",x"87",x"f4"),
   318 => (x"e5",x"c0",x"1e",x"c0"),
   319 => (x"1e",x"c0",x"c1",x"d0"),
   320 => (x"c8",x"87",x"da",x"f5"),
   321 => (x"05",x"a8",x"c1",x"86"),
   322 => (x"c1",x"87",x"c2",x"c0"),
   323 => (x"05",x"ac",x"c2",x"4c"),
   324 => (x"d6",x"87",x"cd",x"c0"),
   325 => (x"c3",x"ed",x"1e",x"c4"),
   326 => (x"c0",x"86",x"c4",x"87"),
   327 => (x"87",x"e0",x"c1",x"48"),
   328 => (x"9c",x"74",x"8c",x"c1"),
   329 => (x"87",x"d9",x"fe",x"05"),
   330 => (x"c1",x"87",x"d6",x"f9"),
   331 => (x"c1",x"58",x"d0",x"d4"),
   332 => (x"05",x"bf",x"cc",x"d4"),
   333 => (x"c1",x"87",x"cd",x"c0"),
   334 => (x"f0",x"ff",x"c0",x"1e"),
   335 => (x"f4",x"1e",x"d0",x"c1"),
   336 => (x"86",x"c8",x"87",x"db"),
   337 => (x"c3",x"48",x"d4",x"ff"),
   338 => (x"c4",x"ca",x"78",x"ff"),
   339 => (x"d4",x"d4",x"c1",x"87"),
   340 => (x"d0",x"d4",x"c1",x"58"),
   341 => (x"cd",x"d6",x"1e",x"bf"),
   342 => (x"87",x"ee",x"ec",x"1e"),
   343 => (x"48",x"6d",x"86",x"c8"),
   344 => (x"a6",x"c4",x"98",x"73"),
   345 => (x"c0",x"02",x"6e",x"58"),
   346 => (x"48",x"6d",x"87",x"cc"),
   347 => (x"a6",x"c4",x"98",x"73"),
   348 => (x"ff",x"05",x"6e",x"58"),
   349 => (x"7d",x"c0",x"87",x"f4"),
   350 => (x"c3",x"48",x"d4",x"ff"),
   351 => (x"48",x"c1",x"78",x"ff"),
   352 => (x"87",x"d1",x"f2",x"26"),
   353 => (x"52",x"52",x"45",x"49"),
   354 => (x"49",x"50",x"53",x"00"),
   355 => (x"20",x"44",x"53",x"00"),
   356 => (x"64",x"72",x"61",x"63"),
   357 => (x"7a",x"69",x"73",x"20"),
   358 => (x"73",x"69",x"20",x"65"),
   359 => (x"0a",x"64",x"25",x"20"),
   360 => (x"5b",x"5e",x"0e",x"00"),
   361 => (x"1e",x"0e",x"5d",x"5c"),
   362 => (x"ff",x"4c",x"ff",x"c3"),
   363 => (x"7b",x"74",x"4b",x"d4"),
   364 => (x"48",x"bf",x"d0",x"ff"),
   365 => (x"98",x"c0",x"c0",x"c8"),
   366 => (x"6e",x"58",x"a6",x"c4"),
   367 => (x"87",x"d0",x"c0",x"02"),
   368 => (x"48",x"bf",x"d0",x"ff"),
   369 => (x"98",x"c0",x"c0",x"c8"),
   370 => (x"6e",x"58",x"a6",x"c4"),
   371 => (x"87",x"f0",x"ff",x"05"),
   372 => (x"c4",x"48",x"d0",x"ff"),
   373 => (x"7b",x"74",x"78",x"c1"),
   374 => (x"c0",x"1e",x"66",x"d4"),
   375 => (x"d8",x"c1",x"f0",x"ff"),
   376 => (x"87",x"f9",x"f1",x"1e"),
   377 => (x"98",x"70",x"86",x"c8"),
   378 => (x"87",x"cd",x"c0",x"02"),
   379 => (x"e9",x"1e",x"c2",x"da"),
   380 => (x"86",x"c4",x"87",x"ea"),
   381 => (x"c5",x"c2",x"48",x"c1"),
   382 => (x"c3",x"7b",x"74",x"87"),
   383 => (x"4d",x"c0",x"7b",x"fe"),
   384 => (x"49",x"bf",x"66",x"d8"),
   385 => (x"b7",x"d8",x"4a",x"71"),
   386 => (x"74",x"48",x"72",x"2a"),
   387 => (x"71",x"7b",x"70",x"98"),
   388 => (x"2a",x"b7",x"d0",x"4a"),
   389 => (x"98",x"74",x"48",x"72"),
   390 => (x"4a",x"71",x"7b",x"70"),
   391 => (x"72",x"2a",x"b7",x"c8"),
   392 => (x"70",x"98",x"74",x"48"),
   393 => (x"74",x"48",x"71",x"7b"),
   394 => (x"d8",x"7b",x"70",x"98"),
   395 => (x"80",x"c4",x"48",x"66"),
   396 => (x"c1",x"58",x"a6",x"dc"),
   397 => (x"b7",x"c0",x"c2",x"85"),
   398 => (x"c3",x"ff",x"04",x"ad"),
   399 => (x"74",x"7b",x"74",x"87"),
   400 => (x"d8",x"7b",x"74",x"7b"),
   401 => (x"74",x"49",x"e0",x"da"),
   402 => (x"c0",x"05",x"6b",x"7b"),
   403 => (x"89",x"c1",x"87",x"c8"),
   404 => (x"ff",x"05",x"99",x"71"),
   405 => (x"7b",x"74",x"87",x"f1"),
   406 => (x"48",x"bf",x"d0",x"ff"),
   407 => (x"98",x"c0",x"c0",x"c8"),
   408 => (x"6e",x"58",x"a6",x"c4"),
   409 => (x"87",x"d0",x"c0",x"02"),
   410 => (x"48",x"bf",x"d0",x"ff"),
   411 => (x"98",x"c0",x"c0",x"c8"),
   412 => (x"6e",x"58",x"a6",x"c4"),
   413 => (x"87",x"f0",x"ff",x"05"),
   414 => (x"c0",x"48",x"d0",x"ff"),
   415 => (x"ee",x"26",x"48",x"78"),
   416 => (x"72",x"57",x"87",x"d3"),
   417 => (x"20",x"65",x"74",x"69"),
   418 => (x"6c",x"69",x"61",x"66"),
   419 => (x"00",x"0a",x"64",x"65"),
   420 => (x"5c",x"5b",x"5e",x"0e"),
   421 => (x"4c",x"66",x"d0",x"0e"),
   422 => (x"c0",x"4b",x"66",x"cc"),
   423 => (x"cd",x"ee",x"c5",x"4a"),
   424 => (x"d4",x"ff",x"49",x"df"),
   425 => (x"78",x"ff",x"c3",x"48"),
   426 => (x"c3",x"48",x"bf",x"70"),
   427 => (x"c1",x"05",x"a8",x"fe"),
   428 => (x"d4",x"c1",x"87",x"d8"),
   429 => (x"78",x"c0",x"48",x"c8"),
   430 => (x"04",x"ac",x"b7",x"c4"),
   431 => (x"ec",x"87",x"dc",x"c0"),
   432 => (x"49",x"70",x"87",x"d1"),
   433 => (x"83",x"c4",x"7b",x"71"),
   434 => (x"bf",x"c8",x"d4",x"c1"),
   435 => (x"c1",x"80",x"71",x"48"),
   436 => (x"c4",x"58",x"cc",x"d4"),
   437 => (x"03",x"ac",x"b7",x"8c"),
   438 => (x"c0",x"87",x"e4",x"ff"),
   439 => (x"c0",x"06",x"ac",x"b7"),
   440 => (x"d4",x"ff",x"87",x"e5"),
   441 => (x"78",x"ff",x"c3",x"48"),
   442 => (x"71",x"49",x"bf",x"70"),
   443 => (x"ff",x"c3",x"7b",x"97"),
   444 => (x"c1",x"83",x"c1",x"98"),
   445 => (x"48",x"bf",x"c8",x"d4"),
   446 => (x"d4",x"c1",x"80",x"71"),
   447 => (x"8c",x"c1",x"58",x"cc"),
   448 => (x"01",x"ac",x"b7",x"c0"),
   449 => (x"c1",x"87",x"db",x"ff"),
   450 => (x"89",x"c1",x"4a",x"49"),
   451 => (x"fe",x"05",x"99",x"71"),
   452 => (x"d4",x"ff",x"87",x"d0"),
   453 => (x"78",x"ff",x"c3",x"48"),
   454 => (x"fa",x"eb",x"48",x"72"),
   455 => (x"5b",x"5e",x"0e",x"87"),
   456 => (x"c8",x"1e",x"0e",x"5c"),
   457 => (x"c0",x"4c",x"c0",x"c0"),
   458 => (x"48",x"d4",x"ff",x"4b"),
   459 => (x"ff",x"78",x"ff",x"c3"),
   460 => (x"74",x"48",x"bf",x"d0"),
   461 => (x"58",x"a6",x"c4",x"98"),
   462 => (x"ce",x"c0",x"02",x"6e"),
   463 => (x"bf",x"d0",x"ff",x"87"),
   464 => (x"c4",x"98",x"74",x"48"),
   465 => (x"05",x"6e",x"58",x"a6"),
   466 => (x"ff",x"87",x"f2",x"ff"),
   467 => (x"c1",x"c4",x"48",x"d0"),
   468 => (x"48",x"d4",x"ff",x"78"),
   469 => (x"d0",x"78",x"ff",x"c3"),
   470 => (x"ff",x"c0",x"1e",x"66"),
   471 => (x"1e",x"d1",x"c1",x"f0"),
   472 => (x"c8",x"87",x"fa",x"eb"),
   473 => (x"71",x"49",x"70",x"86"),
   474 => (x"d0",x"c0",x"02",x"99"),
   475 => (x"d4",x"1e",x"71",x"87"),
   476 => (x"f1",x"de",x"1e",x"66"),
   477 => (x"87",x"d2",x"e4",x"1e"),
   478 => (x"ee",x"c0",x"86",x"cc"),
   479 => (x"1e",x"c0",x"c8",x"87"),
   480 => (x"fc",x"1e",x"66",x"d8"),
   481 => (x"86",x"c8",x"87",x"ca"),
   482 => (x"d0",x"ff",x"4b",x"70"),
   483 => (x"98",x"74",x"48",x"bf"),
   484 => (x"6e",x"58",x"a6",x"c4"),
   485 => (x"87",x"ce",x"c0",x"02"),
   486 => (x"48",x"bf",x"d0",x"ff"),
   487 => (x"a6",x"c4",x"98",x"74"),
   488 => (x"ff",x"05",x"6e",x"58"),
   489 => (x"d0",x"ff",x"87",x"f2"),
   490 => (x"73",x"78",x"c0",x"48"),
   491 => (x"e6",x"e9",x"26",x"48"),
   492 => (x"61",x"65",x"52",x"87"),
   493 => (x"6f",x"63",x"20",x"64"),
   494 => (x"6e",x"61",x"6d",x"6d"),
   495 => (x"61",x"66",x"20",x"64"),
   496 => (x"64",x"65",x"6c",x"69"),
   497 => (x"20",x"74",x"61",x"20"),
   498 => (x"28",x"20",x"64",x"25"),
   499 => (x"0a",x"29",x"64",x"25"),
   500 => (x"5b",x"5e",x"0e",x"00"),
   501 => (x"1e",x"0e",x"5d",x"5c"),
   502 => (x"ff",x"c0",x"1e",x"c0"),
   503 => (x"1e",x"c9",x"c1",x"f0"),
   504 => (x"c8",x"87",x"fa",x"e9"),
   505 => (x"c1",x"1e",x"d2",x"86"),
   506 => (x"fa",x"1e",x"da",x"d4"),
   507 => (x"86",x"c8",x"87",x"e2"),
   508 => (x"85",x"c1",x"4d",x"c0"),
   509 => (x"04",x"ad",x"b7",x"d2"),
   510 => (x"c1",x"87",x"f7",x"ff"),
   511 => (x"bf",x"97",x"da",x"d4"),
   512 => (x"99",x"c0",x"c3",x"49"),
   513 => (x"05",x"a9",x"c0",x"c1"),
   514 => (x"c1",x"87",x"e8",x"c0"),
   515 => (x"bf",x"97",x"e1",x"d4"),
   516 => (x"c1",x"31",x"d0",x"49"),
   517 => (x"bf",x"97",x"e2",x"d4"),
   518 => (x"72",x"32",x"c8",x"4a"),
   519 => (x"e3",x"d4",x"c1",x"b1"),
   520 => (x"72",x"4a",x"bf",x"97"),
   521 => (x"ff",x"ff",x"cf",x"b1"),
   522 => (x"4d",x"71",x"99",x"ff"),
   523 => (x"35",x"ca",x"85",x"c1"),
   524 => (x"c1",x"87",x"f0",x"c2"),
   525 => (x"bf",x"97",x"e3",x"d4"),
   526 => (x"c6",x"33",x"c1",x"4b"),
   527 => (x"e4",x"d4",x"c1",x"9b"),
   528 => (x"c7",x"49",x"bf",x"97"),
   529 => (x"b3",x"71",x"29",x"b7"),
   530 => (x"97",x"df",x"d4",x"c1"),
   531 => (x"48",x"71",x"49",x"bf"),
   532 => (x"a6",x"c4",x"98",x"cf"),
   533 => (x"e0",x"d4",x"c1",x"58"),
   534 => (x"c3",x"4c",x"bf",x"97"),
   535 => (x"c1",x"34",x"ca",x"9c"),
   536 => (x"bf",x"97",x"e1",x"d4"),
   537 => (x"71",x"31",x"c2",x"49"),
   538 => (x"e2",x"d4",x"c1",x"b4"),
   539 => (x"c3",x"49",x"bf",x"97"),
   540 => (x"b7",x"c6",x"99",x"c0"),
   541 => (x"74",x"b4",x"71",x"29"),
   542 => (x"1e",x"66",x"c4",x"1e"),
   543 => (x"e3",x"c0",x"1e",x"73"),
   544 => (x"c5",x"e0",x"1e",x"e9"),
   545 => (x"c2",x"86",x"d0",x"87"),
   546 => (x"73",x"48",x"c1",x"83"),
   547 => (x"73",x"4b",x"70",x"30"),
   548 => (x"d6",x"e4",x"c0",x"1e"),
   549 => (x"f1",x"df",x"ff",x"1e"),
   550 => (x"c1",x"86",x"c8",x"87"),
   551 => (x"c4",x"30",x"6e",x"48"),
   552 => (x"49",x"74",x"58",x"a6"),
   553 => (x"4d",x"71",x"81",x"c1"),
   554 => (x"6e",x"95",x"b7",x"73"),
   555 => (x"c0",x"1e",x"75",x"1e"),
   556 => (x"ff",x"1e",x"df",x"e4"),
   557 => (x"cc",x"87",x"d3",x"df"),
   558 => (x"c8",x"48",x"6e",x"86"),
   559 => (x"06",x"a8",x"b7",x"c0"),
   560 => (x"c1",x"87",x"d4",x"c0"),
   561 => (x"c1",x"48",x"6e",x"35"),
   562 => (x"a6",x"c4",x"28",x"b7"),
   563 => (x"c8",x"48",x"6e",x"58"),
   564 => (x"01",x"a8",x"b7",x"c0"),
   565 => (x"75",x"87",x"ec",x"ff"),
   566 => (x"f5",x"e4",x"c0",x"1e"),
   567 => (x"e9",x"de",x"ff",x"1e"),
   568 => (x"75",x"86",x"c8",x"87"),
   569 => (x"ec",x"e4",x"26",x"48"),
   570 => (x"73",x"5f",x"63",x"87"),
   571 => (x"5f",x"65",x"7a",x"69"),
   572 => (x"74",x"6c",x"75",x"6d"),
   573 => (x"64",x"25",x"20",x"3a"),
   574 => (x"65",x"72",x"20",x"2c"),
   575 => (x"62",x"5f",x"64",x"61"),
   576 => (x"65",x"6c",x"5f",x"6c"),
   577 => (x"25",x"20",x"3a",x"6e"),
   578 => (x"63",x"20",x"2c",x"64"),
   579 => (x"65",x"7a",x"69",x"73"),
   580 => (x"64",x"25",x"20",x"3a"),
   581 => (x"75",x"4d",x"00",x"0a"),
   582 => (x"25",x"20",x"74",x"6c"),
   583 => (x"25",x"00",x"0a",x"64"),
   584 => (x"6c",x"62",x"20",x"64"),
   585 => (x"73",x"6b",x"63",x"6f"),
   586 => (x"20",x"66",x"6f",x"20"),
   587 => (x"65",x"7a",x"69",x"73"),
   588 => (x"0a",x"64",x"25",x"20"),
   589 => (x"20",x"64",x"25",x"00"),
   590 => (x"63",x"6f",x"6c",x"62"),
   591 => (x"6f",x"20",x"73",x"6b"),
   592 => (x"31",x"35",x"20",x"66"),
   593 => (x"79",x"62",x"20",x"32"),
   594 => (x"0a",x"73",x"65",x"74"),
   595 => (x"44",x"4d",x"43",x"00"),
   596 => (x"5b",x"5e",x"0e",x"00"),
   597 => (x"d0",x"4b",x"c0",x"0e"),
   598 => (x"b7",x"c0",x"48",x"66"),
   599 => (x"f6",x"c0",x"06",x"a8"),
   600 => (x"97",x"66",x"c8",x"87"),
   601 => (x"c0",x"fe",x"4a",x"bf"),
   602 => (x"66",x"c8",x"ba",x"82"),
   603 => (x"cc",x"80",x"c1",x"48"),
   604 => (x"66",x"cc",x"58",x"a6"),
   605 => (x"fe",x"49",x"bf",x"97"),
   606 => (x"cc",x"b9",x"81",x"c0"),
   607 => (x"80",x"c1",x"48",x"66"),
   608 => (x"71",x"58",x"a6",x"d0"),
   609 => (x"c4",x"02",x"aa",x"b7"),
   610 => (x"cc",x"48",x"c1",x"87"),
   611 => (x"d0",x"83",x"c1",x"87"),
   612 => (x"04",x"ab",x"b7",x"66"),
   613 => (x"c0",x"87",x"ca",x"ff"),
   614 => (x"26",x"87",x"c4",x"48"),
   615 => (x"26",x"4c",x"26",x"4d"),
   616 => (x"0e",x"4f",x"26",x"4b"),
   617 => (x"5d",x"5c",x"5b",x"5e"),
   618 => (x"f4",x"dc",x"c1",x"0e"),
   619 => (x"c1",x"78",x"c0",x"48"),
   620 => (x"ff",x"1e",x"fd",x"c0"),
   621 => (x"c4",x"87",x"e5",x"da"),
   622 => (x"ec",x"d4",x"c1",x"86"),
   623 => (x"f5",x"1e",x"c0",x"1e"),
   624 => (x"86",x"c8",x"87",x"db"),
   625 => (x"cf",x"05",x"98",x"70"),
   626 => (x"e9",x"fd",x"c0",x"87"),
   627 => (x"cb",x"da",x"ff",x"1e"),
   628 => (x"c0",x"86",x"c4",x"87"),
   629 => (x"87",x"d6",x"cb",x"48"),
   630 => (x"1e",x"ca",x"c1",x"c1"),
   631 => (x"87",x"fc",x"d9",x"ff"),
   632 => (x"4b",x"c0",x"86",x"c4"),
   633 => (x"48",x"e0",x"dd",x"c1"),
   634 => (x"1e",x"c8",x"78",x"c1"),
   635 => (x"1e",x"e1",x"c1",x"c1"),
   636 => (x"1e",x"e2",x"d5",x"c1"),
   637 => (x"cc",x"87",x"da",x"fd"),
   638 => (x"05",x"98",x"70",x"86"),
   639 => (x"dd",x"c1",x"87",x"c6"),
   640 => (x"78",x"c0",x"48",x"e0"),
   641 => (x"c1",x"c1",x"1e",x"c8"),
   642 => (x"d5",x"c1",x"1e",x"ea"),
   643 => (x"c0",x"fd",x"1e",x"fe"),
   644 => (x"70",x"86",x"cc",x"87"),
   645 => (x"87",x"c6",x"05",x"98"),
   646 => (x"48",x"e0",x"dd",x"c1"),
   647 => (x"dd",x"c1",x"78",x"c0"),
   648 => (x"c1",x"1e",x"bf",x"e0"),
   649 => (x"ff",x"1e",x"f3",x"c1"),
   650 => (x"c8",x"87",x"df",x"d9"),
   651 => (x"e0",x"dd",x"c1",x"86"),
   652 => (x"d8",x"c2",x"02",x"bf"),
   653 => (x"ec",x"d4",x"c1",x"87"),
   654 => (x"ea",x"db",x"c1",x"4d"),
   655 => (x"ea",x"dc",x"c1",x"4c"),
   656 => (x"71",x"49",x"bf",x"9f"),
   657 => (x"ea",x"dc",x"c1",x"1e"),
   658 => (x"ec",x"d4",x"c1",x"49"),
   659 => (x"d0",x"1e",x"71",x"89"),
   660 => (x"1e",x"c0",x"c8",x"1e"),
   661 => (x"1e",x"db",x"fe",x"c0"),
   662 => (x"87",x"ee",x"d8",x"ff"),
   663 => (x"49",x"74",x"86",x"d4"),
   664 => (x"4b",x"69",x"81",x"c8"),
   665 => (x"9f",x"ea",x"dc",x"c1"),
   666 => (x"d6",x"c5",x"49",x"bf"),
   667 => (x"c0",x"05",x"a9",x"ea"),
   668 => (x"49",x"74",x"87",x"d0"),
   669 => (x"1e",x"69",x"81",x"c8"),
   670 => (x"c4",x"87",x"d9",x"d9"),
   671 => (x"c0",x"4b",x"70",x"86"),
   672 => (x"49",x"75",x"87",x"df"),
   673 => (x"9f",x"81",x"fe",x"c7"),
   674 => (x"e9",x"ca",x"49",x"69"),
   675 => (x"c0",x"02",x"a9",x"d5"),
   676 => (x"fd",x"c0",x"87",x"cf"),
   677 => (x"d7",x"ff",x"1e",x"fd"),
   678 => (x"86",x"c4",x"87",x"c2"),
   679 => (x"cd",x"c8",x"48",x"c0"),
   680 => (x"c0",x"1e",x"73",x"87"),
   681 => (x"ff",x"1e",x"d8",x"ff"),
   682 => (x"c8",x"87",x"df",x"d7"),
   683 => (x"ec",x"d4",x"c1",x"86"),
   684 => (x"f1",x"1e",x"73",x"1e"),
   685 => (x"86",x"c8",x"87",x"e7"),
   686 => (x"c0",x"05",x"98",x"70"),
   687 => (x"48",x"c0",x"87",x"c5"),
   688 => (x"c0",x"87",x"eb",x"c7"),
   689 => (x"ff",x"1e",x"f0",x"ff"),
   690 => (x"c4",x"87",x"d1",x"d6"),
   691 => (x"c6",x"c2",x"c1",x"86"),
   692 => (x"f5",x"d6",x"ff",x"1e"),
   693 => (x"c8",x"86",x"c4",x"87"),
   694 => (x"de",x"c2",x"c1",x"1e"),
   695 => (x"fe",x"d5",x"c1",x"1e"),
   696 => (x"87",x"ed",x"f9",x"1e"),
   697 => (x"98",x"70",x"86",x"cc"),
   698 => (x"87",x"c9",x"c0",x"05"),
   699 => (x"48",x"f4",x"dc",x"c1"),
   700 => (x"e4",x"c0",x"78",x"c1"),
   701 => (x"c1",x"1e",x"c8",x"87"),
   702 => (x"c1",x"1e",x"e7",x"c2"),
   703 => (x"f9",x"1e",x"e2",x"d5"),
   704 => (x"86",x"cc",x"87",x"cf"),
   705 => (x"c0",x"02",x"98",x"70"),
   706 => (x"c0",x"c1",x"87",x"cf"),
   707 => (x"d5",x"ff",x"1e",x"d7"),
   708 => (x"86",x"c4",x"87",x"f8"),
   709 => (x"d5",x"c6",x"48",x"c0"),
   710 => (x"ea",x"dc",x"c1",x"87"),
   711 => (x"c1",x"49",x"bf",x"97"),
   712 => (x"c0",x"05",x"a9",x"d5"),
   713 => (x"dc",x"c1",x"87",x"cd"),
   714 => (x"49",x"bf",x"97",x"eb"),
   715 => (x"02",x"a9",x"ea",x"c2"),
   716 => (x"c0",x"87",x"c5",x"c0"),
   717 => (x"87",x"f6",x"c5",x"48"),
   718 => (x"97",x"ec",x"d4",x"c1"),
   719 => (x"e9",x"c3",x"49",x"bf"),
   720 => (x"d2",x"c0",x"02",x"a9"),
   721 => (x"ec",x"d4",x"c1",x"87"),
   722 => (x"c3",x"49",x"bf",x"97"),
   723 => (x"c0",x"02",x"a9",x"eb"),
   724 => (x"48",x"c0",x"87",x"c5"),
   725 => (x"c1",x"87",x"d7",x"c5"),
   726 => (x"bf",x"97",x"f7",x"d4"),
   727 => (x"05",x"99",x"71",x"49"),
   728 => (x"c1",x"87",x"cc",x"c0"),
   729 => (x"bf",x"97",x"f8",x"d4"),
   730 => (x"02",x"a9",x"c2",x"49"),
   731 => (x"c0",x"87",x"c5",x"c0"),
   732 => (x"87",x"fa",x"c4",x"48"),
   733 => (x"97",x"f9",x"d4",x"c1"),
   734 => (x"dc",x"c1",x"48",x"bf"),
   735 => (x"dc",x"c1",x"58",x"f0"),
   736 => (x"71",x"49",x"bf",x"ec"),
   737 => (x"c1",x"8a",x"c1",x"4a"),
   738 => (x"72",x"5a",x"f4",x"dc"),
   739 => (x"c1",x"1e",x"71",x"1e"),
   740 => (x"ff",x"1e",x"f0",x"c2"),
   741 => (x"cc",x"87",x"f3",x"d3"),
   742 => (x"fa",x"d4",x"c1",x"86"),
   743 => (x"73",x"49",x"bf",x"97"),
   744 => (x"fb",x"d4",x"c1",x"81"),
   745 => (x"c8",x"4a",x"bf",x"97"),
   746 => (x"71",x"48",x"72",x"32"),
   747 => (x"c4",x"dd",x"c1",x"80"),
   748 => (x"fc",x"d4",x"c1",x"58"),
   749 => (x"c1",x"48",x"bf",x"97"),
   750 => (x"c1",x"58",x"d8",x"dd"),
   751 => (x"02",x"bf",x"f4",x"dc"),
   752 => (x"c8",x"87",x"da",x"c2"),
   753 => (x"f4",x"c0",x"c1",x"1e"),
   754 => (x"fe",x"d5",x"c1",x"1e"),
   755 => (x"87",x"c1",x"f6",x"1e"),
   756 => (x"98",x"70",x"86",x"cc"),
   757 => (x"87",x"c5",x"c0",x"02"),
   758 => (x"d1",x"c3",x"48",x"c0"),
   759 => (x"ec",x"dc",x"c1",x"87"),
   760 => (x"48",x"72",x"4a",x"bf"),
   761 => (x"dd",x"c1",x"30",x"c4"),
   762 => (x"dd",x"c1",x"58",x"dc"),
   763 => (x"d5",x"c1",x"5a",x"d4"),
   764 => (x"49",x"bf",x"97",x"d1"),
   765 => (x"d5",x"c1",x"31",x"c8"),
   766 => (x"4b",x"bf",x"97",x"d0"),
   767 => (x"d5",x"c1",x"81",x"73"),
   768 => (x"4b",x"bf",x"97",x"d2"),
   769 => (x"81",x"73",x"33",x"d0"),
   770 => (x"97",x"d3",x"d5",x"c1"),
   771 => (x"33",x"d8",x"4b",x"bf"),
   772 => (x"dd",x"c1",x"81",x"73"),
   773 => (x"dd",x"c1",x"59",x"e0"),
   774 => (x"c1",x"91",x"bf",x"d4"),
   775 => (x"81",x"bf",x"c0",x"dd"),
   776 => (x"59",x"c8",x"dd",x"c1"),
   777 => (x"97",x"d9",x"d5",x"c1"),
   778 => (x"33",x"c8",x"4b",x"bf"),
   779 => (x"97",x"d8",x"d5",x"c1"),
   780 => (x"83",x"74",x"4c",x"bf"),
   781 => (x"97",x"da",x"d5",x"c1"),
   782 => (x"34",x"d0",x"4c",x"bf"),
   783 => (x"d5",x"c1",x"83",x"74"),
   784 => (x"4c",x"bf",x"97",x"db"),
   785 => (x"34",x"d8",x"9c",x"cf"),
   786 => (x"dd",x"c1",x"83",x"74"),
   787 => (x"8b",x"c2",x"5b",x"cc"),
   788 => (x"48",x"72",x"92",x"73"),
   789 => (x"dd",x"c1",x"80",x"71"),
   790 => (x"cf",x"c1",x"58",x"d0"),
   791 => (x"fe",x"d4",x"c1",x"87"),
   792 => (x"c8",x"49",x"bf",x"97"),
   793 => (x"fd",x"d4",x"c1",x"31"),
   794 => (x"72",x"4a",x"bf",x"97"),
   795 => (x"dc",x"dd",x"c1",x"81"),
   796 => (x"c7",x"31",x"c5",x"59"),
   797 => (x"29",x"c9",x"81",x"ff"),
   798 => (x"59",x"d4",x"dd",x"c1"),
   799 => (x"97",x"c3",x"d5",x"c1"),
   800 => (x"32",x"c8",x"4a",x"bf"),
   801 => (x"97",x"c2",x"d5",x"c1"),
   802 => (x"82",x"73",x"4b",x"bf"),
   803 => (x"5a",x"e0",x"dd",x"c1"),
   804 => (x"bf",x"d4",x"dd",x"c1"),
   805 => (x"c0",x"dd",x"c1",x"92"),
   806 => (x"dd",x"c1",x"82",x"bf"),
   807 => (x"dd",x"c1",x"5a",x"d0"),
   808 => (x"78",x"c0",x"48",x"c8"),
   809 => (x"80",x"71",x"48",x"72"),
   810 => (x"58",x"c8",x"dd",x"c1"),
   811 => (x"ea",x"f3",x"48",x"c1"),
   812 => (x"5b",x"5e",x"0e",x"87"),
   813 => (x"dc",x"c1",x"0e",x"5c"),
   814 => (x"c0",x"02",x"bf",x"f4"),
   815 => (x"66",x"cc",x"87",x"cf"),
   816 => (x"2a",x"b7",x"c7",x"4a"),
   817 => (x"c1",x"4b",x"66",x"cc"),
   818 => (x"cc",x"c0",x"9b",x"ff"),
   819 => (x"4a",x"66",x"cc",x"87"),
   820 => (x"cc",x"2a",x"b7",x"c8"),
   821 => (x"ff",x"c3",x"4b",x"66"),
   822 => (x"ec",x"d4",x"c1",x"9b"),
   823 => (x"c0",x"dd",x"c1",x"1e"),
   824 => (x"81",x"72",x"49",x"bf"),
   825 => (x"f4",x"e8",x"1e",x"71"),
   826 => (x"70",x"86",x"c8",x"87"),
   827 => (x"c5",x"c0",x"05",x"98"),
   828 => (x"c0",x"48",x"c0",x"87"),
   829 => (x"dc",x"c1",x"87",x"ea"),
   830 => (x"c0",x"02",x"bf",x"f4"),
   831 => (x"49",x"73",x"87",x"d4"),
   832 => (x"c1",x"91",x"b7",x"c4"),
   833 => (x"69",x"81",x"ec",x"d4"),
   834 => (x"ff",x"ff",x"cf",x"4c"),
   835 => (x"c0",x"9c",x"ff",x"ff"),
   836 => (x"49",x"73",x"87",x"cc"),
   837 => (x"c1",x"91",x"b7",x"c2"),
   838 => (x"9f",x"81",x"ec",x"d4"),
   839 => (x"48",x"74",x"4c",x"69"),
   840 => (x"0e",x"87",x"fa",x"f1"),
   841 => (x"5d",x"5c",x"5b",x"5e"),
   842 => (x"c0",x"86",x"f4",x"0e"),
   843 => (x"c1",x"48",x"76",x"4b"),
   844 => (x"78",x"bf",x"c8",x"dd"),
   845 => (x"dd",x"c1",x"80",x"c4"),
   846 => (x"c1",x"78",x"bf",x"cc"),
   847 => (x"02",x"bf",x"f4",x"dc"),
   848 => (x"c1",x"87",x"ca",x"c0"),
   849 => (x"49",x"bf",x"ec",x"dc"),
   850 => (x"c7",x"c0",x"31",x"c4"),
   851 => (x"d0",x"dd",x"c1",x"87"),
   852 => (x"31",x"c4",x"49",x"bf"),
   853 => (x"c0",x"59",x"a6",x"cc"),
   854 => (x"48",x"66",x"c8",x"4d"),
   855 => (x"c2",x"06",x"a8",x"c0"),
   856 => (x"49",x"75",x"87",x"f5"),
   857 => (x"99",x"71",x"99",x"cf"),
   858 => (x"87",x"db",x"c0",x"05"),
   859 => (x"1e",x"ec",x"d4",x"c1"),
   860 => (x"48",x"49",x"66",x"c8"),
   861 => (x"a6",x"cc",x"80",x"c1"),
   862 => (x"e6",x"1e",x"71",x"58"),
   863 => (x"86",x"c8",x"87",x"df"),
   864 => (x"4b",x"ec",x"d4",x"c1"),
   865 => (x"c0",x"87",x"c3",x"c0"),
   866 => (x"6b",x"97",x"83",x"e0"),
   867 => (x"02",x"99",x"71",x"49"),
   868 => (x"97",x"87",x"fb",x"c1"),
   869 => (x"e5",x"c3",x"49",x"6b"),
   870 => (x"f1",x"c1",x"02",x"a9"),
   871 => (x"cb",x"49",x"73",x"87"),
   872 => (x"49",x"69",x"97",x"81"),
   873 => (x"99",x"71",x"99",x"d8"),
   874 => (x"87",x"e2",x"c1",x"05"),
   875 => (x"ca",x"ff",x"1e",x"73"),
   876 => (x"86",x"c4",x"87",x"ea"),
   877 => (x"e4",x"c0",x"1e",x"cb"),
   878 => (x"1e",x"73",x"1e",x"66"),
   879 => (x"cc",x"87",x"d2",x"ee"),
   880 => (x"05",x"98",x"70",x"86"),
   881 => (x"73",x"87",x"c7",x"c1"),
   882 => (x"dc",x"82",x"dc",x"4a"),
   883 => (x"81",x"c4",x"49",x"66"),
   884 => (x"4a",x"73",x"79",x"6a"),
   885 => (x"66",x"dc",x"82",x"da"),
   886 => (x"9f",x"81",x"c8",x"49"),
   887 => (x"79",x"70",x"48",x"6a"),
   888 => (x"dc",x"c1",x"4c",x"71"),
   889 => (x"c0",x"02",x"bf",x"f4"),
   890 => (x"49",x"73",x"87",x"d2"),
   891 => (x"69",x"9f",x"81",x"d4"),
   892 => (x"ff",x"ff",x"c0",x"49"),
   893 => (x"d0",x"4a",x"71",x"99"),
   894 => (x"87",x"c2",x"c0",x"32"),
   895 => (x"48",x"72",x"4a",x"c0"),
   896 => (x"7c",x"70",x"80",x"6c"),
   897 => (x"c0",x"48",x"66",x"dc"),
   898 => (x"c1",x"48",x"c1",x"78"),
   899 => (x"85",x"c1",x"87",x"c0"),
   900 => (x"04",x"ad",x"66",x"c8"),
   901 => (x"c1",x"87",x"cb",x"fd"),
   902 => (x"02",x"bf",x"f4",x"dc"),
   903 => (x"6e",x"87",x"ed",x"c0"),
   904 => (x"87",x"cd",x"fa",x"1e"),
   905 => (x"a6",x"c4",x"86",x"c4"),
   906 => (x"cf",x"49",x"6e",x"58"),
   907 => (x"f8",x"ff",x"ff",x"ff"),
   908 => (x"c0",x"02",x"a9",x"99"),
   909 => (x"49",x"6e",x"87",x"d6"),
   910 => (x"dc",x"c1",x"89",x"c2"),
   911 => (x"c1",x"91",x"bf",x"ec"),
   912 => (x"48",x"bf",x"c4",x"dd"),
   913 => (x"a6",x"c8",x"80",x"71"),
   914 => (x"87",x"cb",x"fc",x"58"),
   915 => (x"8e",x"f4",x"48",x"c0"),
   916 => (x"0e",x"87",x"c8",x"ed"),
   917 => (x"c8",x"0e",x"5b",x"5e"),
   918 => (x"c1",x"49",x"bf",x"66"),
   919 => (x"09",x"66",x"c8",x"81"),
   920 => (x"dc",x"c1",x"09",x"79"),
   921 => (x"71",x"99",x"bf",x"f0"),
   922 => (x"d0",x"c0",x"05",x"99"),
   923 => (x"4b",x"66",x"c8",x"87"),
   924 => (x"1e",x"6b",x"83",x"c8"),
   925 => (x"c4",x"87",x"fa",x"f8"),
   926 => (x"71",x"49",x"70",x"86"),
   927 => (x"ec",x"48",x"c1",x"7b"),
   928 => (x"5e",x"0e",x"87",x"dd"),
   929 => (x"c4",x"dd",x"c1",x"0e"),
   930 => (x"66",x"c4",x"49",x"bf"),
   931 => (x"6a",x"82",x"c8",x"4a"),
   932 => (x"c1",x"8a",x"c2",x"4a"),
   933 => (x"92",x"bf",x"ec",x"dc"),
   934 => (x"dc",x"c1",x"81",x"72"),
   935 => (x"c4",x"4a",x"bf",x"f0"),
   936 => (x"72",x"9a",x"bf",x"66"),
   937 => (x"1e",x"66",x"c8",x"81"),
   938 => (x"f0",x"e1",x"1e",x"71"),
   939 => (x"70",x"86",x"c8",x"87"),
   940 => (x"c5",x"c0",x"05",x"98"),
   941 => (x"c0",x"48",x"c0",x"87"),
   942 => (x"48",x"c1",x"87",x"c2"),
   943 => (x"0e",x"87",x"e2",x"eb"),
   944 => (x"0e",x"5c",x"5b",x"5e"),
   945 => (x"c1",x"1e",x"66",x"cc"),
   946 => (x"f9",x"1e",x"e4",x"dd"),
   947 => (x"86",x"c8",x"87",x"d5"),
   948 => (x"c1",x"02",x"98",x"70"),
   949 => (x"dd",x"c1",x"87",x"d4"),
   950 => (x"c7",x"49",x"bf",x"e8"),
   951 => (x"29",x"c9",x"81",x"ff"),
   952 => (x"4b",x"c0",x"4c",x"71"),
   953 => (x"1e",x"c1",x"fd",x"c0"),
   954 => (x"87",x"f0",x"c5",x"ff"),
   955 => (x"b7",x"c0",x"86",x"c4"),
   956 => (x"c7",x"c1",x"06",x"ac"),
   957 => (x"1e",x"66",x"d0",x"87"),
   958 => (x"1e",x"e4",x"dd",x"c1"),
   959 => (x"c8",x"87",x"c3",x"fe"),
   960 => (x"05",x"98",x"70",x"86"),
   961 => (x"c0",x"87",x"c5",x"c0"),
   962 => (x"87",x"f2",x"c0",x"48"),
   963 => (x"1e",x"e4",x"dd",x"c1"),
   964 => (x"c4",x"87",x"c0",x"fd"),
   965 => (x"48",x"66",x"d0",x"86"),
   966 => (x"d4",x"80",x"c0",x"c8"),
   967 => (x"83",x"c1",x"58",x"a6"),
   968 => (x"04",x"ab",x"b7",x"74"),
   969 => (x"c0",x"87",x"ce",x"ff"),
   970 => (x"66",x"cc",x"87",x"d2"),
   971 => (x"da",x"fd",x"c0",x"1e"),
   972 => (x"d5",x"c5",x"ff",x"1e"),
   973 => (x"c0",x"86",x"c8",x"87"),
   974 => (x"87",x"c2",x"c0",x"48"),
   975 => (x"dc",x"e9",x"48",x"c1"),
   976 => (x"65",x"70",x"4f",x"87"),
   977 => (x"20",x"64",x"65",x"6e"),
   978 => (x"65",x"6c",x"69",x"66"),
   979 => (x"6f",x"6c",x"20",x"2c"),
   980 => (x"6e",x"69",x"64",x"61"),
   981 => (x"2e",x"2e",x"2e",x"67"),
   982 => (x"61",x"43",x"00",x"0a"),
   983 => (x"20",x"74",x"27",x"6e"),
   984 => (x"6e",x"65",x"70",x"6f"),
   985 => (x"0a",x"73",x"25",x"20"),
   986 => (x"61",x"65",x"52",x"00"),
   987 => (x"66",x"6f",x"20",x"64"),
   988 => (x"52",x"42",x"4d",x"20"),
   989 => (x"69",x"61",x"66",x"20"),
   990 => (x"0a",x"64",x"65",x"6c"),
   991 => (x"20",x"6f",x"4e",x"00"),
   992 => (x"74",x"72",x"61",x"70"),
   993 => (x"6f",x"69",x"74",x"69"),
   994 => (x"69",x"73",x"20",x"6e"),
   995 => (x"74",x"61",x"6e",x"67"),
   996 => (x"20",x"65",x"72",x"75"),
   997 => (x"6e",x"75",x"6f",x"66"),
   998 => (x"4d",x"00",x"0a",x"64"),
   999 => (x"69",x"73",x"52",x"42"),
  1000 => (x"20",x"3a",x"65",x"7a"),
  1001 => (x"20",x"2c",x"64",x"25"),
  1002 => (x"74",x"72",x"61",x"70"),
  1003 => (x"6f",x"69",x"74",x"69"),
  1004 => (x"7a",x"69",x"73",x"6e"),
  1005 => (x"25",x"20",x"3a",x"65"),
  1006 => (x"6f",x"20",x"2c",x"64"),
  1007 => (x"65",x"73",x"66",x"66"),
  1008 => (x"66",x"6f",x"20",x"74"),
  1009 => (x"67",x"69",x"73",x"20"),
  1010 => (x"64",x"25",x"20",x"3a"),
  1011 => (x"69",x"73",x"20",x"2c"),
  1012 => (x"78",x"30",x"20",x"67"),
  1013 => (x"00",x"0a",x"78",x"25"),
  1014 => (x"64",x"61",x"65",x"52"),
  1015 => (x"20",x"67",x"6e",x"69"),
  1016 => (x"74",x"6f",x"6f",x"62"),
  1017 => (x"63",x"65",x"73",x"20"),
  1018 => (x"20",x"72",x"6f",x"74"),
  1019 => (x"00",x"0a",x"64",x"25"),
  1020 => (x"64",x"61",x"65",x"52"),
  1021 => (x"6f",x"6f",x"62",x"20"),
  1022 => (x"65",x"73",x"20",x"74"),
  1023 => (x"72",x"6f",x"74",x"63"),
  1024 => (x"6f",x"72",x"66",x"20"),
  1025 => (x"69",x"66",x"20",x"6d"),
  1026 => (x"20",x"74",x"73",x"72"),
  1027 => (x"74",x"72",x"61",x"70"),
  1028 => (x"6f",x"69",x"74",x"69"),
  1029 => (x"55",x"00",x"0a",x"6e"),
  1030 => (x"70",x"75",x"73",x"6e"),
  1031 => (x"74",x"72",x"6f",x"70"),
  1032 => (x"70",x"20",x"64",x"65"),
  1033 => (x"69",x"74",x"72",x"61"),
  1034 => (x"6e",x"6f",x"69",x"74"),
  1035 => (x"70",x"79",x"74",x"20"),
  1036 => (x"00",x"0d",x"21",x"65"),
  1037 => (x"33",x"54",x"41",x"46"),
  1038 => (x"20",x"20",x"20",x"32"),
  1039 => (x"61",x"65",x"52",x"00"),
  1040 => (x"67",x"6e",x"69",x"64"),
  1041 => (x"52",x"42",x"4d",x"20"),
  1042 => (x"42",x"4d",x"00",x"0a"),
  1043 => (x"75",x"73",x"20",x"52"),
  1044 => (x"73",x"65",x"63",x"63"),
  1045 => (x"6c",x"75",x"66",x"73"),
  1046 => (x"72",x"20",x"79",x"6c"),
  1047 => (x"0a",x"64",x"61",x"65"),
  1048 => (x"54",x"41",x"46",x"00"),
  1049 => (x"20",x"20",x"36",x"31"),
  1050 => (x"41",x"46",x"00",x"20"),
  1051 => (x"20",x"32",x"33",x"54"),
  1052 => (x"50",x"00",x"20",x"20"),
  1053 => (x"69",x"74",x"72",x"61"),
  1054 => (x"6e",x"6f",x"69",x"74"),
  1055 => (x"6e",x"75",x"6f",x"63"),
  1056 => (x"64",x"25",x"20",x"74"),
  1057 => (x"75",x"48",x"00",x"0a"),
  1058 => (x"6e",x"69",x"74",x"6e"),
  1059 => (x"6f",x"66",x"20",x"67"),
  1060 => (x"69",x"66",x"20",x"72"),
  1061 => (x"79",x"73",x"65",x"6c"),
  1062 => (x"6d",x"65",x"74",x"73"),
  1063 => (x"41",x"46",x"00",x"0a"),
  1064 => (x"20",x"32",x"33",x"54"),
  1065 => (x"46",x"00",x"20",x"20"),
  1066 => (x"36",x"31",x"54",x"41"),
  1067 => (x"00",x"20",x"20",x"20"),
  1068 => (x"73",x"75",x"6c",x"43"),
  1069 => (x"20",x"72",x"65",x"74"),
  1070 => (x"65",x"7a",x"69",x"73"),
  1071 => (x"64",x"25",x"20",x"3a"),
  1072 => (x"6c",x"43",x"20",x"2c"),
  1073 => (x"65",x"74",x"73",x"75"),
  1074 => (x"61",x"6d",x"20",x"72"),
  1075 => (x"20",x"2c",x"6b",x"73"),
  1076 => (x"00",x"0a",x"64",x"25"),
  1077 => (x"c4",x"0e",x"5e",x"0e"),
  1078 => (x"29",x"d8",x"49",x"66"),
  1079 => (x"c4",x"99",x"ff",x"c3"),
  1080 => (x"2a",x"c8",x"4a",x"66"),
  1081 => (x"9a",x"c0",x"fc",x"cf"),
  1082 => (x"66",x"c4",x"b1",x"72"),
  1083 => (x"c0",x"32",x"c8",x"4a"),
  1084 => (x"c0",x"c0",x"f0",x"ff"),
  1085 => (x"c4",x"b1",x"72",x"9a"),
  1086 => (x"32",x"d8",x"4a",x"66"),
  1087 => (x"c0",x"c0",x"c0",x"ff"),
  1088 => (x"b1",x"72",x"9a",x"c0"),
  1089 => (x"87",x"c6",x"48",x"71"),
  1090 => (x"4c",x"26",x"4d",x"26"),
  1091 => (x"4f",x"26",x"4b",x"26"),
  1092 => (x"c4",x"0e",x"5e",x"0e"),
  1093 => (x"2a",x"c8",x"4a",x"66"),
  1094 => (x"cf",x"9a",x"ff",x"c3"),
  1095 => (x"c4",x"9a",x"ff",x"ff"),
  1096 => (x"31",x"c8",x"49",x"66"),
  1097 => (x"99",x"c0",x"fc",x"cf"),
  1098 => (x"ff",x"cf",x"b1",x"72"),
  1099 => (x"48",x"71",x"99",x"ff"),
  1100 => (x"0e",x"87",x"db",x"ff"),
  1101 => (x"66",x"c4",x"0e",x"5e"),
  1102 => (x"cf",x"29",x"d0",x"49"),
  1103 => (x"c4",x"99",x"ff",x"ff"),
  1104 => (x"32",x"d0",x"4a",x"66"),
  1105 => (x"9a",x"c0",x"c0",x"f0"),
  1106 => (x"48",x"71",x"b1",x"72"),
  1107 => (x"1e",x"87",x"ff",x"fe"),
  1108 => (x"c0",x"d0",x"1e",x"73"),
  1109 => (x"4b",x"c0",x"c0",x"c0"),
  1110 => (x"87",x"fe",x"0f",x"73"),
  1111 => (x"4d",x"26",x"87",x"c4"),
  1112 => (x"4b",x"26",x"4c",x"26"),
  1113 => (x"c8",x"1e",x"4f",x"26"),
  1114 => (x"df",x"c3",x"49",x"66"),
  1115 => (x"89",x"f7",x"c0",x"99"),
  1116 => (x"03",x"a9",x"b7",x"c0"),
  1117 => (x"e7",x"c0",x"87",x"c3"),
  1118 => (x"48",x"66",x"c4",x"81"),
  1119 => (x"a6",x"c8",x"30",x"c4"),
  1120 => (x"48",x"66",x"c4",x"58"),
  1121 => (x"a6",x"c8",x"b0",x"71"),
  1122 => (x"48",x"66",x"c4",x"58"),
  1123 => (x"0e",x"87",x"d5",x"ff"),
  1124 => (x"0e",x"5c",x"5b",x"5e"),
  1125 => (x"c0",x"c0",x"c0",x"d0"),
  1126 => (x"dd",x"c1",x"4c",x"c0"),
  1127 => (x"c1",x"48",x"bf",x"f0"),
  1128 => (x"f4",x"dd",x"c1",x"80"),
  1129 => (x"66",x"cc",x"97",x"58"),
  1130 => (x"81",x"c0",x"fe",x"49"),
  1131 => (x"a9",x"d3",x"c1",x"b9"),
  1132 => (x"87",x"e1",x"c0",x"05"),
  1133 => (x"48",x"f0",x"dd",x"c1"),
  1134 => (x"dd",x"c1",x"78",x"c0"),
  1135 => (x"78",x"c0",x"48",x"f4"),
  1136 => (x"48",x"fc",x"dd",x"c1"),
  1137 => (x"de",x"c1",x"78",x"c0"),
  1138 => (x"78",x"c0",x"48",x"c0"),
  1139 => (x"c1",x"48",x"c0",x"ff"),
  1140 => (x"ee",x"c7",x"78",x"d3"),
  1141 => (x"f0",x"dd",x"c1",x"87"),
  1142 => (x"a8",x"c1",x"48",x"bf"),
  1143 => (x"87",x"c8",x"c1",x"05"),
  1144 => (x"c1",x"48",x"c0",x"ff"),
  1145 => (x"cc",x"97",x"78",x"f4"),
  1146 => (x"c0",x"fe",x"49",x"66"),
  1147 => (x"1e",x"71",x"b9",x"81"),
  1148 => (x"bf",x"c0",x"de",x"c1"),
  1149 => (x"87",x"ee",x"fd",x"1e"),
  1150 => (x"de",x"c1",x"86",x"c8"),
  1151 => (x"de",x"c1",x"58",x"c4"),
  1152 => (x"c3",x"4a",x"bf",x"c0"),
  1153 => (x"c6",x"06",x"aa",x"b7"),
  1154 => (x"72",x"48",x"ca",x"87"),
  1155 => (x"72",x"4a",x"70",x"88"),
  1156 => (x"71",x"81",x"c1",x"49"),
  1157 => (x"c1",x"30",x"c1",x"48"),
  1158 => (x"72",x"58",x"fc",x"dd"),
  1159 => (x"80",x"f0",x"c0",x"48"),
  1160 => (x"78",x"08",x"c0",x"ff"),
  1161 => (x"87",x"db",x"c6",x"08"),
  1162 => (x"bf",x"c0",x"de",x"c1"),
  1163 => (x"a8",x"b7",x"c9",x"48"),
  1164 => (x"87",x"cf",x"c6",x"01"),
  1165 => (x"bf",x"c0",x"de",x"c1"),
  1166 => (x"a8",x"b7",x"c0",x"48"),
  1167 => (x"87",x"c3",x"c6",x"06"),
  1168 => (x"bf",x"c0",x"de",x"c1"),
  1169 => (x"80",x"f0",x"c0",x"48"),
  1170 => (x"78",x"08",x"c0",x"ff"),
  1171 => (x"f0",x"dd",x"c1",x"08"),
  1172 => (x"b7",x"c3",x"48",x"bf"),
  1173 => (x"87",x"db",x"01",x"a8"),
  1174 => (x"49",x"66",x"cc",x"97"),
  1175 => (x"b9",x"81",x"c0",x"fe"),
  1176 => (x"dd",x"c1",x"1e",x"71"),
  1177 => (x"fb",x"1e",x"bf",x"fc"),
  1178 => (x"86",x"c8",x"87",x"fc"),
  1179 => (x"58",x"c0",x"de",x"c1"),
  1180 => (x"c1",x"87",x"d0",x"c5"),
  1181 => (x"49",x"bf",x"f8",x"dd"),
  1182 => (x"dd",x"c1",x"81",x"c3"),
  1183 => (x"a9",x"b7",x"bf",x"f0"),
  1184 => (x"87",x"e1",x"c0",x"04"),
  1185 => (x"49",x"66",x"cc",x"97"),
  1186 => (x"b9",x"81",x"c0",x"fe"),
  1187 => (x"dd",x"c1",x"1e",x"71"),
  1188 => (x"fb",x"1e",x"bf",x"f4"),
  1189 => (x"86",x"c8",x"87",x"d0"),
  1190 => (x"58",x"f8",x"dd",x"c1"),
  1191 => (x"48",x"c4",x"de",x"c1"),
  1192 => (x"de",x"c4",x"78",x"c1"),
  1193 => (x"c0",x"de",x"c1",x"87"),
  1194 => (x"b7",x"c0",x"48",x"bf"),
  1195 => (x"db",x"c2",x"06",x"a8"),
  1196 => (x"c0",x"de",x"c1",x"87"),
  1197 => (x"b7",x"c3",x"48",x"bf"),
  1198 => (x"cf",x"c2",x"01",x"a8"),
  1199 => (x"fc",x"dd",x"c1",x"87"),
  1200 => (x"31",x"c1",x"49",x"bf"),
  1201 => (x"f0",x"dd",x"c1",x"81"),
  1202 => (x"04",x"a9",x"b7",x"bf"),
  1203 => (x"97",x"87",x"df",x"c1"),
  1204 => (x"fe",x"49",x"66",x"cc"),
  1205 => (x"71",x"b9",x"81",x"c0"),
  1206 => (x"c8",x"de",x"c1",x"1e"),
  1207 => (x"c5",x"fa",x"1e",x"bf"),
  1208 => (x"c1",x"86",x"c8",x"87"),
  1209 => (x"c1",x"58",x"cc",x"de"),
  1210 => (x"49",x"bf",x"c4",x"de"),
  1211 => (x"de",x"c1",x"89",x"c1"),
  1212 => (x"b7",x"c0",x"59",x"c8"),
  1213 => (x"ca",x"c3",x"03",x"a9"),
  1214 => (x"f4",x"dd",x"c1",x"87"),
  1215 => (x"de",x"c1",x"49",x"bf"),
  1216 => (x"51",x"bf",x"97",x"c8"),
  1217 => (x"c1",x"98",x"ff",x"c3"),
  1218 => (x"49",x"bf",x"f4",x"dd"),
  1219 => (x"dd",x"c1",x"81",x"c1"),
  1220 => (x"de",x"c1",x"59",x"f8"),
  1221 => (x"a9",x"b7",x"bf",x"cc"),
  1222 => (x"87",x"c9",x"c0",x"06"),
  1223 => (x"48",x"cc",x"de",x"c1"),
  1224 => (x"bf",x"f4",x"dd",x"c1"),
  1225 => (x"c4",x"de",x"c1",x"78"),
  1226 => (x"c2",x"78",x"c1",x"48"),
  1227 => (x"de",x"c1",x"87",x"d5"),
  1228 => (x"c2",x"05",x"bf",x"c4"),
  1229 => (x"de",x"c1",x"87",x"cd"),
  1230 => (x"c4",x"49",x"bf",x"c8"),
  1231 => (x"cc",x"de",x"c1",x"31"),
  1232 => (x"f4",x"dd",x"c1",x"59"),
  1233 => (x"79",x"97",x"09",x"bf"),
  1234 => (x"87",x"f7",x"c1",x"09"),
  1235 => (x"bf",x"c0",x"de",x"c1"),
  1236 => (x"a8",x"b7",x"c7",x"48"),
  1237 => (x"87",x"de",x"c1",x"04"),
  1238 => (x"f4",x"fe",x"4b",x"c0"),
  1239 => (x"c1",x"78",x"c1",x"48"),
  1240 => (x"1e",x"bf",x"cc",x"de"),
  1241 => (x"d3",x"c1",x"1e",x"74"),
  1242 => (x"f4",x"fe",x"1e",x"e2"),
  1243 => (x"86",x"cc",x"87",x"dc"),
  1244 => (x"5c",x"f8",x"dd",x"c1"),
  1245 => (x"bf",x"f4",x"dd",x"c1"),
  1246 => (x"cc",x"de",x"c1",x"48"),
  1247 => (x"03",x"a8",x"b7",x"bf"),
  1248 => (x"c1",x"87",x"db",x"c0"),
  1249 => (x"bf",x"bf",x"f4",x"dd"),
  1250 => (x"f4",x"dd",x"c1",x"83"),
  1251 => (x"81",x"c4",x"49",x"bf"),
  1252 => (x"59",x"f8",x"dd",x"c1"),
  1253 => (x"bf",x"cc",x"de",x"c1"),
  1254 => (x"ff",x"04",x"a9",x"b7"),
  1255 => (x"1e",x"73",x"87",x"e5"),
  1256 => (x"1e",x"c1",x"d4",x"c1"),
  1257 => (x"87",x"e2",x"f3",x"fe"),
  1258 => (x"c0",x"ff",x"86",x"c8"),
  1259 => (x"78",x"c2",x"c1",x"48"),
  1260 => (x"c0",x"87",x"dc",x"f6"),
  1261 => (x"de",x"c1",x"87",x"cd"),
  1262 => (x"c0",x"48",x"bf",x"c0"),
  1263 => (x"c0",x"ff",x"80",x"f0"),
  1264 => (x"f6",x"08",x"78",x"08"),
  1265 => (x"5e",x"0e",x"87",x"da"),
  1266 => (x"0e",x"5d",x"5c",x"5b"),
  1267 => (x"1e",x"e4",x"d2",x"c1"),
  1268 => (x"87",x"c8",x"f2",x"fe"),
  1269 => (x"c3",x"ff",x"86",x"c4"),
  1270 => (x"98",x"70",x"87",x"c9"),
  1271 => (x"87",x"cf",x"c0",x"02"),
  1272 => (x"87",x"ff",x"d6",x"ff"),
  1273 => (x"c0",x"02",x"98",x"70"),
  1274 => (x"49",x"c1",x"87",x"c5"),
  1275 => (x"c0",x"87",x"c2",x"c0"),
  1276 => (x"c1",x"4d",x"71",x"49"),
  1277 => (x"fe",x"1e",x"fa",x"d2"),
  1278 => (x"c4",x"87",x"e1",x"f1"),
  1279 => (x"cc",x"de",x"c1",x"86"),
  1280 => (x"c0",x"78",x"c0",x"48"),
  1281 => (x"f0",x"fe",x"1e",x"ee"),
  1282 => (x"86",x"c4",x"87",x"f2"),
  1283 => (x"ff",x"c8",x"f4",x"c3"),
  1284 => (x"bf",x"c0",x"ff",x"4a"),
  1285 => (x"c8",x"49",x"74",x"4c"),
  1286 => (x"99",x"71",x"99",x"c0"),
  1287 => (x"87",x"cc",x"c1",x"02"),
  1288 => (x"ff",x"c3",x"4b",x"74"),
  1289 => (x"05",x"ab",x"db",x"9b"),
  1290 => (x"75",x"87",x"f5",x"c0"),
  1291 => (x"e5",x"c0",x"02",x"9d"),
  1292 => (x"c0",x"c0",x"d0",x"87"),
  1293 => (x"c1",x"1e",x"c0",x"c0"),
  1294 => (x"ea",x"1e",x"c8",x"d2"),
  1295 => (x"86",x"c8",x"87",x"c1"),
  1296 => (x"c0",x"02",x"98",x"70"),
  1297 => (x"d1",x"c1",x"87",x"d0"),
  1298 => (x"f0",x"fe",x"1e",x"fc"),
  1299 => (x"86",x"c4",x"87",x"ce"),
  1300 => (x"c0",x"87",x"fc",x"f3"),
  1301 => (x"d2",x"c1",x"87",x"ca"),
  1302 => (x"ef",x"fe",x"1e",x"d4"),
  1303 => (x"86",x"c4",x"87",x"fe"),
  1304 => (x"ea",x"f4",x"1e",x"73"),
  1305 => (x"c3",x"86",x"c4",x"87"),
  1306 => (x"4a",x"c0",x"c9",x"f4"),
  1307 => (x"8a",x"c1",x"49",x"72"),
  1308 => (x"fe",x"05",x"99",x"71"),
  1309 => (x"ca",x"fe",x"87",x"db"),
  1310 => (x"87",x"e2",x"f3",x"87"),
  1311 => (x"74",x"6f",x"6f",x"42"),
  1312 => (x"2e",x"67",x"6e",x"69"),
  1313 => (x"00",x"0a",x"2e",x"2e"),
  1314 => (x"54",x"4f",x"4f",x"42"),
  1315 => (x"20",x"32",x"33",x"38"),
  1316 => (x"00",x"4e",x"49",x"42"),
  1317 => (x"62",x"20",x"44",x"53"),
  1318 => (x"20",x"74",x"6f",x"6f"),
  1319 => (x"6c",x"69",x"61",x"66"),
  1320 => (x"00",x"0a",x"64",x"65"),
  1321 => (x"74",x"69",x"6e",x"49"),
  1322 => (x"69",x"6c",x"61",x"69"),
  1323 => (x"67",x"6e",x"69",x"7a"),
  1324 => (x"20",x"44",x"53",x"20"),
  1325 => (x"64",x"72",x"61",x"63"),
  1326 => (x"53",x"52",x"00",x"0a"),
  1327 => (x"20",x"32",x"33",x"32"),
  1328 => (x"74",x"6f",x"6f",x"62"),
  1329 => (x"70",x"20",x"2d",x"20"),
  1330 => (x"73",x"73",x"65",x"72"),
  1331 => (x"43",x"53",x"45",x"20"),
  1332 => (x"20",x"6f",x"74",x"20"),
  1333 => (x"74",x"6f",x"6f",x"62"),
  1334 => (x"6f",x"72",x"66",x"20"),
  1335 => (x"44",x"53",x"20",x"6d"),
  1336 => (x"68",x"43",x"00",x"2e"),
  1337 => (x"73",x"6b",x"63",x"65"),
  1338 => (x"69",x"6d",x"6d",x"75"),
  1339 => (x"66",x"20",x"67",x"6e"),
  1340 => (x"20",x"6d",x"6f",x"72"),
  1341 => (x"74",x"20",x"64",x"25"),
  1342 => (x"64",x"25",x"20",x"6f"),
  1343 => (x"20",x"2e",x"2e",x"2e"),
  1344 => (x"0a",x"64",x"25",x"00"),
  1345 => (x"0a",x"64",x"25",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
