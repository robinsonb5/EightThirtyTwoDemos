
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"2c",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"29"),
    10 => (x"87",x"fd",x"00",x"4f"),
    11 => (x"c8",x"f4",x"c3",x"4f"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"c8",x"f4",x"c3"),
    14 => (x"48",x"d0",x"d1",x"c1"),
    15 => (x"03",x"89",x"d0",x"89"),
    16 => (x"40",x"40",x"40",x"c0"),
    17 => (x"d0",x"87",x"f6",x"40"),
    18 => (x"50",x"c0",x"05",x"81"),
    19 => (x"f9",x"05",x"89",x"c1"),
    20 => (x"cf",x"d1",x"c1",x"87"),
    21 => (x"cf",x"d1",x"c1",x"4d"),
    22 => (x"02",x"ad",x"74",x"4c"),
    23 => (x"0f",x"24",x"87",x"c4"),
    24 => (x"cd",x"cd",x"87",x"f7"),
    25 => (x"cf",x"d1",x"c1",x"87"),
    26 => (x"cf",x"d1",x"c1",x"4d"),
    27 => (x"02",x"ad",x"74",x"4c"),
    28 => (x"8c",x"c4",x"87",x"c6"),
    29 => (x"87",x"f5",x"0f",x"6c"),
    30 => (x"1e",x"87",x"fd",x"00"),
    31 => (x"c0",x"ff",x"86",x"fc"),
    32 => (x"49",x"bf",x"6e",x"7e"),
    33 => (x"02",x"99",x"c0",x"c4"),
    34 => (x"48",x"6e",x"87",x"f7"),
    35 => (x"48",x"78",x"66",x"c8"),
    36 => (x"4f",x"26",x"8e",x"fc"),
    37 => (x"c1",x"86",x"f0",x"1e"),
    38 => (x"c4",x"7e",x"d0",x"d1"),
    39 => (x"f4",x"c4",x"48",x"a6"),
    40 => (x"c0",x"80",x"c4",x"78"),
    41 => (x"05",x"66",x"d4",x"78"),
    42 => (x"49",x"6e",x"87",x"ce"),
    43 => (x"c4",x"80",x"c1",x"48"),
    44 => (x"f0",x"c0",x"58",x"a6"),
    45 => (x"87",x"c5",x"c1",x"51"),
    46 => (x"71",x"87",x"fc",x"c0"),
    47 => (x"dc",x"1e",x"72",x"1e"),
    48 => (x"e0",x"c0",x"49",x"66"),
    49 => (x"f3",x"c9",x"4a",x"66"),
    50 => (x"26",x"48",x"71",x"87"),
    51 => (x"d0",x"49",x"26",x"4a"),
    52 => (x"66",x"c4",x"58",x"a6"),
    53 => (x"81",x"66",x"cc",x"49"),
    54 => (x"c1",x"48",x"4a",x"6e"),
    55 => (x"58",x"a6",x"c4",x"80"),
    56 => (x"1e",x"71",x"52",x"11"),
    57 => (x"66",x"dc",x"1e",x"72"),
    58 => (x"66",x"e0",x"c0",x"49"),
    59 => (x"87",x"cc",x"c9",x"4a"),
    60 => (x"49",x"26",x"4a",x"26"),
    61 => (x"d4",x"58",x"a6",x"d8"),
    62 => (x"fe",x"fe",x"05",x"66"),
    63 => (x"87",x"e3",x"c0",x"87"),
    64 => (x"1e",x"66",x"e0",x"c0"),
    65 => (x"c1",x"48",x"66",x"c4"),
    66 => (x"58",x"a6",x"c8",x"88"),
    67 => (x"bf",x"97",x"66",x"c4"),
    68 => (x"c0",x"1e",x"71",x"49"),
    69 => (x"c8",x"0f",x"66",x"e4"),
    70 => (x"c8",x"49",x"70",x"86"),
    71 => (x"80",x"c1",x"48",x"66"),
    72 => (x"6e",x"58",x"a6",x"cc"),
    73 => (x"d0",x"d1",x"c1",x"48"),
    74 => (x"d3",x"ff",x"05",x"a8"),
    75 => (x"48",x"66",x"c8",x"87"),
    76 => (x"4f",x"26",x"8e",x"f0"),
    77 => (x"33",x"32",x"31",x"30"),
    78 => (x"37",x"36",x"35",x"34"),
    79 => (x"42",x"41",x"39",x"38"),
    80 => (x"46",x"45",x"44",x"43"),
    81 => (x"86",x"f4",x"1e",x"00"),
    82 => (x"a6",x"c8",x"7e",x"ff"),
    83 => (x"dc",x"78",x"c1",x"48"),
    84 => (x"c1",x"48",x"6e",x"87"),
    85 => (x"58",x"a6",x"c4",x"80"),
    86 => (x"c8",x"1e",x"66",x"d8"),
    87 => (x"66",x"dc",x"1e",x"66"),
    88 => (x"c4",x"86",x"c8",x"0f"),
    89 => (x"c4",x"02",x"a8",x"66"),
    90 => (x"d6",x"48",x"6e",x"87"),
    91 => (x"49",x"66",x"d0",x"87"),
    92 => (x"d4",x"80",x"c1",x"48"),
    93 => (x"48",x"11",x"58",x"a6"),
    94 => (x"c4",x"58",x"a6",x"c8"),
    95 => (x"d0",x"ff",x"05",x"66"),
    96 => (x"f4",x"48",x"6e",x"87"),
    97 => (x"1e",x"4f",x"26",x"8e"),
    98 => (x"7e",x"c0",x"86",x"e8"),
    99 => (x"c0",x"48",x"a6",x"cc"),
   100 => (x"87",x"e6",x"c5",x"78"),
   101 => (x"c5",x"02",x"66",x"cc"),
   102 => (x"a6",x"d4",x"87",x"c1"),
   103 => (x"f4",x"78",x"c0",x"48"),
   104 => (x"cc",x"78",x"c0",x"80"),
   105 => (x"78",x"c0",x"48",x"a6"),
   106 => (x"c0",x"49",x"66",x"c4"),
   107 => (x"c1",x"02",x"a9",x"f0"),
   108 => (x"e3",x"c1",x"87",x"eb"),
   109 => (x"ec",x"c1",x"02",x"a9"),
   110 => (x"a9",x"e4",x"c1",x"87"),
   111 => (x"87",x"e2",x"c0",x"02"),
   112 => (x"02",x"a9",x"ec",x"c1"),
   113 => (x"c1",x"87",x"d6",x"c1"),
   114 => (x"dd",x"02",x"a9",x"f0"),
   115 => (x"a9",x"f3",x"c1",x"87"),
   116 => (x"c1",x"87",x"df",x"02"),
   117 => (x"c9",x"02",x"a9",x"f5"),
   118 => (x"a9",x"f8",x"c1",x"87"),
   119 => (x"c1",x"87",x"cb",x"02"),
   120 => (x"a6",x"d4",x"87",x"eb"),
   121 => (x"c2",x"78",x"ca",x"48"),
   122 => (x"a6",x"d4",x"87",x"d1"),
   123 => (x"c2",x"78",x"d0",x"48"),
   124 => (x"e8",x"c0",x"87",x"c9"),
   125 => (x"e8",x"c0",x"1e",x"66"),
   126 => (x"e8",x"c0",x"1e",x"66"),
   127 => (x"80",x"c4",x"48",x"66"),
   128 => (x"58",x"a6",x"ec",x"c0"),
   129 => (x"49",x"66",x"e8",x"c0"),
   130 => (x"1e",x"69",x"81",x"fc"),
   131 => (x"cc",x"87",x"f6",x"fc"),
   132 => (x"71",x"49",x"70",x"86"),
   133 => (x"c4",x"80",x"6e",x"48"),
   134 => (x"de",x"c1",x"58",x"a6"),
   135 => (x"48",x"a6",x"cc",x"87"),
   136 => (x"d6",x"c1",x"78",x"c1"),
   137 => (x"66",x"e8",x"c0",x"87"),
   138 => (x"66",x"e4",x"c0",x"1e"),
   139 => (x"c0",x"80",x"c4",x"48"),
   140 => (x"c0",x"58",x"a6",x"e8"),
   141 => (x"fc",x"49",x"66",x"e4"),
   142 => (x"c0",x"1e",x"69",x"81"),
   143 => (x"c8",x"0f",x"66",x"ec"),
   144 => (x"6e",x"49",x"70",x"86"),
   145 => (x"c4",x"80",x"c1",x"48"),
   146 => (x"ee",x"c0",x"58",x"a6"),
   147 => (x"48",x"66",x"c4",x"87"),
   148 => (x"02",x"a8",x"e5",x"c0"),
   149 => (x"e8",x"c0",x"87",x"cf"),
   150 => (x"e5",x"c0",x"1e",x"66"),
   151 => (x"66",x"ec",x"c0",x"1e"),
   152 => (x"70",x"86",x"c8",x"0f"),
   153 => (x"66",x"e8",x"c0",x"49"),
   154 => (x"1e",x"66",x"c8",x"1e"),
   155 => (x"0f",x"66",x"ec",x"c0"),
   156 => (x"49",x"70",x"86",x"c8"),
   157 => (x"80",x"c1",x"48",x"6e"),
   158 => (x"d4",x"58",x"a6",x"c4"),
   159 => (x"d8",x"c1",x"02",x"66"),
   160 => (x"66",x"e0",x"c0",x"87"),
   161 => (x"c0",x"80",x"c4",x"48"),
   162 => (x"c0",x"58",x"a6",x"e4"),
   163 => (x"fc",x"49",x"66",x"e0"),
   164 => (x"48",x"a6",x"d0",x"81"),
   165 => (x"66",x"c4",x"78",x"69"),
   166 => (x"a8",x"e4",x"c1",x"48"),
   167 => (x"d0",x"87",x"dc",x"05"),
   168 => (x"b7",x"c0",x"48",x"66"),
   169 => (x"87",x"d3",x"03",x"a8"),
   170 => (x"f7",x"1e",x"ed",x"c0"),
   171 => (x"86",x"c4",x"87",x"cd"),
   172 => (x"66",x"d0",x"49",x"70"),
   173 => (x"88",x"08",x"c0",x"48"),
   174 => (x"c0",x"58",x"a6",x"d4"),
   175 => (x"c0",x"1e",x"66",x"e8"),
   176 => (x"dc",x"1e",x"66",x"e8"),
   177 => (x"66",x"dc",x"1e",x"66"),
   178 => (x"87",x"c8",x"f7",x"1e"),
   179 => (x"a6",x"cc",x"86",x"d0"),
   180 => (x"c8",x"48",x"6e",x"58"),
   181 => (x"a6",x"c4",x"80",x"66"),
   182 => (x"c4",x"87",x"df",x"58"),
   183 => (x"e5",x"c0",x"48",x"66"),
   184 => (x"87",x"c7",x"05",x"a8"),
   185 => (x"c1",x"48",x"a6",x"cc"),
   186 => (x"c0",x"87",x"cf",x"78"),
   187 => (x"c8",x"1e",x"66",x"e8"),
   188 => (x"ec",x"c0",x"1e",x"66"),
   189 => (x"86",x"c8",x"0f",x"66"),
   190 => (x"66",x"dc",x"49",x"70"),
   191 => (x"80",x"c1",x"48",x"49"),
   192 => (x"58",x"a6",x"e0",x"c0"),
   193 => (x"a6",x"c8",x"48",x"11"),
   194 => (x"05",x"66",x"c4",x"58"),
   195 => (x"6e",x"87",x"c5",x"fa"),
   196 => (x"26",x"8e",x"e8",x"48"),
   197 => (x"86",x"f8",x"1e",x"4f"),
   198 => (x"c8",x"48",x"a6",x"d0"),
   199 => (x"1e",x"c0",x"58",x"a6"),
   200 => (x"cc",x"1e",x"fb",x"c1"),
   201 => (x"66",x"d8",x"1e",x"66"),
   202 => (x"87",x"db",x"f9",x"1e"),
   203 => (x"a6",x"c4",x"86",x"d0"),
   204 => (x"48",x"a6",x"c4",x"58"),
   205 => (x"48",x"6e",x"78",x"c0"),
   206 => (x"4f",x"26",x"8e",x"f8"),
   207 => (x"72",x"1e",x"73",x"1e"),
   208 => (x"e7",x"c0",x"02",x"9a"),
   209 => (x"c1",x"48",x"c0",x"87"),
   210 => (x"06",x"a9",x"72",x"4b"),
   211 => (x"82",x"72",x"87",x"d1"),
   212 => (x"73",x"87",x"c9",x"06"),
   213 => (x"01",x"a9",x"72",x"83"),
   214 => (x"87",x"c3",x"87",x"f4"),
   215 => (x"72",x"3a",x"b2",x"c1"),
   216 => (x"73",x"89",x"03",x"a9"),
   217 => (x"2a",x"c1",x"07",x"80"),
   218 => (x"87",x"f3",x"05",x"2b"),
   219 => (x"4f",x"26",x"4b",x"26"),
   220 => (x"c4",x"1e",x"75",x"1e"),
   221 => (x"a1",x"b7",x"71",x"4d"),
   222 => (x"c1",x"b9",x"ff",x"04"),
   223 => (x"07",x"bd",x"c3",x"81"),
   224 => (x"04",x"a2",x"b7",x"72"),
   225 => (x"82",x"c1",x"ba",x"ff"),
   226 => (x"fe",x"07",x"bd",x"c1"),
   227 => (x"2d",x"c1",x"87",x"ee"),
   228 => (x"c1",x"b8",x"ff",x"04"),
   229 => (x"04",x"2d",x"07",x"80"),
   230 => (x"81",x"c1",x"b9",x"ff"),
   231 => (x"26",x"4d",x"26",x"07"),
   232 => (x"1e",x"72",x"1e",x"4f"),
   233 => (x"02",x"11",x"48",x"12"),
   234 => (x"02",x"88",x"87",x"c4"),
   235 => (x"4a",x"26",x"87",x"f6"),
   236 => (x"73",x"1e",x"4f",x"26"),
   237 => (x"75",x"1e",x"74",x"1e"),
   238 => (x"86",x"dc",x"ff",x"1e"),
   239 => (x"48",x"e4",x"d1",x"c1"),
   240 => (x"78",x"e8",x"f1",x"c3"),
   241 => (x"48",x"e0",x"d1",x"c1"),
   242 => (x"78",x"d8",x"f2",x"c3"),
   243 => (x"e8",x"f1",x"c3",x"48"),
   244 => (x"dc",x"f2",x"c3",x"78"),
   245 => (x"c4",x"78",x"c0",x"48"),
   246 => (x"c3",x"78",x"c2",x"80"),
   247 => (x"c0",x"48",x"e4",x"f2"),
   248 => (x"1e",x"71",x"78",x"e8"),
   249 => (x"49",x"e8",x"f2",x"c3"),
   250 => (x"48",x"f8",x"ef",x"c0"),
   251 => (x"41",x"20",x"41",x"20"),
   252 => (x"41",x"20",x"41",x"20"),
   253 => (x"41",x"20",x"41",x"20"),
   254 => (x"51",x"10",x"41",x"20"),
   255 => (x"51",x"10",x"51",x"10"),
   256 => (x"1e",x"71",x"49",x"26"),
   257 => (x"49",x"c8",x"f3",x"c3"),
   258 => (x"48",x"d8",x"f0",x"c0"),
   259 => (x"41",x"20",x"41",x"20"),
   260 => (x"41",x"20",x"41",x"20"),
   261 => (x"41",x"20",x"41",x"20"),
   262 => (x"51",x"10",x"41",x"20"),
   263 => (x"51",x"10",x"51",x"10"),
   264 => (x"ee",x"c1",x"49",x"26"),
   265 => (x"78",x"ca",x"48",x"dc"),
   266 => (x"1e",x"f8",x"f0",x"c0"),
   267 => (x"c4",x"87",x"e6",x"fb"),
   268 => (x"fc",x"f0",x"c0",x"86"),
   269 => (x"87",x"dd",x"fb",x"1e"),
   270 => (x"f1",x"c0",x"86",x"c4"),
   271 => (x"d4",x"fb",x"1e",x"ec"),
   272 => (x"c0",x"86",x"c4",x"87"),
   273 => (x"02",x"bf",x"dc",x"e9"),
   274 => (x"e9",x"c0",x"87",x"d4"),
   275 => (x"c4",x"fb",x"1e",x"e4"),
   276 => (x"c0",x"86",x"c4",x"87"),
   277 => (x"fa",x"1e",x"d0",x"ea"),
   278 => (x"86",x"c4",x"87",x"fb"),
   279 => (x"ea",x"c0",x"87",x"d2"),
   280 => (x"f0",x"fa",x"1e",x"d4"),
   281 => (x"c0",x"86",x"c4",x"87"),
   282 => (x"fa",x"1e",x"c4",x"eb"),
   283 => (x"86",x"c4",x"87",x"e7"),
   284 => (x"bf",x"e0",x"e9",x"c0"),
   285 => (x"f0",x"f1",x"c0",x"1e"),
   286 => (x"87",x"d9",x"fa",x"1e"),
   287 => (x"f1",x"c3",x"86",x"c8"),
   288 => (x"c8",x"ff",x"48",x"d0"),
   289 => (x"a6",x"c8",x"78",x"bf"),
   290 => (x"c0",x"78",x"c1",x"48"),
   291 => (x"48",x"bf",x"e0",x"e9"),
   292 => (x"06",x"a8",x"b7",x"c0"),
   293 => (x"cc",x"87",x"f5",x"c8"),
   294 => (x"a6",x"d4",x"48",x"a6"),
   295 => (x"dc",x"80",x"c8",x"58"),
   296 => (x"a6",x"dc",x"58",x"a6"),
   297 => (x"58",x"a6",x"c8",x"48"),
   298 => (x"48",x"f0",x"d1",x"c1"),
   299 => (x"c1",x"50",x"c1",x"c1"),
   300 => (x"c0",x"48",x"ec",x"d1"),
   301 => (x"f0",x"d1",x"c1",x"78"),
   302 => (x"c1",x"49",x"bf",x"97"),
   303 => (x"c0",x"02",x"a9",x"c1"),
   304 => (x"7e",x"c0",x"87",x"c5"),
   305 => (x"c1",x"87",x"c2",x"c0"),
   306 => (x"ec",x"d1",x"c1",x"7e"),
   307 => (x"b0",x"6e",x"48",x"bf"),
   308 => (x"58",x"f0",x"d1",x"c1"),
   309 => (x"48",x"f4",x"d1",x"c1"),
   310 => (x"dc",x"50",x"c2",x"c1"),
   311 => (x"78",x"c2",x"48",x"a6"),
   312 => (x"78",x"c3",x"80",x"c4"),
   313 => (x"49",x"e8",x"f3",x"c3"),
   314 => (x"48",x"e8",x"eb",x"c0"),
   315 => (x"41",x"20",x"41",x"20"),
   316 => (x"41",x"20",x"41",x"20"),
   317 => (x"41",x"20",x"41",x"20"),
   318 => (x"51",x"10",x"41",x"20"),
   319 => (x"51",x"10",x"51",x"10"),
   320 => (x"c1",x"48",x"a6",x"d4"),
   321 => (x"e8",x"f3",x"c3",x"78"),
   322 => (x"c8",x"f3",x"c3",x"1e"),
   323 => (x"cd",x"fb",x"c0",x"1e"),
   324 => (x"70",x"86",x"c8",x"87"),
   325 => (x"c5",x"c0",x"05",x"98"),
   326 => (x"c0",x"49",x"c1",x"87"),
   327 => (x"49",x"c0",x"87",x"c2"),
   328 => (x"59",x"f0",x"d1",x"c1"),
   329 => (x"c3",x"48",x"66",x"dc"),
   330 => (x"c0",x"03",x"a8",x"b7"),
   331 => (x"66",x"dc",x"87",x"ee"),
   332 => (x"71",x"91",x"c5",x"49"),
   333 => (x"d0",x"88",x"c3",x"48"),
   334 => (x"66",x"d0",x"58",x"a6"),
   335 => (x"c0",x"1e",x"c3",x"1e"),
   336 => (x"c0",x"1e",x"66",x"e4"),
   337 => (x"cc",x"87",x"c4",x"f7"),
   338 => (x"48",x"66",x"dc",x"86"),
   339 => (x"e0",x"c0",x"80",x"c1"),
   340 => (x"66",x"dc",x"58",x"a6"),
   341 => (x"a8",x"b7",x"c3",x"48"),
   342 => (x"87",x"d2",x"ff",x"04"),
   343 => (x"c0",x"1e",x"66",x"cc"),
   344 => (x"c1",x"1e",x"66",x"e0"),
   345 => (x"c1",x"1e",x"c0",x"d5"),
   346 => (x"c0",x"1e",x"f8",x"d1"),
   347 => (x"d0",x"87",x"ee",x"f6"),
   348 => (x"e0",x"d1",x"c1",x"86"),
   349 => (x"d1",x"c1",x"4c",x"bf"),
   350 => (x"4b",x"bf",x"bf",x"e0"),
   351 => (x"49",x"73",x"1e",x"72"),
   352 => (x"bf",x"e0",x"d1",x"c1"),
   353 => (x"a1",x"f0",x"c0",x"48"),
   354 => (x"71",x"41",x"20",x"4a"),
   355 => (x"f8",x"ff",x"05",x"aa"),
   356 => (x"c8",x"4a",x"26",x"87"),
   357 => (x"a4",x"cc",x"7e",x"a4"),
   358 => (x"cc",x"79",x"c5",x"49"),
   359 => (x"7d",x"69",x"4d",x"a3"),
   360 => (x"1e",x"73",x"7b",x"6c"),
   361 => (x"c4",x"87",x"c9",x"d2"),
   362 => (x"49",x"a3",x"c4",x"86"),
   363 => (x"e6",x"c0",x"05",x"69"),
   364 => (x"49",x"a3",x"c8",x"87"),
   365 => (x"1e",x"71",x"7d",x"c6"),
   366 => (x"1e",x"bf",x"66",x"c4"),
   367 => (x"87",x"ef",x"f3",x"c0"),
   368 => (x"d1",x"c1",x"86",x"c8"),
   369 => (x"7b",x"bf",x"bf",x"e0"),
   370 => (x"1e",x"ca",x"1e",x"75"),
   371 => (x"f4",x"c0",x"1e",x"6d"),
   372 => (x"86",x"cc",x"87",x"f9"),
   373 => (x"6c",x"87",x"d9",x"c0"),
   374 => (x"72",x"1e",x"71",x"49"),
   375 => (x"48",x"49",x"74",x"1e"),
   376 => (x"4a",x"a1",x"f0",x"c0"),
   377 => (x"aa",x"71",x"41",x"20"),
   378 => (x"87",x"f8",x"ff",x"05"),
   379 => (x"49",x"26",x"4a",x"26"),
   380 => (x"7e",x"97",x"c1",x"c1"),
   381 => (x"97",x"f4",x"d1",x"c1"),
   382 => (x"c1",x"c1",x"49",x"bf"),
   383 => (x"c1",x"04",x"a9",x"b7"),
   384 => (x"6e",x"97",x"87",x"e1"),
   385 => (x"1e",x"c3",x"c1",x"4b"),
   386 => (x"1e",x"71",x"49",x"73"),
   387 => (x"87",x"ec",x"f6",x"c0"),
   388 => (x"66",x"d4",x"86",x"c8"),
   389 => (x"f9",x"c0",x"05",x"a8"),
   390 => (x"1e",x"66",x"d8",x"87"),
   391 => (x"f2",x"c0",x"1e",x"c0"),
   392 => (x"86",x"c8",x"87",x"cd"),
   393 => (x"f3",x"c3",x"1e",x"71"),
   394 => (x"eb",x"c0",x"49",x"e8"),
   395 => (x"41",x"20",x"48",x"c8"),
   396 => (x"41",x"20",x"41",x"20"),
   397 => (x"41",x"20",x"41",x"20"),
   398 => (x"41",x"20",x"41",x"20"),
   399 => (x"51",x"10",x"51",x"10"),
   400 => (x"49",x"26",x"51",x"10"),
   401 => (x"48",x"a6",x"e0",x"c0"),
   402 => (x"c1",x"78",x"66",x"c8"),
   403 => (x"c8",x"48",x"e8",x"d1"),
   404 => (x"83",x"c1",x"78",x"66"),
   405 => (x"d1",x"c1",x"4a",x"73"),
   406 => (x"49",x"bf",x"97",x"f4"),
   407 => (x"06",x"aa",x"b7",x"71"),
   408 => (x"c0",x"87",x"e2",x"fe"),
   409 => (x"dc",x"48",x"66",x"e0"),
   410 => (x"e4",x"c0",x"90",x"66"),
   411 => (x"1e",x"71",x"58",x"a6"),
   412 => (x"e8",x"c0",x"1e",x"72"),
   413 => (x"66",x"d4",x"49",x"66"),
   414 => (x"87",x"f4",x"f3",x"4a"),
   415 => (x"49",x"26",x"4a",x"26"),
   416 => (x"58",x"a6",x"e0",x"c0"),
   417 => (x"49",x"66",x"e0",x"c0"),
   418 => (x"c7",x"89",x"66",x"cc"),
   419 => (x"dc",x"48",x"71",x"91"),
   420 => (x"e4",x"c0",x"88",x"66"),
   421 => (x"66",x"c4",x"58",x"a6"),
   422 => (x"82",x"ca",x"4a",x"bf"),
   423 => (x"97",x"f0",x"d1",x"c1"),
   424 => (x"c1",x"c1",x"49",x"bf"),
   425 => (x"ce",x"c0",x"05",x"a9"),
   426 => (x"72",x"8a",x"c1",x"87"),
   427 => (x"e8",x"d1",x"c1",x"48"),
   428 => (x"66",x"c4",x"88",x"bf"),
   429 => (x"c8",x"08",x"78",x"08"),
   430 => (x"80",x"c1",x"48",x"66"),
   431 => (x"c8",x"58",x"a6",x"cc"),
   432 => (x"e9",x"c0",x"48",x"66"),
   433 => (x"a8",x"b7",x"bf",x"e0"),
   434 => (x"87",x"dc",x"f7",x"06"),
   435 => (x"48",x"d4",x"f1",x"c3"),
   436 => (x"78",x"bf",x"c8",x"ff"),
   437 => (x"1e",x"e0",x"f2",x"c0"),
   438 => (x"c4",x"87",x"fa",x"f0"),
   439 => (x"f0",x"f2",x"c0",x"86"),
   440 => (x"87",x"f1",x"f0",x"1e"),
   441 => (x"f2",x"c0",x"86",x"c4"),
   442 => (x"e8",x"f0",x"1e",x"f4"),
   443 => (x"c0",x"86",x"c4",x"87"),
   444 => (x"f0",x"1e",x"ec",x"f3"),
   445 => (x"86",x"c4",x"87",x"df"),
   446 => (x"bf",x"e8",x"d1",x"c1"),
   447 => (x"f0",x"f3",x"c0",x"1e"),
   448 => (x"87",x"d1",x"f0",x"1e"),
   449 => (x"1e",x"c5",x"86",x"c8"),
   450 => (x"1e",x"cc",x"f4",x"c0"),
   451 => (x"c8",x"87",x"c6",x"f0"),
   452 => (x"ec",x"d1",x"c1",x"86"),
   453 => (x"f4",x"c0",x"1e",x"bf"),
   454 => (x"f8",x"ef",x"1e",x"e8"),
   455 => (x"c1",x"86",x"c8",x"87"),
   456 => (x"c4",x"f5",x"c0",x"1e"),
   457 => (x"87",x"ed",x"ef",x"1e"),
   458 => (x"d1",x"c1",x"86",x"c8"),
   459 => (x"49",x"bf",x"97",x"f0"),
   460 => (x"f5",x"c0",x"1e",x"71"),
   461 => (x"dc",x"ef",x"1e",x"e0"),
   462 => (x"c1",x"86",x"c8",x"87"),
   463 => (x"f5",x"c0",x"1e",x"c1"),
   464 => (x"d0",x"ef",x"1e",x"fc"),
   465 => (x"c1",x"86",x"c8",x"87"),
   466 => (x"bf",x"97",x"f4",x"d1"),
   467 => (x"c0",x"1e",x"71",x"49"),
   468 => (x"ee",x"1e",x"d8",x"f6"),
   469 => (x"86",x"c8",x"87",x"ff"),
   470 => (x"c0",x"1e",x"c2",x"c1"),
   471 => (x"ee",x"1e",x"f4",x"f6"),
   472 => (x"86",x"c8",x"87",x"f3"),
   473 => (x"bf",x"d8",x"d2",x"c1"),
   474 => (x"d0",x"f7",x"c0",x"1e"),
   475 => (x"87",x"e5",x"ee",x"1e"),
   476 => (x"1e",x"c7",x"86",x"c8"),
   477 => (x"1e",x"ec",x"f7",x"c0"),
   478 => (x"c8",x"87",x"da",x"ee"),
   479 => (x"dc",x"ee",x"c1",x"86"),
   480 => (x"f8",x"c0",x"1e",x"bf"),
   481 => (x"cc",x"ee",x"1e",x"c8"),
   482 => (x"c0",x"86",x"c8",x"87"),
   483 => (x"ee",x"1e",x"e4",x"f8"),
   484 => (x"86",x"c4",x"87",x"c3"),
   485 => (x"1e",x"d0",x"f9",x"c0"),
   486 => (x"c4",x"87",x"fa",x"ed"),
   487 => (x"e0",x"d1",x"c1",x"86"),
   488 => (x"c0",x"1e",x"bf",x"bf"),
   489 => (x"ed",x"1e",x"dc",x"f9"),
   490 => (x"86",x"c8",x"87",x"eb"),
   491 => (x"1e",x"f8",x"f9",x"c0"),
   492 => (x"c4",x"87",x"e2",x"ed"),
   493 => (x"e0",x"d1",x"c1",x"86"),
   494 => (x"81",x"c4",x"49",x"bf"),
   495 => (x"fa",x"c0",x"1e",x"69"),
   496 => (x"d0",x"ed",x"1e",x"ec"),
   497 => (x"c0",x"86",x"c8",x"87"),
   498 => (x"c8",x"fb",x"c0",x"1e"),
   499 => (x"87",x"c5",x"ed",x"1e"),
   500 => (x"d1",x"c1",x"86",x"c8"),
   501 => (x"c8",x"49",x"bf",x"e0"),
   502 => (x"c0",x"1e",x"69",x"81"),
   503 => (x"ec",x"1e",x"e4",x"fb"),
   504 => (x"86",x"c8",x"87",x"f3"),
   505 => (x"fc",x"c0",x"1e",x"c2"),
   506 => (x"e8",x"ec",x"1e",x"c0"),
   507 => (x"c1",x"86",x"c8",x"87"),
   508 => (x"49",x"bf",x"e0",x"d1"),
   509 => (x"1e",x"69",x"81",x"cc"),
   510 => (x"1e",x"dc",x"fc",x"c0"),
   511 => (x"c8",x"87",x"d6",x"ec"),
   512 => (x"c0",x"1e",x"d1",x"86"),
   513 => (x"ec",x"1e",x"f8",x"fc"),
   514 => (x"86",x"c8",x"87",x"cb"),
   515 => (x"bf",x"e0",x"d1",x"c1"),
   516 => (x"71",x"81",x"d0",x"49"),
   517 => (x"d4",x"fd",x"c0",x"1e"),
   518 => (x"87",x"f9",x"eb",x"1e"),
   519 => (x"fd",x"c0",x"86",x"c8"),
   520 => (x"f0",x"eb",x"1e",x"f0"),
   521 => (x"c0",x"86",x"c4",x"87"),
   522 => (x"eb",x"1e",x"e8",x"fe"),
   523 => (x"86",x"c4",x"87",x"e7"),
   524 => (x"bf",x"e4",x"d1",x"c1"),
   525 => (x"fe",x"c0",x"1e",x"bf"),
   526 => (x"d8",x"eb",x"1e",x"fc"),
   527 => (x"c0",x"86",x"c8",x"87"),
   528 => (x"eb",x"1e",x"d8",x"ff"),
   529 => (x"86",x"c4",x"87",x"cf"),
   530 => (x"bf",x"e4",x"d1",x"c1"),
   531 => (x"69",x"81",x"c4",x"49"),
   532 => (x"d8",x"c0",x"c1",x"1e"),
   533 => (x"87",x"fd",x"ea",x"1e"),
   534 => (x"1e",x"c0",x"86",x"c8"),
   535 => (x"1e",x"f4",x"c0",x"c1"),
   536 => (x"c8",x"87",x"f2",x"ea"),
   537 => (x"e4",x"d1",x"c1",x"86"),
   538 => (x"81",x"c8",x"49",x"bf"),
   539 => (x"c1",x"c1",x"1e",x"69"),
   540 => (x"e0",x"ea",x"1e",x"d0"),
   541 => (x"c1",x"86",x"c8",x"87"),
   542 => (x"ec",x"c1",x"c1",x"1e"),
   543 => (x"87",x"d5",x"ea",x"1e"),
   544 => (x"d1",x"c1",x"86",x"c8"),
   545 => (x"cc",x"49",x"bf",x"e4"),
   546 => (x"c1",x"1e",x"69",x"81"),
   547 => (x"ea",x"1e",x"c8",x"c2"),
   548 => (x"86",x"c8",x"87",x"c3"),
   549 => (x"c2",x"c1",x"1e",x"d2"),
   550 => (x"f8",x"e9",x"1e",x"e4"),
   551 => (x"c1",x"86",x"c8",x"87"),
   552 => (x"49",x"bf",x"e4",x"d1"),
   553 => (x"1e",x"71",x"81",x"d0"),
   554 => (x"1e",x"c0",x"c3",x"c1"),
   555 => (x"c8",x"87",x"e6",x"e9"),
   556 => (x"dc",x"c3",x"c1",x"86"),
   557 => (x"87",x"dd",x"e9",x"1e"),
   558 => (x"66",x"dc",x"86",x"c4"),
   559 => (x"d4",x"c4",x"c1",x"1e"),
   560 => (x"87",x"d1",x"e9",x"1e"),
   561 => (x"1e",x"c5",x"86",x"c8"),
   562 => (x"1e",x"f0",x"c4",x"c1"),
   563 => (x"c8",x"87",x"c6",x"e9"),
   564 => (x"66",x"e0",x"c0",x"86"),
   565 => (x"cc",x"c5",x"c1",x"1e"),
   566 => (x"87",x"f9",x"e8",x"1e"),
   567 => (x"1e",x"cd",x"86",x"c8"),
   568 => (x"1e",x"e8",x"c5",x"c1"),
   569 => (x"c8",x"87",x"ee",x"e8"),
   570 => (x"1e",x"66",x"cc",x"86"),
   571 => (x"1e",x"c4",x"c6",x"c1"),
   572 => (x"c8",x"87",x"e2",x"e8"),
   573 => (x"c1",x"1e",x"c7",x"86"),
   574 => (x"e8",x"1e",x"e0",x"c6"),
   575 => (x"86",x"c8",x"87",x"d7"),
   576 => (x"c1",x"1e",x"66",x"d4"),
   577 => (x"e8",x"1e",x"fc",x"c6"),
   578 => (x"86",x"c8",x"87",x"cb"),
   579 => (x"c7",x"c1",x"1e",x"c1"),
   580 => (x"c0",x"e8",x"1e",x"d8"),
   581 => (x"c3",x"86",x"c8",x"87"),
   582 => (x"c1",x"1e",x"c8",x"f3"),
   583 => (x"e7",x"1e",x"f4",x"c7"),
   584 => (x"86",x"c8",x"87",x"f3"),
   585 => (x"1e",x"d0",x"c8",x"c1"),
   586 => (x"c4",x"87",x"ea",x"e7"),
   587 => (x"e8",x"f3",x"c3",x"86"),
   588 => (x"c8",x"c9",x"c1",x"1e"),
   589 => (x"87",x"dd",x"e7",x"1e"),
   590 => (x"c9",x"c1",x"86",x"c8"),
   591 => (x"d4",x"e7",x"1e",x"e4"),
   592 => (x"c1",x"86",x"c4",x"87"),
   593 => (x"e7",x"1e",x"dc",x"ca"),
   594 => (x"86",x"c4",x"87",x"cb"),
   595 => (x"bf",x"d4",x"f1",x"c3"),
   596 => (x"d0",x"f1",x"c3",x"49"),
   597 => (x"f1",x"c3",x"89",x"bf"),
   598 => (x"1e",x"71",x"59",x"dc"),
   599 => (x"1e",x"e0",x"ca",x"c1"),
   600 => (x"c8",x"87",x"f2",x"e6"),
   601 => (x"d8",x"f1",x"c3",x"86"),
   602 => (x"f8",x"c1",x"48",x"bf"),
   603 => (x"c0",x"03",x"a8",x"b7"),
   604 => (x"ec",x"c0",x"87",x"db"),
   605 => (x"dc",x"e6",x"1e",x"c8"),
   606 => (x"c0",x"86",x"c4",x"87"),
   607 => (x"e6",x"1e",x"c0",x"ed"),
   608 => (x"86",x"c4",x"87",x"d3"),
   609 => (x"1e",x"e0",x"ed",x"c0"),
   610 => (x"c4",x"87",x"ca",x"e6"),
   611 => (x"d8",x"f1",x"c3",x"86"),
   612 => (x"4a",x"71",x"49",x"bf"),
   613 => (x"71",x"92",x"e8",x"cf"),
   614 => (x"72",x"1e",x"72",x"1e"),
   615 => (x"e0",x"e9",x"c0",x"49"),
   616 => (x"cb",x"e7",x"4a",x"bf"),
   617 => (x"26",x"4a",x"26",x"87"),
   618 => (x"e0",x"f1",x"c3",x"49"),
   619 => (x"e0",x"e9",x"c0",x"58"),
   620 => (x"4b",x"72",x"4a",x"bf"),
   621 => (x"71",x"93",x"e8",x"cf"),
   622 => (x"73",x"1e",x"72",x"1e"),
   623 => (x"ef",x"e6",x"4a",x"09"),
   624 => (x"26",x"4a",x"26",x"87"),
   625 => (x"e4",x"f1",x"c3",x"49"),
   626 => (x"92",x"f9",x"c8",x"58"),
   627 => (x"1e",x"72",x"1e",x"71"),
   628 => (x"e6",x"4a",x"09",x"72"),
   629 => (x"4a",x"26",x"87",x"da"),
   630 => (x"f1",x"c3",x"49",x"26"),
   631 => (x"ed",x"c0",x"58",x"e8"),
   632 => (x"f0",x"e4",x"1e",x"e4"),
   633 => (x"c3",x"86",x"c4",x"87"),
   634 => (x"1e",x"bf",x"dc",x"f1"),
   635 => (x"1e",x"d4",x"ee",x"c0"),
   636 => (x"c8",x"87",x"e2",x"e4"),
   637 => (x"dc",x"ee",x"c0",x"86"),
   638 => (x"87",x"d9",x"e4",x"1e"),
   639 => (x"f1",x"c3",x"86",x"c4"),
   640 => (x"c0",x"1e",x"bf",x"e0"),
   641 => (x"e4",x"1e",x"cc",x"ef"),
   642 => (x"86",x"c8",x"87",x"cb"),
   643 => (x"bf",x"e4",x"f1",x"c3"),
   644 => (x"d4",x"ef",x"c0",x"1e"),
   645 => (x"87",x"fd",x"e3",x"1e"),
   646 => (x"ef",x"c0",x"86",x"c8"),
   647 => (x"f4",x"e3",x"1e",x"f4"),
   648 => (x"c0",x"86",x"c4",x"87"),
   649 => (x"8e",x"dc",x"ff",x"48"),
   650 => (x"4c",x"26",x"4d",x"26"),
   651 => (x"4f",x"26",x"4b",x"26"),
   652 => (x"e0",x"d1",x"c1",x"1e"),
   653 => (x"87",x"c9",x"02",x"bf"),
   654 => (x"c1",x"48",x"66",x"c4"),
   655 => (x"bf",x"bf",x"e0",x"d1"),
   656 => (x"e0",x"d1",x"c1",x"78"),
   657 => (x"81",x"cc",x"49",x"bf"),
   658 => (x"d1",x"c1",x"1e",x"71"),
   659 => (x"ca",x"1e",x"bf",x"e8"),
   660 => (x"f6",x"e2",x"c0",x"1e"),
   661 => (x"26",x"86",x"cc",x"87"),
   662 => (x"00",x"00",x"00",x"4f"),
   663 => (x"00",x"00",x"00",x"00"),
   664 => (x"00",x"00",x"61",x"a8"),
   665 => (x"67",x"6f",x"72",x"50"),
   666 => (x"20",x"6d",x"61",x"72"),
   667 => (x"70",x"6d",x"6f",x"63"),
   668 => (x"64",x"65",x"6c",x"69"),
   669 => (x"74",x"69",x"77",x"20"),
   670 => (x"72",x"27",x"20",x"68"),
   671 => (x"73",x"69",x"67",x"65"),
   672 => (x"27",x"72",x"65",x"74"),
   673 => (x"74",x"74",x"61",x"20"),
   674 => (x"75",x"62",x"69",x"72"),
   675 => (x"00",x"0a",x"65",x"74"),
   676 => (x"00",x"00",x"00",x"0a"),
   677 => (x"67",x"6f",x"72",x"50"),
   678 => (x"20",x"6d",x"61",x"72"),
   679 => (x"70",x"6d",x"6f",x"63"),
   680 => (x"64",x"65",x"6c",x"69"),
   681 => (x"74",x"69",x"77",x"20"),
   682 => (x"74",x"75",x"6f",x"68"),
   683 => (x"65",x"72",x"27",x"20"),
   684 => (x"74",x"73",x"69",x"67"),
   685 => (x"20",x"27",x"72",x"65"),
   686 => (x"72",x"74",x"74",x"61"),
   687 => (x"74",x"75",x"62",x"69"),
   688 => (x"00",x"00",x"0a",x"65"),
   689 => (x"00",x"00",x"00",x"0a"),
   690 => (x"59",x"52",x"48",x"44"),
   691 => (x"4e",x"4f",x"54",x"53"),
   692 => (x"52",x"50",x"20",x"45"),
   693 => (x"41",x"52",x"47",x"4f"),
   694 => (x"33",x"20",x"2c",x"4d"),
   695 => (x"20",x"44",x"52",x"27"),
   696 => (x"49",x"52",x"54",x"53"),
   697 => (x"00",x"00",x"47",x"4e"),
   698 => (x"59",x"52",x"48",x"44"),
   699 => (x"4e",x"4f",x"54",x"53"),
   700 => (x"52",x"50",x"20",x"45"),
   701 => (x"41",x"52",x"47",x"4f"),
   702 => (x"32",x"20",x"2c",x"4d"),
   703 => (x"20",x"44",x"4e",x"27"),
   704 => (x"49",x"52",x"54",x"53"),
   705 => (x"00",x"00",x"47",x"4e"),
   706 => (x"73",x"61",x"65",x"4d"),
   707 => (x"64",x"65",x"72",x"75"),
   708 => (x"6d",x"69",x"74",x"20"),
   709 => (x"6f",x"74",x"20",x"65"),
   710 => (x"6d",x"73",x"20",x"6f"),
   711 => (x"20",x"6c",x"6c",x"61"),
   712 => (x"6f",x"20",x"6f",x"74"),
   713 => (x"69",x"61",x"74",x"62"),
   714 => (x"65",x"6d",x"20",x"6e"),
   715 => (x"6e",x"69",x"6e",x"61"),
   716 => (x"6c",x"75",x"66",x"67"),
   717 => (x"73",x"65",x"72",x"20"),
   718 => (x"73",x"74",x"6c",x"75"),
   719 => (x"00",x"00",x"00",x"0a"),
   720 => (x"61",x"65",x"6c",x"50"),
   721 => (x"69",x"20",x"65",x"73"),
   722 => (x"65",x"72",x"63",x"6e"),
   723 => (x"20",x"65",x"73",x"61"),
   724 => (x"62",x"6d",x"75",x"6e"),
   725 => (x"6f",x"20",x"72",x"65"),
   726 => (x"75",x"72",x"20",x"66"),
   727 => (x"00",x"0a",x"73",x"6e"),
   728 => (x"00",x"00",x"00",x"0a"),
   729 => (x"72",x"63",x"69",x"4d"),
   730 => (x"63",x"65",x"73",x"6f"),
   731 => (x"73",x"64",x"6e",x"6f"),
   732 => (x"72",x"6f",x"66",x"20"),
   733 => (x"65",x"6e",x"6f",x"20"),
   734 => (x"6e",x"75",x"72",x"20"),
   735 => (x"72",x"68",x"74",x"20"),
   736 => (x"68",x"67",x"75",x"6f"),
   737 => (x"72",x"68",x"44",x"20"),
   738 => (x"6f",x"74",x"73",x"79"),
   739 => (x"20",x"3a",x"65",x"6e"),
   740 => (x"00",x"00",x"00",x"00"),
   741 => (x"0a",x"20",x"64",x"25"),
   742 => (x"00",x"00",x"00",x"00"),
   743 => (x"79",x"72",x"68",x"44"),
   744 => (x"6e",x"6f",x"74",x"73"),
   745 => (x"70",x"20",x"73",x"65"),
   746 => (x"53",x"20",x"72",x"65"),
   747 => (x"6e",x"6f",x"63",x"65"),
   748 => (x"20",x"20",x"3a",x"64"),
   749 => (x"20",x"20",x"20",x"20"),
   750 => (x"20",x"20",x"20",x"20"),
   751 => (x"20",x"20",x"20",x"20"),
   752 => (x"20",x"20",x"20",x"20"),
   753 => (x"20",x"20",x"20",x"20"),
   754 => (x"00",x"00",x"00",x"00"),
   755 => (x"0a",x"20",x"64",x"25"),
   756 => (x"00",x"00",x"00",x"00"),
   757 => (x"20",x"58",x"41",x"56"),
   758 => (x"53",x"50",x"49",x"4d"),
   759 => (x"74",x"61",x"72",x"20"),
   760 => (x"20",x"67",x"6e",x"69"),
   761 => (x"30",x"31",x"20",x"2a"),
   762 => (x"3d",x"20",x"30",x"30"),
   763 => (x"20",x"64",x"25",x"20"),
   764 => (x"00",x"00",x"00",x"0a"),
   765 => (x"00",x"00",x"00",x"0a"),
   766 => (x"59",x"52",x"48",x"44"),
   767 => (x"4e",x"4f",x"54",x"53"),
   768 => (x"52",x"50",x"20",x"45"),
   769 => (x"41",x"52",x"47",x"4f"),
   770 => (x"53",x"20",x"2c",x"4d"),
   771 => (x"20",x"45",x"4d",x"4f"),
   772 => (x"49",x"52",x"54",x"53"),
   773 => (x"00",x"00",x"47",x"4e"),
   774 => (x"59",x"52",x"48",x"44"),
   775 => (x"4e",x"4f",x"54",x"53"),
   776 => (x"52",x"50",x"20",x"45"),
   777 => (x"41",x"52",x"47",x"4f"),
   778 => (x"31",x"20",x"2c",x"4d"),
   779 => (x"20",x"54",x"53",x"27"),
   780 => (x"49",x"52",x"54",x"53"),
   781 => (x"00",x"00",x"47",x"4e"),
   782 => (x"00",x"00",x"00",x"0a"),
   783 => (x"79",x"72",x"68",x"44"),
   784 => (x"6e",x"6f",x"74",x"73"),
   785 => (x"65",x"42",x"20",x"65"),
   786 => (x"6d",x"68",x"63",x"6e"),
   787 => (x"2c",x"6b",x"72",x"61"),
   788 => (x"72",x"65",x"56",x"20"),
   789 => (x"6e",x"6f",x"69",x"73"),
   790 => (x"31",x"2e",x"32",x"20"),
   791 => (x"61",x"4c",x"28",x"20"),
   792 => (x"61",x"75",x"67",x"6e"),
   793 => (x"20",x"3a",x"65",x"67"),
   794 => (x"00",x"0a",x"29",x"43"),
   795 => (x"00",x"00",x"00",x"0a"),
   796 => (x"63",x"65",x"78",x"45"),
   797 => (x"6f",x"69",x"74",x"75"),
   798 => (x"74",x"73",x"20",x"6e"),
   799 => (x"73",x"74",x"72",x"61"),
   800 => (x"64",x"25",x"20",x"2c"),
   801 => (x"6e",x"75",x"72",x"20"),
   802 => (x"68",x"74",x"20",x"73"),
   803 => (x"67",x"75",x"6f",x"72"),
   804 => (x"68",x"44",x"20",x"68"),
   805 => (x"74",x"73",x"79",x"72"),
   806 => (x"0a",x"65",x"6e",x"6f"),
   807 => (x"00",x"00",x"00",x"00"),
   808 => (x"63",x"65",x"78",x"45"),
   809 => (x"6f",x"69",x"74",x"75"),
   810 => (x"6e",x"65",x"20",x"6e"),
   811 => (x"00",x"0a",x"73",x"64"),
   812 => (x"00",x"00",x"00",x"0a"),
   813 => (x"61",x"6e",x"69",x"46"),
   814 => (x"61",x"76",x"20",x"6c"),
   815 => (x"73",x"65",x"75",x"6c"),
   816 => (x"20",x"66",x"6f",x"20"),
   817 => (x"20",x"65",x"68",x"74"),
   818 => (x"69",x"72",x"61",x"76"),
   819 => (x"65",x"6c",x"62",x"61"),
   820 => (x"73",x"75",x"20",x"73"),
   821 => (x"69",x"20",x"64",x"65"),
   822 => (x"68",x"74",x"20",x"6e"),
   823 => (x"65",x"62",x"20",x"65"),
   824 => (x"6d",x"68",x"63",x"6e"),
   825 => (x"3a",x"6b",x"72",x"61"),
   826 => (x"00",x"00",x"00",x"0a"),
   827 => (x"00",x"00",x"00",x"0a"),
   828 => (x"5f",x"74",x"6e",x"49"),
   829 => (x"62",x"6f",x"6c",x"47"),
   830 => (x"20",x"20",x"20",x"3a"),
   831 => (x"20",x"20",x"20",x"20"),
   832 => (x"20",x"20",x"20",x"20"),
   833 => (x"0a",x"64",x"25",x"20"),
   834 => (x"00",x"00",x"00",x"00"),
   835 => (x"20",x"20",x"20",x"20"),
   836 => (x"20",x"20",x"20",x"20"),
   837 => (x"75",x"6f",x"68",x"73"),
   838 => (x"62",x"20",x"64",x"6c"),
   839 => (x"20",x"20",x"3a",x"65"),
   840 => (x"0a",x"64",x"25",x"20"),
   841 => (x"00",x"00",x"00",x"00"),
   842 => (x"6c",x"6f",x"6f",x"42"),
   843 => (x"6f",x"6c",x"47",x"5f"),
   844 => (x"20",x"20",x"3a",x"62"),
   845 => (x"20",x"20",x"20",x"20"),
   846 => (x"20",x"20",x"20",x"20"),
   847 => (x"0a",x"64",x"25",x"20"),
   848 => (x"00",x"00",x"00",x"00"),
   849 => (x"20",x"20",x"20",x"20"),
   850 => (x"20",x"20",x"20",x"20"),
   851 => (x"75",x"6f",x"68",x"73"),
   852 => (x"62",x"20",x"64",x"6c"),
   853 => (x"20",x"20",x"3a",x"65"),
   854 => (x"0a",x"64",x"25",x"20"),
   855 => (x"00",x"00",x"00",x"00"),
   856 => (x"31",x"5f",x"68",x"43"),
   857 => (x"6f",x"6c",x"47",x"5f"),
   858 => (x"20",x"20",x"3a",x"62"),
   859 => (x"20",x"20",x"20",x"20"),
   860 => (x"20",x"20",x"20",x"20"),
   861 => (x"0a",x"63",x"25",x"20"),
   862 => (x"00",x"00",x"00",x"00"),
   863 => (x"20",x"20",x"20",x"20"),
   864 => (x"20",x"20",x"20",x"20"),
   865 => (x"75",x"6f",x"68",x"73"),
   866 => (x"62",x"20",x"64",x"6c"),
   867 => (x"20",x"20",x"3a",x"65"),
   868 => (x"0a",x"63",x"25",x"20"),
   869 => (x"00",x"00",x"00",x"00"),
   870 => (x"32",x"5f",x"68",x"43"),
   871 => (x"6f",x"6c",x"47",x"5f"),
   872 => (x"20",x"20",x"3a",x"62"),
   873 => (x"20",x"20",x"20",x"20"),
   874 => (x"20",x"20",x"20",x"20"),
   875 => (x"0a",x"63",x"25",x"20"),
   876 => (x"00",x"00",x"00",x"00"),
   877 => (x"20",x"20",x"20",x"20"),
   878 => (x"20",x"20",x"20",x"20"),
   879 => (x"75",x"6f",x"68",x"73"),
   880 => (x"62",x"20",x"64",x"6c"),
   881 => (x"20",x"20",x"3a",x"65"),
   882 => (x"0a",x"63",x"25",x"20"),
   883 => (x"00",x"00",x"00",x"00"),
   884 => (x"5f",x"72",x"72",x"41"),
   885 => (x"6c",x"47",x"5f",x"31"),
   886 => (x"38",x"5b",x"62",x"6f"),
   887 => (x"20",x"20",x"3a",x"5d"),
   888 => (x"20",x"20",x"20",x"20"),
   889 => (x"0a",x"64",x"25",x"20"),
   890 => (x"00",x"00",x"00",x"00"),
   891 => (x"20",x"20",x"20",x"20"),
   892 => (x"20",x"20",x"20",x"20"),
   893 => (x"75",x"6f",x"68",x"73"),
   894 => (x"62",x"20",x"64",x"6c"),
   895 => (x"20",x"20",x"3a",x"65"),
   896 => (x"0a",x"64",x"25",x"20"),
   897 => (x"00",x"00",x"00",x"00"),
   898 => (x"5f",x"72",x"72",x"41"),
   899 => (x"6c",x"47",x"5f",x"32"),
   900 => (x"38",x"5b",x"62",x"6f"),
   901 => (x"5d",x"37",x"5b",x"5d"),
   902 => (x"20",x"20",x"20",x"3a"),
   903 => (x"0a",x"64",x"25",x"20"),
   904 => (x"00",x"00",x"00",x"00"),
   905 => (x"20",x"20",x"20",x"20"),
   906 => (x"20",x"20",x"20",x"20"),
   907 => (x"75",x"6f",x"68",x"73"),
   908 => (x"62",x"20",x"64",x"6c"),
   909 => (x"20",x"20",x"3a",x"65"),
   910 => (x"6d",x"75",x"4e",x"20"),
   911 => (x"5f",x"72",x"65",x"62"),
   912 => (x"52",x"5f",x"66",x"4f"),
   913 => (x"20",x"73",x"6e",x"75"),
   914 => (x"30",x"31",x"20",x"2b"),
   915 => (x"00",x"00",x"00",x"0a"),
   916 => (x"5f",x"72",x"74",x"50"),
   917 => (x"62",x"6f",x"6c",x"47"),
   918 => (x"00",x"0a",x"3e",x"2d"),
   919 => (x"74",x"50",x"20",x"20"),
   920 => (x"6f",x"43",x"5f",x"72"),
   921 => (x"20",x"3a",x"70",x"6d"),
   922 => (x"20",x"20",x"20",x"20"),
   923 => (x"20",x"20",x"20",x"20"),
   924 => (x"0a",x"64",x"25",x"20"),
   925 => (x"00",x"00",x"00",x"00"),
   926 => (x"20",x"20",x"20",x"20"),
   927 => (x"20",x"20",x"20",x"20"),
   928 => (x"75",x"6f",x"68",x"73"),
   929 => (x"62",x"20",x"64",x"6c"),
   930 => (x"20",x"20",x"3a",x"65"),
   931 => (x"6d",x"69",x"28",x"20"),
   932 => (x"6d",x"65",x"6c",x"70"),
   933 => (x"61",x"74",x"6e",x"65"),
   934 => (x"6e",x"6f",x"69",x"74"),
   935 => (x"70",x"65",x"64",x"2d"),
   936 => (x"65",x"64",x"6e",x"65"),
   937 => (x"0a",x"29",x"74",x"6e"),
   938 => (x"00",x"00",x"00",x"00"),
   939 => (x"69",x"44",x"20",x"20"),
   940 => (x"3a",x"72",x"63",x"73"),
   941 => (x"20",x"20",x"20",x"20"),
   942 => (x"20",x"20",x"20",x"20"),
   943 => (x"20",x"20",x"20",x"20"),
   944 => (x"0a",x"64",x"25",x"20"),
   945 => (x"00",x"00",x"00",x"00"),
   946 => (x"20",x"20",x"20",x"20"),
   947 => (x"20",x"20",x"20",x"20"),
   948 => (x"75",x"6f",x"68",x"73"),
   949 => (x"62",x"20",x"64",x"6c"),
   950 => (x"20",x"20",x"3a",x"65"),
   951 => (x"0a",x"64",x"25",x"20"),
   952 => (x"00",x"00",x"00",x"00"),
   953 => (x"6e",x"45",x"20",x"20"),
   954 => (x"43",x"5f",x"6d",x"75"),
   955 => (x"3a",x"70",x"6d",x"6f"),
   956 => (x"20",x"20",x"20",x"20"),
   957 => (x"20",x"20",x"20",x"20"),
   958 => (x"0a",x"64",x"25",x"20"),
   959 => (x"00",x"00",x"00",x"00"),
   960 => (x"20",x"20",x"20",x"20"),
   961 => (x"20",x"20",x"20",x"20"),
   962 => (x"75",x"6f",x"68",x"73"),
   963 => (x"62",x"20",x"64",x"6c"),
   964 => (x"20",x"20",x"3a",x"65"),
   965 => (x"0a",x"64",x"25",x"20"),
   966 => (x"00",x"00",x"00",x"00"),
   967 => (x"6e",x"49",x"20",x"20"),
   968 => (x"6f",x"43",x"5f",x"74"),
   969 => (x"20",x"3a",x"70",x"6d"),
   970 => (x"20",x"20",x"20",x"20"),
   971 => (x"20",x"20",x"20",x"20"),
   972 => (x"0a",x"64",x"25",x"20"),
   973 => (x"00",x"00",x"00",x"00"),
   974 => (x"20",x"20",x"20",x"20"),
   975 => (x"20",x"20",x"20",x"20"),
   976 => (x"75",x"6f",x"68",x"73"),
   977 => (x"62",x"20",x"64",x"6c"),
   978 => (x"20",x"20",x"3a",x"65"),
   979 => (x"0a",x"64",x"25",x"20"),
   980 => (x"00",x"00",x"00",x"00"),
   981 => (x"74",x"53",x"20",x"20"),
   982 => (x"6f",x"43",x"5f",x"72"),
   983 => (x"20",x"3a",x"70",x"6d"),
   984 => (x"20",x"20",x"20",x"20"),
   985 => (x"20",x"20",x"20",x"20"),
   986 => (x"0a",x"73",x"25",x"20"),
   987 => (x"00",x"00",x"00",x"00"),
   988 => (x"20",x"20",x"20",x"20"),
   989 => (x"20",x"20",x"20",x"20"),
   990 => (x"75",x"6f",x"68",x"73"),
   991 => (x"62",x"20",x"64",x"6c"),
   992 => (x"20",x"20",x"3a",x"65"),
   993 => (x"52",x"48",x"44",x"20"),
   994 => (x"4f",x"54",x"53",x"59"),
   995 => (x"50",x"20",x"45",x"4e"),
   996 => (x"52",x"47",x"4f",x"52"),
   997 => (x"20",x"2c",x"4d",x"41"),
   998 => (x"45",x"4d",x"4f",x"53"),
   999 => (x"52",x"54",x"53",x"20"),
  1000 => (x"0a",x"47",x"4e",x"49"),
  1001 => (x"00",x"00",x"00",x"00"),
  1002 => (x"74",x"78",x"65",x"4e"),
  1003 => (x"72",x"74",x"50",x"5f"),
  1004 => (x"6f",x"6c",x"47",x"5f"),
  1005 => (x"0a",x"3e",x"2d",x"62"),
  1006 => (x"00",x"00",x"00",x"00"),
  1007 => (x"74",x"50",x"20",x"20"),
  1008 => (x"6f",x"43",x"5f",x"72"),
  1009 => (x"20",x"3a",x"70",x"6d"),
  1010 => (x"20",x"20",x"20",x"20"),
  1011 => (x"20",x"20",x"20",x"20"),
  1012 => (x"0a",x"64",x"25",x"20"),
  1013 => (x"00",x"00",x"00",x"00"),
  1014 => (x"20",x"20",x"20",x"20"),
  1015 => (x"20",x"20",x"20",x"20"),
  1016 => (x"75",x"6f",x"68",x"73"),
  1017 => (x"62",x"20",x"64",x"6c"),
  1018 => (x"20",x"20",x"3a",x"65"),
  1019 => (x"6d",x"69",x"28",x"20"),
  1020 => (x"6d",x"65",x"6c",x"70"),
  1021 => (x"61",x"74",x"6e",x"65"),
  1022 => (x"6e",x"6f",x"69",x"74"),
  1023 => (x"70",x"65",x"64",x"2d"),
  1024 => (x"65",x"64",x"6e",x"65"),
  1025 => (x"2c",x"29",x"74",x"6e"),
  1026 => (x"6d",x"61",x"73",x"20"),
  1027 => (x"73",x"61",x"20",x"65"),
  1028 => (x"6f",x"62",x"61",x"20"),
  1029 => (x"00",x"0a",x"65",x"76"),
  1030 => (x"69",x"44",x"20",x"20"),
  1031 => (x"3a",x"72",x"63",x"73"),
  1032 => (x"20",x"20",x"20",x"20"),
  1033 => (x"20",x"20",x"20",x"20"),
  1034 => (x"20",x"20",x"20",x"20"),
  1035 => (x"0a",x"64",x"25",x"20"),
  1036 => (x"00",x"00",x"00",x"00"),
  1037 => (x"20",x"20",x"20",x"20"),
  1038 => (x"20",x"20",x"20",x"20"),
  1039 => (x"75",x"6f",x"68",x"73"),
  1040 => (x"62",x"20",x"64",x"6c"),
  1041 => (x"20",x"20",x"3a",x"65"),
  1042 => (x"0a",x"64",x"25",x"20"),
  1043 => (x"00",x"00",x"00",x"00"),
  1044 => (x"6e",x"45",x"20",x"20"),
  1045 => (x"43",x"5f",x"6d",x"75"),
  1046 => (x"3a",x"70",x"6d",x"6f"),
  1047 => (x"20",x"20",x"20",x"20"),
  1048 => (x"20",x"20",x"20",x"20"),
  1049 => (x"0a",x"64",x"25",x"20"),
  1050 => (x"00",x"00",x"00",x"00"),
  1051 => (x"20",x"20",x"20",x"20"),
  1052 => (x"20",x"20",x"20",x"20"),
  1053 => (x"75",x"6f",x"68",x"73"),
  1054 => (x"62",x"20",x"64",x"6c"),
  1055 => (x"20",x"20",x"3a",x"65"),
  1056 => (x"0a",x"64",x"25",x"20"),
  1057 => (x"00",x"00",x"00",x"00"),
  1058 => (x"6e",x"49",x"20",x"20"),
  1059 => (x"6f",x"43",x"5f",x"74"),
  1060 => (x"20",x"3a",x"70",x"6d"),
  1061 => (x"20",x"20",x"20",x"20"),
  1062 => (x"20",x"20",x"20",x"20"),
  1063 => (x"0a",x"64",x"25",x"20"),
  1064 => (x"00",x"00",x"00",x"00"),
  1065 => (x"20",x"20",x"20",x"20"),
  1066 => (x"20",x"20",x"20",x"20"),
  1067 => (x"75",x"6f",x"68",x"73"),
  1068 => (x"62",x"20",x"64",x"6c"),
  1069 => (x"20",x"20",x"3a",x"65"),
  1070 => (x"0a",x"64",x"25",x"20"),
  1071 => (x"00",x"00",x"00",x"00"),
  1072 => (x"74",x"53",x"20",x"20"),
  1073 => (x"6f",x"43",x"5f",x"72"),
  1074 => (x"20",x"3a",x"70",x"6d"),
  1075 => (x"20",x"20",x"20",x"20"),
  1076 => (x"20",x"20",x"20",x"20"),
  1077 => (x"0a",x"73",x"25",x"20"),
  1078 => (x"00",x"00",x"00",x"00"),
  1079 => (x"20",x"20",x"20",x"20"),
  1080 => (x"20",x"20",x"20",x"20"),
  1081 => (x"75",x"6f",x"68",x"73"),
  1082 => (x"62",x"20",x"64",x"6c"),
  1083 => (x"20",x"20",x"3a",x"65"),
  1084 => (x"52",x"48",x"44",x"20"),
  1085 => (x"4f",x"54",x"53",x"59"),
  1086 => (x"50",x"20",x"45",x"4e"),
  1087 => (x"52",x"47",x"4f",x"52"),
  1088 => (x"20",x"2c",x"4d",x"41"),
  1089 => (x"45",x"4d",x"4f",x"53"),
  1090 => (x"52",x"54",x"53",x"20"),
  1091 => (x"0a",x"47",x"4e",x"49"),
  1092 => (x"00",x"00",x"00",x"00"),
  1093 => (x"5f",x"74",x"6e",x"49"),
  1094 => (x"6f",x"4c",x"5f",x"31"),
  1095 => (x"20",x"20",x"3a",x"63"),
  1096 => (x"20",x"20",x"20",x"20"),
  1097 => (x"20",x"20",x"20",x"20"),
  1098 => (x"0a",x"64",x"25",x"20"),
  1099 => (x"00",x"00",x"00",x"00"),
  1100 => (x"20",x"20",x"20",x"20"),
  1101 => (x"20",x"20",x"20",x"20"),
  1102 => (x"75",x"6f",x"68",x"73"),
  1103 => (x"62",x"20",x"64",x"6c"),
  1104 => (x"20",x"20",x"3a",x"65"),
  1105 => (x"0a",x"64",x"25",x"20"),
  1106 => (x"00",x"00",x"00",x"00"),
  1107 => (x"5f",x"74",x"6e",x"49"),
  1108 => (x"6f",x"4c",x"5f",x"32"),
  1109 => (x"20",x"20",x"3a",x"63"),
  1110 => (x"20",x"20",x"20",x"20"),
  1111 => (x"20",x"20",x"20",x"20"),
  1112 => (x"0a",x"64",x"25",x"20"),
  1113 => (x"00",x"00",x"00",x"00"),
  1114 => (x"20",x"20",x"20",x"20"),
  1115 => (x"20",x"20",x"20",x"20"),
  1116 => (x"75",x"6f",x"68",x"73"),
  1117 => (x"62",x"20",x"64",x"6c"),
  1118 => (x"20",x"20",x"3a",x"65"),
  1119 => (x"0a",x"64",x"25",x"20"),
  1120 => (x"00",x"00",x"00",x"00"),
  1121 => (x"5f",x"74",x"6e",x"49"),
  1122 => (x"6f",x"4c",x"5f",x"33"),
  1123 => (x"20",x"20",x"3a",x"63"),
  1124 => (x"20",x"20",x"20",x"20"),
  1125 => (x"20",x"20",x"20",x"20"),
  1126 => (x"0a",x"64",x"25",x"20"),
  1127 => (x"00",x"00",x"00",x"00"),
  1128 => (x"20",x"20",x"20",x"20"),
  1129 => (x"20",x"20",x"20",x"20"),
  1130 => (x"75",x"6f",x"68",x"73"),
  1131 => (x"62",x"20",x"64",x"6c"),
  1132 => (x"20",x"20",x"3a",x"65"),
  1133 => (x"0a",x"64",x"25",x"20"),
  1134 => (x"00",x"00",x"00",x"00"),
  1135 => (x"6d",x"75",x"6e",x"45"),
  1136 => (x"63",x"6f",x"4c",x"5f"),
  1137 => (x"20",x"20",x"20",x"3a"),
  1138 => (x"20",x"20",x"20",x"20"),
  1139 => (x"20",x"20",x"20",x"20"),
  1140 => (x"0a",x"64",x"25",x"20"),
  1141 => (x"00",x"00",x"00",x"00"),
  1142 => (x"20",x"20",x"20",x"20"),
  1143 => (x"20",x"20",x"20",x"20"),
  1144 => (x"75",x"6f",x"68",x"73"),
  1145 => (x"62",x"20",x"64",x"6c"),
  1146 => (x"20",x"20",x"3a",x"65"),
  1147 => (x"0a",x"64",x"25",x"20"),
  1148 => (x"00",x"00",x"00",x"00"),
  1149 => (x"5f",x"72",x"74",x"53"),
  1150 => (x"6f",x"4c",x"5f",x"31"),
  1151 => (x"20",x"20",x"3a",x"63"),
  1152 => (x"20",x"20",x"20",x"20"),
  1153 => (x"20",x"20",x"20",x"20"),
  1154 => (x"0a",x"73",x"25",x"20"),
  1155 => (x"00",x"00",x"00",x"00"),
  1156 => (x"20",x"20",x"20",x"20"),
  1157 => (x"20",x"20",x"20",x"20"),
  1158 => (x"75",x"6f",x"68",x"73"),
  1159 => (x"62",x"20",x"64",x"6c"),
  1160 => (x"20",x"20",x"3a",x"65"),
  1161 => (x"52",x"48",x"44",x"20"),
  1162 => (x"4f",x"54",x"53",x"59"),
  1163 => (x"50",x"20",x"45",x"4e"),
  1164 => (x"52",x"47",x"4f",x"52"),
  1165 => (x"20",x"2c",x"4d",x"41"),
  1166 => (x"54",x"53",x"27",x"31"),
  1167 => (x"52",x"54",x"53",x"20"),
  1168 => (x"0a",x"47",x"4e",x"49"),
  1169 => (x"00",x"00",x"00",x"00"),
  1170 => (x"5f",x"72",x"74",x"53"),
  1171 => (x"6f",x"4c",x"5f",x"32"),
  1172 => (x"20",x"20",x"3a",x"63"),
  1173 => (x"20",x"20",x"20",x"20"),
  1174 => (x"20",x"20",x"20",x"20"),
  1175 => (x"0a",x"73",x"25",x"20"),
  1176 => (x"00",x"00",x"00",x"00"),
  1177 => (x"20",x"20",x"20",x"20"),
  1178 => (x"20",x"20",x"20",x"20"),
  1179 => (x"75",x"6f",x"68",x"73"),
  1180 => (x"62",x"20",x"64",x"6c"),
  1181 => (x"20",x"20",x"3a",x"65"),
  1182 => (x"52",x"48",x"44",x"20"),
  1183 => (x"4f",x"54",x"53",x"59"),
  1184 => (x"50",x"20",x"45",x"4e"),
  1185 => (x"52",x"47",x"4f",x"52"),
  1186 => (x"20",x"2c",x"4d",x"41"),
  1187 => (x"44",x"4e",x"27",x"32"),
  1188 => (x"52",x"54",x"53",x"20"),
  1189 => (x"0a",x"47",x"4e",x"49"),
  1190 => (x"00",x"00",x"00",x"00"),
  1191 => (x"00",x"00",x"00",x"0a"),
  1192 => (x"72",x"65",x"73",x"55"),
  1193 => (x"6d",x"69",x"74",x"20"),
  1194 => (x"25",x"20",x"3a",x"65"),
  1195 => (x"1e",x"00",x"0a",x"64"),
  1196 => (x"66",x"c8",x"1e",x"73"),
  1197 => (x"49",x"66",x"cc",x"4b"),
  1198 => (x"ab",x"c2",x"79",x"73"),
  1199 => (x"c1",x"87",x"c4",x"05"),
  1200 => (x"c0",x"87",x"c2",x"4a"),
  1201 => (x"05",x"9a",x"72",x"4a"),
  1202 => (x"79",x"c3",x"87",x"c2"),
  1203 => (x"d8",x"02",x"ab",x"c0"),
  1204 => (x"02",x"ab",x"c1",x"87"),
  1205 => (x"ab",x"c2",x"87",x"d7"),
  1206 => (x"87",x"e5",x"c0",x"02"),
  1207 => (x"c0",x"02",x"ab",x"c3"),
  1208 => (x"ab",x"c4",x"87",x"e5"),
  1209 => (x"de",x"87",x"de",x"02"),
  1210 => (x"da",x"79",x"c0",x"87"),
  1211 => (x"e8",x"d1",x"c1",x"87"),
  1212 => (x"e4",x"c1",x"48",x"bf"),
  1213 => (x"c4",x"06",x"a8",x"b7"),
  1214 => (x"ca",x"79",x"c0",x"87"),
  1215 => (x"c6",x"79",x"c3",x"87"),
  1216 => (x"c2",x"79",x"c1",x"87"),
  1217 => (x"26",x"79",x"c2",x"87"),
  1218 => (x"1e",x"4f",x"26",x"4b"),
  1219 => (x"c2",x"49",x"66",x"c4"),
  1220 => (x"48",x"66",x"c8",x"81"),
  1221 => (x"66",x"cc",x"80",x"71"),
  1222 => (x"26",x"08",x"78",x"08"),
  1223 => (x"1e",x"73",x"1e",x"4f"),
  1224 => (x"1e",x"75",x"1e",x"74"),
  1225 => (x"e4",x"c0",x"86",x"f4"),
  1226 => (x"84",x"c5",x"4c",x"66"),
  1227 => (x"90",x"c4",x"48",x"74"),
  1228 => (x"dc",x"58",x"a6",x"c8"),
  1229 => (x"66",x"c4",x"48",x"66"),
  1230 => (x"58",x"a6",x"c4",x"80"),
  1231 => (x"e8",x"c0",x"48",x"6e"),
  1232 => (x"a6",x"c8",x"78",x"66"),
  1233 => (x"78",x"a4",x"c1",x"48"),
  1234 => (x"dc",x"91",x"c4",x"49"),
  1235 => (x"e8",x"c0",x"81",x"66"),
  1236 => (x"a4",x"de",x"79",x"66"),
  1237 => (x"dc",x"91",x"c4",x"49"),
  1238 => (x"79",x"74",x"81",x"66"),
  1239 => (x"ac",x"b7",x"66",x"c8"),
  1240 => (x"87",x"e0",x"c0",x"01"),
  1241 => (x"c8",x"c3",x"49",x"74"),
  1242 => (x"66",x"e0",x"c0",x"91"),
  1243 => (x"71",x"4d",x"c4",x"81"),
  1244 => (x"82",x"66",x"c4",x"4a"),
  1245 => (x"74",x"4b",x"66",x"c8"),
  1246 => (x"74",x"83",x"c1",x"8b"),
  1247 => (x"c1",x"82",x"75",x"7a"),
  1248 => (x"87",x"f7",x"01",x"8b"),
  1249 => (x"c8",x"c3",x"4a",x"74"),
  1250 => (x"66",x"e0",x"c0",x"92"),
  1251 => (x"c1",x"49",x"74",x"82"),
  1252 => (x"72",x"91",x"c4",x"89"),
  1253 => (x"48",x"69",x"49",x"a1"),
  1254 => (x"79",x"70",x"80",x"c1"),
  1255 => (x"c3",x"49",x"a4",x"d4"),
  1256 => (x"e0",x"c0",x"91",x"c8"),
  1257 => (x"66",x"c4",x"81",x"66"),
  1258 => (x"79",x"bf",x"6e",x"81"),
  1259 => (x"48",x"e8",x"d1",x"c1"),
  1260 => (x"8e",x"f4",x"78",x"c5"),
  1261 => (x"4c",x"26",x"4d",x"26"),
  1262 => (x"4f",x"26",x"4b",x"26"),
  1263 => (x"97",x"1e",x"73",x"1e"),
  1264 => (x"73",x"4b",x"66",x"c8"),
  1265 => (x"66",x"cc",x"97",x"4a"),
  1266 => (x"aa",x"b7",x"71",x"49"),
  1267 => (x"c0",x"87",x"c4",x"02"),
  1268 => (x"c1",x"87",x"c7",x"48"),
  1269 => (x"5b",x"97",x"f4",x"d1"),
  1270 => (x"4b",x"26",x"48",x"c1"),
  1271 => (x"73",x"1e",x"4f",x"26"),
  1272 => (x"75",x"1e",x"74",x"1e"),
  1273 => (x"c2",x"86",x"f8",x"1e"),
  1274 => (x"49",x"66",x"dc",x"4d"),
  1275 => (x"66",x"d8",x"81",x"c1"),
  1276 => (x"a1",x"84",x"c2",x"4c"),
  1277 => (x"49",x"6b",x"97",x"4b"),
  1278 => (x"7e",x"97",x"6c",x"97"),
  1279 => (x"71",x"4a",x"6e",x"97"),
  1280 => (x"c7",x"02",x"aa",x"b7"),
  1281 => (x"48",x"a6",x"c4",x"87"),
  1282 => (x"87",x"cc",x"78",x"c0"),
  1283 => (x"48",x"f0",x"d1",x"c1"),
  1284 => (x"c4",x"50",x"6e",x"97"),
  1285 => (x"78",x"c1",x"48",x"a6"),
  1286 => (x"c4",x"05",x"66",x"c4"),
  1287 => (x"83",x"85",x"c1",x"87"),
  1288 => (x"ad",x"b7",x"c2",x"84"),
  1289 => (x"87",x"cd",x"ff",x"06"),
  1290 => (x"dc",x"4a",x"66",x"d8"),
  1291 => (x"fd",x"fe",x"49",x"66"),
  1292 => (x"b7",x"c0",x"87",x"ef"),
  1293 => (x"87",x"cb",x"06",x"a8"),
  1294 => (x"48",x"e8",x"d1",x"c1"),
  1295 => (x"c1",x"78",x"a5",x"c7"),
  1296 => (x"c0",x"87",x"c2",x"48"),
  1297 => (x"26",x"8e",x"f8",x"48"),
  1298 => (x"26",x"4c",x"26",x"4d"),
  1299 => (x"26",x"4f",x"26",x"4b"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
