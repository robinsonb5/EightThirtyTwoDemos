
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"3b",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"38"),
    10 => (x"20",x"00",x"27",x"4f"),
    11 => (x"27",x"4e",x"00",x"00"),
    12 => (x"00",x"00",x"13",x"97"),
    13 => (x"87",x"fd",x"00",x"0f"),
    14 => (x"4f",x"87",x"fd",x"00"),
    15 => (x"ff",x"86",x"fc",x"1e"),
    16 => (x"48",x"69",x"49",x"c0"),
    17 => (x"c4",x"98",x"c0",x"c4"),
    18 => (x"02",x"6e",x"58",x"a6"),
    19 => (x"66",x"c8",x"87",x"f4"),
    20 => (x"8e",x"fc",x"48",x"79"),
    21 => (x"5e",x"0e",x"4f",x"26"),
    22 => (x"cc",x"0e",x"5c",x"5b"),
    23 => (x"4c",x"c0",x"4b",x"66"),
    24 => (x"ff",x"c3",x"4a",x"13"),
    25 => (x"02",x"9a",x"72",x"9a"),
    26 => (x"49",x"72",x"87",x"d5"),
    27 => (x"cb",x"ff",x"1e",x"71"),
    28 => (x"c1",x"86",x"c4",x"87"),
    29 => (x"c3",x"4a",x"13",x"84"),
    30 => (x"9a",x"72",x"9a",x"ff"),
    31 => (x"74",x"87",x"eb",x"05"),
    32 => (x"26",x"4c",x"26",x"48"),
    33 => (x"0e",x"4f",x"26",x"4b"),
    34 => (x"5d",x"5c",x"5b",x"5e"),
    35 => (x"c0",x"86",x"f0",x"0e"),
    36 => (x"48",x"a6",x"c4",x"4b"),
    37 => (x"e4",x"c0",x"78",x"c0"),
    38 => (x"e0",x"c0",x"4c",x"a6"),
    39 => (x"c1",x"48",x"49",x"66"),
    40 => (x"a6",x"e4",x"c0",x"80"),
    41 => (x"fe",x"4a",x"11",x"58"),
    42 => (x"72",x"ba",x"82",x"c0"),
    43 => (x"d3",x"c4",x"02",x"9a"),
    44 => (x"02",x"66",x"c4",x"87"),
    45 => (x"c4",x"87",x"e2",x"c3"),
    46 => (x"78",x"c0",x"48",x"a6"),
    47 => (x"f0",x"c0",x"49",x"72"),
    48 => (x"f2",x"c2",x"02",x"aa"),
    49 => (x"a9",x"e3",x"c1",x"87"),
    50 => (x"87",x"f3",x"c2",x"02"),
    51 => (x"02",x"a9",x"e4",x"c1"),
    52 => (x"c1",x"87",x"e1",x"c0"),
    53 => (x"c2",x"02",x"a9",x"ec"),
    54 => (x"f0",x"c1",x"87",x"dd"),
    55 => (x"87",x"d4",x"02",x"a9"),
    56 => (x"02",x"a9",x"f3",x"c1"),
    57 => (x"c1",x"87",x"fc",x"c1"),
    58 => (x"c7",x"02",x"a9",x"f5"),
    59 => (x"a9",x"f8",x"c1",x"87"),
    60 => (x"87",x"dc",x"c2",x"05"),
    61 => (x"49",x"74",x"84",x"c4"),
    62 => (x"48",x"76",x"89",x"c4"),
    63 => (x"02",x"6e",x"78",x"69"),
    64 => (x"c8",x"87",x"d3",x"c1"),
    65 => (x"cc",x"78",x"c0",x"80"),
    66 => (x"78",x"c0",x"48",x"a6"),
    67 => (x"b7",x"dc",x"49",x"6e"),
    68 => (x"cf",x"4a",x"71",x"29"),
    69 => (x"c4",x"48",x"6e",x"9a"),
    70 => (x"58",x"a6",x"c4",x"30"),
    71 => (x"c5",x"02",x"9a",x"72"),
    72 => (x"48",x"a6",x"c8",x"87"),
    73 => (x"aa",x"c9",x"78",x"c1"),
    74 => (x"c0",x"87",x"c5",x"06"),
    75 => (x"87",x"c3",x"82",x"f7"),
    76 => (x"c8",x"82",x"f0",x"c0"),
    77 => (x"87",x"c9",x"02",x"66"),
    78 => (x"ff",x"fb",x"1e",x"72"),
    79 => (x"c1",x"86",x"c4",x"87"),
    80 => (x"48",x"66",x"cc",x"83"),
    81 => (x"a6",x"d0",x"80",x"c1"),
    82 => (x"48",x"66",x"cc",x"58"),
    83 => (x"04",x"a8",x"b7",x"c8"),
    84 => (x"c1",x"87",x"f9",x"fe"),
    85 => (x"f0",x"c0",x"87",x"d7"),
    86 => (x"87",x"e0",x"fb",x"1e"),
    87 => (x"83",x"c1",x"86",x"c4"),
    88 => (x"c4",x"87",x"ca",x"c1"),
    89 => (x"c4",x"49",x"74",x"84"),
    90 => (x"fb",x"1e",x"69",x"89"),
    91 => (x"86",x"c4",x"87",x"e8"),
    92 => (x"83",x"71",x"49",x"70"),
    93 => (x"c4",x"87",x"f6",x"c0"),
    94 => (x"78",x"c1",x"48",x"a6"),
    95 => (x"c4",x"87",x"ee",x"c0"),
    96 => (x"c4",x"49",x"74",x"84"),
    97 => (x"fa",x"1e",x"69",x"89"),
    98 => (x"86",x"c4",x"87",x"f2"),
    99 => (x"87",x"dd",x"83",x"c1"),
   100 => (x"e7",x"fa",x"1e",x"72"),
   101 => (x"d4",x"86",x"c4",x"87"),
   102 => (x"aa",x"e5",x"c0",x"87"),
   103 => (x"c4",x"87",x"c7",x"05"),
   104 => (x"78",x"c1",x"48",x"a6"),
   105 => (x"1e",x"72",x"87",x"c7"),
   106 => (x"c4",x"87",x"d1",x"fa"),
   107 => (x"66",x"e0",x"c0",x"86"),
   108 => (x"80",x"c1",x"48",x"49"),
   109 => (x"58",x"a6",x"e4",x"c0"),
   110 => (x"c0",x"fe",x"4a",x"11"),
   111 => (x"9a",x"72",x"ba",x"82"),
   112 => (x"87",x"ed",x"fb",x"05"),
   113 => (x"8e",x"f0",x"48",x"73"),
   114 => (x"4c",x"26",x"4d",x"26"),
   115 => (x"4f",x"26",x"4b",x"26"),
   116 => (x"e8",x"0e",x"5e",x"0e"),
   117 => (x"4a",x"d4",x"ff",x"86"),
   118 => (x"6a",x"7a",x"ff",x"c3"),
   119 => (x"7a",x"ff",x"c3",x"49"),
   120 => (x"30",x"c8",x"48",x"6a"),
   121 => (x"c8",x"58",x"a6",x"c4"),
   122 => (x"b1",x"6e",x"59",x"a6"),
   123 => (x"6a",x"7a",x"ff",x"c3"),
   124 => (x"cc",x"30",x"d0",x"48"),
   125 => (x"a6",x"d0",x"58",x"a6"),
   126 => (x"b1",x"66",x"c8",x"59"),
   127 => (x"6a",x"7a",x"ff",x"c3"),
   128 => (x"d4",x"30",x"d8",x"48"),
   129 => (x"a6",x"d8",x"58",x"a6"),
   130 => (x"b1",x"66",x"d0",x"59"),
   131 => (x"8e",x"e8",x"48",x"71"),
   132 => (x"5e",x"0e",x"4f",x"26"),
   133 => (x"ff",x"86",x"f4",x"0e"),
   134 => (x"ff",x"c3",x"4a",x"d4"),
   135 => (x"c3",x"49",x"6a",x"7a"),
   136 => (x"48",x"71",x"7a",x"ff"),
   137 => (x"a6",x"c4",x"30",x"c8"),
   138 => (x"6e",x"49",x"6a",x"58"),
   139 => (x"7a",x"ff",x"c3",x"b1"),
   140 => (x"30",x"c8",x"48",x"71"),
   141 => (x"6a",x"58",x"a6",x"c8"),
   142 => (x"b1",x"66",x"c4",x"49"),
   143 => (x"71",x"7a",x"ff",x"c3"),
   144 => (x"cc",x"30",x"c8",x"48"),
   145 => (x"49",x"6a",x"58",x"a6"),
   146 => (x"71",x"b1",x"66",x"c8"),
   147 => (x"26",x"8e",x"f4",x"48"),
   148 => (x"5b",x"5e",x"0e",x"4f"),
   149 => (x"c3",x"0e",x"5d",x"5c"),
   150 => (x"d4",x"ff",x"4d",x"ff"),
   151 => (x"48",x"66",x"d0",x"4c"),
   152 => (x"70",x"98",x"ff",x"c3"),
   153 => (x"d8",x"d3",x"c1",x"7c"),
   154 => (x"87",x"c8",x"05",x"bf"),
   155 => (x"c9",x"48",x"66",x"d4"),
   156 => (x"58",x"a6",x"d8",x"30"),
   157 => (x"d8",x"49",x"66",x"d4"),
   158 => (x"c3",x"48",x"71",x"29"),
   159 => (x"7c",x"70",x"98",x"ff"),
   160 => (x"d0",x"49",x"66",x"d4"),
   161 => (x"c3",x"48",x"71",x"29"),
   162 => (x"7c",x"70",x"98",x"ff"),
   163 => (x"c8",x"49",x"66",x"d4"),
   164 => (x"c3",x"48",x"71",x"29"),
   165 => (x"7c",x"70",x"98",x"ff"),
   166 => (x"c3",x"48",x"66",x"d4"),
   167 => (x"7c",x"70",x"98",x"ff"),
   168 => (x"d0",x"49",x"66",x"d0"),
   169 => (x"c3",x"48",x"71",x"29"),
   170 => (x"7c",x"70",x"98",x"ff"),
   171 => (x"f0",x"c9",x"4b",x"6c"),
   172 => (x"ab",x"75",x"4a",x"ff"),
   173 => (x"75",x"87",x"ce",x"05"),
   174 => (x"c1",x"4b",x"6c",x"7c"),
   175 => (x"87",x"c5",x"02",x"8a"),
   176 => (x"f2",x"02",x"ab",x"75"),
   177 => (x"26",x"48",x"73",x"87"),
   178 => (x"26",x"4c",x"26",x"4d"),
   179 => (x"1e",x"4f",x"26",x"4b"),
   180 => (x"d4",x"ff",x"49",x"c0"),
   181 => (x"78",x"ff",x"c3",x"48"),
   182 => (x"c8",x"c3",x"81",x"c1"),
   183 => (x"f1",x"04",x"a9",x"b7"),
   184 => (x"0e",x"4f",x"26",x"87"),
   185 => (x"5d",x"5c",x"5b",x"5e"),
   186 => (x"f0",x"ff",x"c0",x"0e"),
   187 => (x"c1",x"4d",x"f7",x"c1"),
   188 => (x"c0",x"c0",x"c0",x"c0"),
   189 => (x"d6",x"ff",x"4b",x"c0"),
   190 => (x"df",x"f8",x"c4",x"87"),
   191 => (x"75",x"1e",x"c0",x"4c"),
   192 => (x"87",x"cd",x"fd",x"1e"),
   193 => (x"a8",x"c1",x"86",x"c8"),
   194 => (x"87",x"e5",x"c0",x"05"),
   195 => (x"c3",x"48",x"d4",x"ff"),
   196 => (x"1e",x"73",x"78",x"ff"),
   197 => (x"c1",x"f0",x"e1",x"c0"),
   198 => (x"f4",x"fc",x"1e",x"e9"),
   199 => (x"70",x"86",x"c8",x"87"),
   200 => (x"87",x"ca",x"05",x"98"),
   201 => (x"c3",x"48",x"d4",x"ff"),
   202 => (x"48",x"c1",x"78",x"ff"),
   203 => (x"de",x"fe",x"87",x"cb"),
   204 => (x"05",x"8c",x"c1",x"87"),
   205 => (x"c0",x"87",x"c6",x"ff"),
   206 => (x"26",x"4d",x"26",x"48"),
   207 => (x"26",x"4b",x"26",x"4c"),
   208 => (x"5b",x"5e",x"0e",x"4f"),
   209 => (x"ff",x"c0",x"0e",x"5c"),
   210 => (x"4c",x"c1",x"c1",x"f0"),
   211 => (x"c3",x"48",x"d4",x"ff"),
   212 => (x"e5",x"c0",x"78",x"ff"),
   213 => (x"fd",x"f3",x"1e",x"d8"),
   214 => (x"d3",x"86",x"c4",x"87"),
   215 => (x"74",x"1e",x"c0",x"4b"),
   216 => (x"87",x"ed",x"fb",x"1e"),
   217 => (x"98",x"70",x"86",x"c8"),
   218 => (x"ff",x"87",x"ca",x"05"),
   219 => (x"ff",x"c3",x"48",x"d4"),
   220 => (x"cb",x"48",x"c1",x"78"),
   221 => (x"87",x"d7",x"fd",x"87"),
   222 => (x"ff",x"05",x"8b",x"c1"),
   223 => (x"48",x"c0",x"87",x"df"),
   224 => (x"4b",x"26",x"4c",x"26"),
   225 => (x"5e",x"0e",x"4f",x"26"),
   226 => (x"0e",x"5d",x"5c",x"5b"),
   227 => (x"fc",x"4c",x"d4",x"ff"),
   228 => (x"ea",x"c6",x"87",x"fd"),
   229 => (x"f0",x"e1",x"c0",x"1e"),
   230 => (x"fa",x"1e",x"c8",x"c1"),
   231 => (x"86",x"c8",x"87",x"f3"),
   232 => (x"1e",x"73",x"4b",x"70"),
   233 => (x"f3",x"1e",x"d2",x"d2"),
   234 => (x"86",x"c8",x"87",x"dd"),
   235 => (x"c8",x"02",x"ab",x"c1"),
   236 => (x"87",x"cd",x"fe",x"87"),
   237 => (x"cf",x"c2",x"48",x"c0"),
   238 => (x"87",x"d6",x"f9",x"87"),
   239 => (x"ff",x"cf",x"49",x"70"),
   240 => (x"ea",x"c6",x"99",x"ff"),
   241 => (x"87",x"c8",x"02",x"a9"),
   242 => (x"c0",x"87",x"f6",x"fd"),
   243 => (x"87",x"f8",x"c1",x"48"),
   244 => (x"c0",x"7c",x"ff",x"c3"),
   245 => (x"ca",x"fc",x"4d",x"f1"),
   246 => (x"02",x"98",x"70",x"87"),
   247 => (x"c0",x"87",x"d0",x"c1"),
   248 => (x"f0",x"ff",x"c0",x"1e"),
   249 => (x"f9",x"1e",x"fa",x"c1"),
   250 => (x"86",x"c8",x"87",x"e7"),
   251 => (x"9b",x"73",x"4b",x"70"),
   252 => (x"87",x"f1",x"c0",x"05"),
   253 => (x"d0",x"d1",x"1e",x"73"),
   254 => (x"87",x"cb",x"f2",x"1e"),
   255 => (x"ff",x"c3",x"86",x"c8"),
   256 => (x"73",x"4b",x"6c",x"7c"),
   257 => (x"1e",x"dc",x"d1",x"1e"),
   258 => (x"c8",x"87",x"fc",x"f1"),
   259 => (x"7c",x"ff",x"c3",x"86"),
   260 => (x"73",x"7c",x"7c",x"7c"),
   261 => (x"99",x"c0",x"c1",x"49"),
   262 => (x"c1",x"87",x"c5",x"02"),
   263 => (x"87",x"e8",x"c0",x"48"),
   264 => (x"e3",x"c0",x"48",x"c0"),
   265 => (x"d1",x"1e",x"73",x"87"),
   266 => (x"da",x"f1",x"1e",x"ea"),
   267 => (x"c2",x"86",x"c8",x"87"),
   268 => (x"87",x"cc",x"05",x"ad"),
   269 => (x"f1",x"1e",x"f6",x"d1"),
   270 => (x"86",x"c4",x"87",x"cd"),
   271 => (x"87",x"c8",x"48",x"c0"),
   272 => (x"fe",x"05",x"8d",x"c1"),
   273 => (x"48",x"c0",x"87",x"d0"),
   274 => (x"4c",x"26",x"4d",x"26"),
   275 => (x"4f",x"26",x"4b",x"26"),
   276 => (x"35",x"44",x"4d",x"43"),
   277 => (x"64",x"25",x"20",x"38"),
   278 => (x"00",x"20",x"20",x"0a"),
   279 => (x"35",x"44",x"4d",x"43"),
   280 => (x"20",x"32",x"5f",x"38"),
   281 => (x"20",x"0a",x"64",x"25"),
   282 => (x"4d",x"43",x"00",x"20"),
   283 => (x"20",x"38",x"35",x"44"),
   284 => (x"20",x"0a",x"64",x"25"),
   285 => (x"44",x"53",x"00",x"20"),
   286 => (x"49",x"20",x"43",x"48"),
   287 => (x"69",x"74",x"69",x"6e"),
   288 => (x"7a",x"69",x"6c",x"61"),
   289 => (x"6f",x"69",x"74",x"61"),
   290 => (x"72",x"65",x"20",x"6e"),
   291 => (x"21",x"72",x"6f",x"72"),
   292 => (x"6d",x"63",x"00",x"0a"),
   293 => (x"4d",x"43",x"5f",x"64"),
   294 => (x"72",x"20",x"38",x"44"),
   295 => (x"6f",x"70",x"73",x"65"),
   296 => (x"3a",x"65",x"73",x"6e"),
   297 => (x"0a",x"64",x"25",x"20"),
   298 => (x"5b",x"5e",x"0e",x"00"),
   299 => (x"fc",x"0e",x"5d",x"5c"),
   300 => (x"4c",x"d0",x"ff",x"86"),
   301 => (x"4b",x"c0",x"c0",x"c8"),
   302 => (x"48",x"d8",x"d3",x"c1"),
   303 => (x"d2",x"d6",x"78",x"c1"),
   304 => (x"87",x"d2",x"ee",x"1e"),
   305 => (x"4d",x"c7",x"86",x"c4"),
   306 => (x"98",x"73",x"48",x"6c"),
   307 => (x"6e",x"58",x"a6",x"c4"),
   308 => (x"6c",x"87",x"cc",x"02"),
   309 => (x"c4",x"98",x"73",x"48"),
   310 => (x"05",x"6e",x"58",x"a6"),
   311 => (x"c0",x"87",x"f4",x"ff"),
   312 => (x"87",x"eb",x"f7",x"7c"),
   313 => (x"98",x"73",x"48",x"6c"),
   314 => (x"6e",x"58",x"a6",x"c4"),
   315 => (x"6c",x"87",x"cc",x"02"),
   316 => (x"c4",x"98",x"73",x"48"),
   317 => (x"05",x"6e",x"58",x"a6"),
   318 => (x"c1",x"87",x"f4",x"ff"),
   319 => (x"c0",x"1e",x"c0",x"7c"),
   320 => (x"c0",x"c1",x"d0",x"e5"),
   321 => (x"87",x"c9",x"f5",x"1e"),
   322 => (x"a8",x"c1",x"86",x"c8"),
   323 => (x"87",x"c2",x"c0",x"05"),
   324 => (x"ad",x"c2",x"4d",x"c1"),
   325 => (x"87",x"cd",x"c0",x"05"),
   326 => (x"ec",x"1e",x"cd",x"d6"),
   327 => (x"86",x"c4",x"87",x"f8"),
   328 => (x"de",x"c1",x"48",x"c0"),
   329 => (x"05",x"8d",x"c1",x"87"),
   330 => (x"f9",x"87",x"dd",x"fe"),
   331 => (x"d3",x"c1",x"87",x"d8"),
   332 => (x"d3",x"c1",x"58",x"dc"),
   333 => (x"c0",x"05",x"bf",x"d8"),
   334 => (x"1e",x"c1",x"87",x"cd"),
   335 => (x"c1",x"f0",x"ff",x"c0"),
   336 => (x"cc",x"f4",x"1e",x"d0"),
   337 => (x"ff",x"86",x"c8",x"87"),
   338 => (x"ff",x"c3",x"48",x"d4"),
   339 => (x"87",x"ca",x"ca",x"78"),
   340 => (x"58",x"e0",x"d3",x"c1"),
   341 => (x"bf",x"dc",x"d3",x"c1"),
   342 => (x"1e",x"d6",x"d6",x"1e"),
   343 => (x"c8",x"87",x"e8",x"ec"),
   344 => (x"73",x"48",x"6c",x"86"),
   345 => (x"58",x"a6",x"c4",x"98"),
   346 => (x"cc",x"c0",x"02",x"6e"),
   347 => (x"73",x"48",x"6c",x"87"),
   348 => (x"58",x"a6",x"c4",x"98"),
   349 => (x"f4",x"ff",x"05",x"6e"),
   350 => (x"ff",x"7c",x"c0",x"87"),
   351 => (x"ff",x"c3",x"48",x"d4"),
   352 => (x"fc",x"48",x"c1",x"78"),
   353 => (x"26",x"4d",x"26",x"8e"),
   354 => (x"26",x"4b",x"26",x"4c"),
   355 => (x"52",x"45",x"49",x"4f"),
   356 => (x"50",x"53",x"00",x"52"),
   357 => (x"44",x"53",x"00",x"49"),
   358 => (x"72",x"61",x"63",x"20"),
   359 => (x"69",x"73",x"20",x"64"),
   360 => (x"69",x"20",x"65",x"7a"),
   361 => (x"64",x"25",x"20",x"73"),
   362 => (x"5e",x"0e",x"00",x"0a"),
   363 => (x"0e",x"5d",x"5c",x"5b"),
   364 => (x"c0",x"c8",x"86",x"fc"),
   365 => (x"ff",x"c3",x"4d",x"c0"),
   366 => (x"4b",x"d4",x"ff",x"4c"),
   367 => (x"d0",x"ff",x"7b",x"74"),
   368 => (x"98",x"75",x"48",x"bf"),
   369 => (x"6e",x"58",x"a6",x"c4"),
   370 => (x"87",x"ce",x"c0",x"02"),
   371 => (x"48",x"bf",x"d0",x"ff"),
   372 => (x"a6",x"c4",x"98",x"75"),
   373 => (x"ff",x"05",x"6e",x"58"),
   374 => (x"d0",x"ff",x"87",x"f2"),
   375 => (x"78",x"c1",x"c4",x"48"),
   376 => (x"66",x"d4",x"7b",x"74"),
   377 => (x"f0",x"ff",x"c0",x"1e"),
   378 => (x"f1",x"1e",x"d8",x"c1"),
   379 => (x"86",x"c8",x"87",x"e3"),
   380 => (x"c0",x"02",x"98",x"70"),
   381 => (x"d2",x"da",x"87",x"cd"),
   382 => (x"87",x"da",x"e9",x"1e"),
   383 => (x"48",x"c1",x"86",x"c4"),
   384 => (x"74",x"87",x"c5",x"c2"),
   385 => (x"7b",x"fe",x"c3",x"7b"),
   386 => (x"78",x"c0",x"48",x"76"),
   387 => (x"25",x"4d",x"66",x"d8"),
   388 => (x"d8",x"4a",x"71",x"49"),
   389 => (x"48",x"72",x"2a",x"b7"),
   390 => (x"7b",x"70",x"98",x"74"),
   391 => (x"b7",x"d0",x"4a",x"71"),
   392 => (x"74",x"48",x"72",x"2a"),
   393 => (x"71",x"7b",x"70",x"98"),
   394 => (x"2a",x"b7",x"c8",x"4a"),
   395 => (x"98",x"74",x"48",x"72"),
   396 => (x"48",x"71",x"7b",x"70"),
   397 => (x"7b",x"70",x"98",x"74"),
   398 => (x"80",x"c1",x"48",x"6e"),
   399 => (x"6e",x"58",x"a6",x"c4"),
   400 => (x"b7",x"c0",x"c2",x"48"),
   401 => (x"c6",x"ff",x"04",x"a8"),
   402 => (x"c0",x"c0",x"c8",x"87"),
   403 => (x"74",x"7b",x"74",x"4d"),
   404 => (x"d8",x"7b",x"74",x"7b"),
   405 => (x"74",x"49",x"e0",x"da"),
   406 => (x"c0",x"05",x"6b",x"7b"),
   407 => (x"89",x"c1",x"87",x"c6"),
   408 => (x"87",x"f3",x"ff",x"05"),
   409 => (x"d0",x"ff",x"7b",x"74"),
   410 => (x"98",x"75",x"48",x"bf"),
   411 => (x"6e",x"58",x"a6",x"c4"),
   412 => (x"87",x"ce",x"c0",x"02"),
   413 => (x"48",x"bf",x"d0",x"ff"),
   414 => (x"a6",x"c4",x"98",x"75"),
   415 => (x"ff",x"05",x"6e",x"58"),
   416 => (x"d0",x"ff",x"87",x"f2"),
   417 => (x"48",x"78",x"c0",x"48"),
   418 => (x"4d",x"26",x"8e",x"fc"),
   419 => (x"4b",x"26",x"4c",x"26"),
   420 => (x"72",x"57",x"4f",x"26"),
   421 => (x"20",x"65",x"74",x"69"),
   422 => (x"6c",x"69",x"61",x"66"),
   423 => (x"00",x"0a",x"64",x"65"),
   424 => (x"5c",x"5b",x"5e",x"0e"),
   425 => (x"d4",x"ff",x"0e",x"5d"),
   426 => (x"4c",x"66",x"d4",x"4d"),
   427 => (x"c0",x"4b",x"66",x"d0"),
   428 => (x"cd",x"ee",x"c5",x"4a"),
   429 => (x"ff",x"c3",x"49",x"df"),
   430 => (x"c3",x"48",x"6d",x"7d"),
   431 => (x"c1",x"05",x"a8",x"fe"),
   432 => (x"d3",x"c1",x"87",x"d4"),
   433 => (x"78",x"c0",x"48",x"d4"),
   434 => (x"04",x"ac",x"b7",x"c4"),
   435 => (x"eb",x"87",x"dc",x"c0"),
   436 => (x"49",x"70",x"87",x"fe"),
   437 => (x"83",x"c4",x"7b",x"71"),
   438 => (x"bf",x"d4",x"d3",x"c1"),
   439 => (x"c1",x"80",x"71",x"48"),
   440 => (x"c4",x"58",x"d8",x"d3"),
   441 => (x"03",x"ac",x"b7",x"8c"),
   442 => (x"c0",x"87",x"e4",x"ff"),
   443 => (x"c0",x"06",x"ac",x"b7"),
   444 => (x"ff",x"c3",x"87",x"e1"),
   445 => (x"71",x"49",x"6d",x"7d"),
   446 => (x"ff",x"c3",x"7b",x"97"),
   447 => (x"c1",x"83",x"c1",x"98"),
   448 => (x"48",x"bf",x"d4",x"d3"),
   449 => (x"d3",x"c1",x"80",x"71"),
   450 => (x"8c",x"c1",x"58",x"d8"),
   451 => (x"01",x"ac",x"b7",x"c0"),
   452 => (x"c1",x"87",x"df",x"ff"),
   453 => (x"89",x"c1",x"4a",x"49"),
   454 => (x"87",x"da",x"fe",x"05"),
   455 => (x"72",x"7d",x"ff",x"c3"),
   456 => (x"26",x"4d",x"26",x"48"),
   457 => (x"26",x"4b",x"26",x"4c"),
   458 => (x"5b",x"5e",x"0e",x"4f"),
   459 => (x"fc",x"0e",x"5d",x"5c"),
   460 => (x"4c",x"d0",x"ff",x"86"),
   461 => (x"4b",x"c0",x"c0",x"c8"),
   462 => (x"d4",x"ff",x"4d",x"c0"),
   463 => (x"78",x"ff",x"c3",x"48"),
   464 => (x"98",x"73",x"48",x"6c"),
   465 => (x"6e",x"58",x"a6",x"c4"),
   466 => (x"87",x"cc",x"c0",x"02"),
   467 => (x"98",x"73",x"48",x"6c"),
   468 => (x"6e",x"58",x"a6",x"c4"),
   469 => (x"87",x"f4",x"ff",x"05"),
   470 => (x"ff",x"7c",x"c1",x"c4"),
   471 => (x"ff",x"c3",x"48",x"d4"),
   472 => (x"1e",x"66",x"d4",x"78"),
   473 => (x"c1",x"f0",x"ff",x"c0"),
   474 => (x"e4",x"eb",x"1e",x"d1"),
   475 => (x"70",x"86",x"c8",x"87"),
   476 => (x"02",x"99",x"71",x"49"),
   477 => (x"71",x"87",x"d0",x"c0"),
   478 => (x"1e",x"66",x"d8",x"1e"),
   479 => (x"e4",x"1e",x"fa",x"de"),
   480 => (x"86",x"cc",x"87",x"c5"),
   481 => (x"c8",x"87",x"e7",x"c0"),
   482 => (x"66",x"dc",x"1e",x"c0"),
   483 => (x"87",x"d0",x"fc",x"1e"),
   484 => (x"4d",x"70",x"86",x"c8"),
   485 => (x"98",x"73",x"48",x"6c"),
   486 => (x"6e",x"58",x"a6",x"c4"),
   487 => (x"87",x"cc",x"c0",x"02"),
   488 => (x"98",x"73",x"48",x"6c"),
   489 => (x"6e",x"58",x"a6",x"c4"),
   490 => (x"87",x"f4",x"ff",x"05"),
   491 => (x"48",x"75",x"7c",x"c0"),
   492 => (x"4d",x"26",x"8e",x"fc"),
   493 => (x"4b",x"26",x"4c",x"26"),
   494 => (x"65",x"52",x"4f",x"26"),
   495 => (x"63",x"20",x"64",x"61"),
   496 => (x"61",x"6d",x"6d",x"6f"),
   497 => (x"66",x"20",x"64",x"6e"),
   498 => (x"65",x"6c",x"69",x"61"),
   499 => (x"74",x"61",x"20",x"64"),
   500 => (x"20",x"64",x"25",x"20"),
   501 => (x"29",x"64",x"25",x"28"),
   502 => (x"5e",x"0e",x"00",x"0a"),
   503 => (x"0e",x"5d",x"5c",x"5b"),
   504 => (x"1e",x"c0",x"86",x"fc"),
   505 => (x"c1",x"f0",x"ff",x"c0"),
   506 => (x"e4",x"e9",x"1e",x"c9"),
   507 => (x"d2",x"86",x"c8",x"87"),
   508 => (x"e6",x"d3",x"c1",x"1e"),
   509 => (x"87",x"e8",x"fa",x"1e"),
   510 => (x"4d",x"c0",x"86",x"c8"),
   511 => (x"b7",x"d2",x"85",x"c1"),
   512 => (x"f7",x"ff",x"04",x"ad"),
   513 => (x"e6",x"d3",x"c1",x"87"),
   514 => (x"c3",x"49",x"bf",x"97"),
   515 => (x"c0",x"c1",x"99",x"c0"),
   516 => (x"e8",x"c0",x"05",x"a9"),
   517 => (x"ed",x"d3",x"c1",x"87"),
   518 => (x"d0",x"49",x"bf",x"97"),
   519 => (x"ee",x"d3",x"c1",x"31"),
   520 => (x"c8",x"4a",x"bf",x"97"),
   521 => (x"c1",x"b1",x"72",x"32"),
   522 => (x"bf",x"97",x"ef",x"d3"),
   523 => (x"cf",x"b1",x"72",x"4a"),
   524 => (x"99",x"ff",x"ff",x"ff"),
   525 => (x"85",x"c1",x"4d",x"71"),
   526 => (x"eb",x"c2",x"35",x"ca"),
   527 => (x"ef",x"d3",x"c1",x"87"),
   528 => (x"c1",x"4b",x"bf",x"97"),
   529 => (x"c1",x"9b",x"c6",x"33"),
   530 => (x"bf",x"97",x"f0",x"d3"),
   531 => (x"29",x"b7",x"c7",x"49"),
   532 => (x"d3",x"c1",x"b3",x"71"),
   533 => (x"49",x"bf",x"97",x"eb"),
   534 => (x"98",x"cf",x"48",x"71"),
   535 => (x"c1",x"58",x"a6",x"c4"),
   536 => (x"bf",x"97",x"ec",x"d3"),
   537 => (x"ca",x"9c",x"c3",x"4c"),
   538 => (x"ed",x"d3",x"c1",x"34"),
   539 => (x"c2",x"49",x"bf",x"97"),
   540 => (x"c1",x"b4",x"71",x"31"),
   541 => (x"bf",x"97",x"ee",x"d3"),
   542 => (x"99",x"c0",x"c3",x"49"),
   543 => (x"71",x"29",x"b7",x"c6"),
   544 => (x"c4",x"1e",x"74",x"b4"),
   545 => (x"1e",x"73",x"1e",x"66"),
   546 => (x"1e",x"f4",x"e3",x"c0"),
   547 => (x"87",x"f7",x"df",x"ff"),
   548 => (x"83",x"c2",x"86",x"d0"),
   549 => (x"30",x"73",x"48",x"c1"),
   550 => (x"1e",x"73",x"4b",x"70"),
   551 => (x"1e",x"e1",x"e4",x"c0"),
   552 => (x"87",x"e3",x"df",x"ff"),
   553 => (x"48",x"c1",x"86",x"c8"),
   554 => (x"a6",x"c4",x"30",x"6e"),
   555 => (x"c1",x"49",x"74",x"58"),
   556 => (x"73",x"4d",x"71",x"81"),
   557 => (x"1e",x"6e",x"95",x"b7"),
   558 => (x"e4",x"c0",x"1e",x"75"),
   559 => (x"df",x"ff",x"1e",x"ea"),
   560 => (x"86",x"cc",x"87",x"c5"),
   561 => (x"c0",x"c8",x"48",x"6e"),
   562 => (x"c0",x"06",x"a8",x"b7"),
   563 => (x"4b",x"6e",x"87",x"ce"),
   564 => (x"2b",x"b7",x"35",x"c1"),
   565 => (x"ab",x"b7",x"c0",x"c8"),
   566 => (x"87",x"f4",x"ff",x"01"),
   567 => (x"e5",x"c0",x"1e",x"75"),
   568 => (x"de",x"ff",x"1e",x"c0"),
   569 => (x"86",x"c8",x"87",x"e1"),
   570 => (x"8e",x"fc",x"48",x"75"),
   571 => (x"4c",x"26",x"4d",x"26"),
   572 => (x"4f",x"26",x"4b",x"26"),
   573 => (x"69",x"73",x"5f",x"63"),
   574 => (x"6d",x"5f",x"65",x"7a"),
   575 => (x"3a",x"74",x"6c",x"75"),
   576 => (x"2c",x"64",x"25",x"20"),
   577 => (x"61",x"65",x"72",x"20"),
   578 => (x"6c",x"62",x"5f",x"64"),
   579 => (x"6e",x"65",x"6c",x"5f"),
   580 => (x"64",x"25",x"20",x"3a"),
   581 => (x"73",x"63",x"20",x"2c"),
   582 => (x"3a",x"65",x"7a",x"69"),
   583 => (x"0a",x"64",x"25",x"20"),
   584 => (x"6c",x"75",x"4d",x"00"),
   585 => (x"64",x"25",x"20",x"74"),
   586 => (x"64",x"25",x"00",x"0a"),
   587 => (x"6f",x"6c",x"62",x"20"),
   588 => (x"20",x"73",x"6b",x"63"),
   589 => (x"73",x"20",x"66",x"6f"),
   590 => (x"20",x"65",x"7a",x"69"),
   591 => (x"00",x"0a",x"64",x"25"),
   592 => (x"62",x"20",x"64",x"25"),
   593 => (x"6b",x"63",x"6f",x"6c"),
   594 => (x"66",x"6f",x"20",x"73"),
   595 => (x"32",x"31",x"35",x"20"),
   596 => (x"74",x"79",x"62",x"20"),
   597 => (x"00",x"0a",x"73",x"65"),
   598 => (x"00",x"44",x"4d",x"43"),
   599 => (x"0e",x"5b",x"5e",x"0e"),
   600 => (x"66",x"d0",x"4b",x"c0"),
   601 => (x"a8",x"b7",x"c0",x"48"),
   602 => (x"87",x"f6",x"c0",x"06"),
   603 => (x"bf",x"97",x"66",x"c8"),
   604 => (x"82",x"c0",x"fe",x"4a"),
   605 => (x"48",x"66",x"c8",x"ba"),
   606 => (x"a6",x"cc",x"80",x"c1"),
   607 => (x"97",x"66",x"cc",x"58"),
   608 => (x"c0",x"fe",x"49",x"bf"),
   609 => (x"66",x"cc",x"b9",x"81"),
   610 => (x"d0",x"80",x"c1",x"48"),
   611 => (x"b7",x"71",x"58",x"a6"),
   612 => (x"87",x"c4",x"02",x"aa"),
   613 => (x"87",x"cc",x"48",x"c1"),
   614 => (x"66",x"d0",x"83",x"c1"),
   615 => (x"ff",x"04",x"ab",x"b7"),
   616 => (x"48",x"c0",x"87",x"ca"),
   617 => (x"4d",x"26",x"87",x"c4"),
   618 => (x"4b",x"26",x"4c",x"26"),
   619 => (x"5e",x"0e",x"4f",x"26"),
   620 => (x"0e",x"5d",x"5c",x"5b"),
   621 => (x"48",x"c0",x"dc",x"c1"),
   622 => (x"c1",x"c1",x"78",x"c0"),
   623 => (x"da",x"ff",x"1e",x"c8"),
   624 => (x"86",x"c4",x"87",x"d4"),
   625 => (x"1e",x"f8",x"d3",x"c1"),
   626 => (x"dc",x"f5",x"1e",x"c0"),
   627 => (x"70",x"86",x"c8",x"87"),
   628 => (x"87",x"cf",x"05",x"98"),
   629 => (x"1e",x"f4",x"fd",x"c0"),
   630 => (x"87",x"fa",x"d9",x"ff"),
   631 => (x"48",x"c0",x"86",x"c4"),
   632 => (x"c1",x"87",x"d6",x"cb"),
   633 => (x"ff",x"1e",x"d5",x"c1"),
   634 => (x"c4",x"87",x"eb",x"d9"),
   635 => (x"c1",x"4b",x"c0",x"86"),
   636 => (x"c1",x"48",x"ec",x"dc"),
   637 => (x"c1",x"1e",x"c8",x"78"),
   638 => (x"c1",x"1e",x"ec",x"c1"),
   639 => (x"fd",x"1e",x"ee",x"d4"),
   640 => (x"86",x"cc",x"87",x"da"),
   641 => (x"c6",x"05",x"98",x"70"),
   642 => (x"ec",x"dc",x"c1",x"87"),
   643 => (x"c8",x"78",x"c0",x"48"),
   644 => (x"f5",x"c1",x"c1",x"1e"),
   645 => (x"ca",x"d5",x"c1",x"1e"),
   646 => (x"87",x"c0",x"fd",x"1e"),
   647 => (x"98",x"70",x"86",x"cc"),
   648 => (x"c1",x"87",x"c6",x"05"),
   649 => (x"c0",x"48",x"ec",x"dc"),
   650 => (x"ec",x"dc",x"c1",x"78"),
   651 => (x"c1",x"c1",x"1e",x"bf"),
   652 => (x"d9",x"ff",x"1e",x"fe"),
   653 => (x"86",x"c8",x"87",x"d1"),
   654 => (x"bf",x"ec",x"dc",x"c1"),
   655 => (x"87",x"d8",x"c2",x"02"),
   656 => (x"4d",x"f8",x"d3",x"c1"),
   657 => (x"4c",x"f6",x"da",x"c1"),
   658 => (x"9f",x"f6",x"db",x"c1"),
   659 => (x"1e",x"71",x"49",x"bf"),
   660 => (x"49",x"f6",x"db",x"c1"),
   661 => (x"89",x"f8",x"d3",x"c1"),
   662 => (x"1e",x"d0",x"1e",x"71"),
   663 => (x"c0",x"1e",x"c0",x"c8"),
   664 => (x"ff",x"1e",x"e6",x"fe"),
   665 => (x"d4",x"87",x"e0",x"d8"),
   666 => (x"c8",x"49",x"74",x"86"),
   667 => (x"c1",x"4b",x"69",x"81"),
   668 => (x"bf",x"9f",x"f6",x"db"),
   669 => (x"ea",x"d6",x"c5",x"49"),
   670 => (x"d0",x"c0",x"05",x"a9"),
   671 => (x"c8",x"49",x"74",x"87"),
   672 => (x"d9",x"1e",x"69",x"81"),
   673 => (x"86",x"c4",x"87",x"d9"),
   674 => (x"df",x"c0",x"4b",x"70"),
   675 => (x"c7",x"49",x"75",x"87"),
   676 => (x"69",x"9f",x"81",x"fe"),
   677 => (x"d5",x"e9",x"ca",x"49"),
   678 => (x"cf",x"c0",x"02",x"a9"),
   679 => (x"c8",x"fe",x"c0",x"87"),
   680 => (x"f1",x"d6",x"ff",x"1e"),
   681 => (x"c0",x"86",x"c4",x"87"),
   682 => (x"87",x"cd",x"c8",x"48"),
   683 => (x"ff",x"c0",x"1e",x"73"),
   684 => (x"d7",x"ff",x"1e",x"e3"),
   685 => (x"86",x"c8",x"87",x"d1"),
   686 => (x"1e",x"f8",x"d3",x"c1"),
   687 => (x"e8",x"f1",x"1e",x"73"),
   688 => (x"70",x"86",x"c8",x"87"),
   689 => (x"c5",x"c0",x"05",x"98"),
   690 => (x"c7",x"48",x"c0",x"87"),
   691 => (x"ff",x"c0",x"87",x"eb"),
   692 => (x"d6",x"ff",x"1e",x"fb"),
   693 => (x"86",x"c4",x"87",x"c0"),
   694 => (x"1e",x"d1",x"c2",x"c1"),
   695 => (x"87",x"e7",x"d6",x"ff"),
   696 => (x"1e",x"c8",x"86",x"c4"),
   697 => (x"1e",x"e9",x"c2",x"c1"),
   698 => (x"1e",x"ca",x"d5",x"c1"),
   699 => (x"cc",x"87",x"ed",x"f9"),
   700 => (x"05",x"98",x"70",x"86"),
   701 => (x"c1",x"87",x"c9",x"c0"),
   702 => (x"c1",x"48",x"c0",x"dc"),
   703 => (x"87",x"e4",x"c0",x"78"),
   704 => (x"c2",x"c1",x"1e",x"c8"),
   705 => (x"d4",x"c1",x"1e",x"f2"),
   706 => (x"cf",x"f9",x"1e",x"ee"),
   707 => (x"70",x"86",x"cc",x"87"),
   708 => (x"cf",x"c0",x"02",x"98"),
   709 => (x"e2",x"c0",x"c1",x"87"),
   710 => (x"ea",x"d5",x"ff",x"1e"),
   711 => (x"c0",x"86",x"c4",x"87"),
   712 => (x"87",x"d5",x"c6",x"48"),
   713 => (x"97",x"f6",x"db",x"c1"),
   714 => (x"d5",x"c1",x"49",x"bf"),
   715 => (x"cd",x"c0",x"05",x"a9"),
   716 => (x"f7",x"db",x"c1",x"87"),
   717 => (x"c2",x"49",x"bf",x"97"),
   718 => (x"c0",x"02",x"a9",x"ea"),
   719 => (x"48",x"c0",x"87",x"c5"),
   720 => (x"c1",x"87",x"f6",x"c5"),
   721 => (x"bf",x"97",x"f8",x"d3"),
   722 => (x"a9",x"e9",x"c3",x"49"),
   723 => (x"87",x"d2",x"c0",x"02"),
   724 => (x"97",x"f8",x"d3",x"c1"),
   725 => (x"eb",x"c3",x"49",x"bf"),
   726 => (x"c5",x"c0",x"02",x"a9"),
   727 => (x"c5",x"48",x"c0",x"87"),
   728 => (x"d4",x"c1",x"87",x"d7"),
   729 => (x"49",x"bf",x"97",x"c3"),
   730 => (x"c0",x"05",x"99",x"71"),
   731 => (x"d4",x"c1",x"87",x"cc"),
   732 => (x"49",x"bf",x"97",x"c4"),
   733 => (x"c0",x"02",x"a9",x"c2"),
   734 => (x"48",x"c0",x"87",x"c5"),
   735 => (x"c1",x"87",x"fa",x"c4"),
   736 => (x"bf",x"97",x"c5",x"d4"),
   737 => (x"fc",x"db",x"c1",x"48"),
   738 => (x"f8",x"db",x"c1",x"58"),
   739 => (x"4a",x"71",x"49",x"bf"),
   740 => (x"dc",x"c1",x"8a",x"c1"),
   741 => (x"1e",x"72",x"5a",x"c0"),
   742 => (x"c2",x"c1",x"1e",x"71"),
   743 => (x"d3",x"ff",x"1e",x"fb"),
   744 => (x"86",x"cc",x"87",x"e5"),
   745 => (x"97",x"c6",x"d4",x"c1"),
   746 => (x"81",x"73",x"49",x"bf"),
   747 => (x"97",x"c7",x"d4",x"c1"),
   748 => (x"32",x"c8",x"4a",x"bf"),
   749 => (x"80",x"71",x"48",x"72"),
   750 => (x"58",x"d0",x"dc",x"c1"),
   751 => (x"97",x"c8",x"d4",x"c1"),
   752 => (x"dc",x"c1",x"48",x"bf"),
   753 => (x"dc",x"c1",x"58",x"e4"),
   754 => (x"c2",x"02",x"bf",x"c0"),
   755 => (x"1e",x"c8",x"87",x"da"),
   756 => (x"1e",x"ff",x"c0",x"c1"),
   757 => (x"1e",x"ca",x"d5",x"c1"),
   758 => (x"cc",x"87",x"c1",x"f6"),
   759 => (x"02",x"98",x"70",x"86"),
   760 => (x"c0",x"87",x"c5",x"c0"),
   761 => (x"87",x"d1",x"c3",x"48"),
   762 => (x"bf",x"f8",x"db",x"c1"),
   763 => (x"c4",x"48",x"72",x"4a"),
   764 => (x"e8",x"dc",x"c1",x"30"),
   765 => (x"e0",x"dc",x"c1",x"58"),
   766 => (x"dd",x"d4",x"c1",x"5a"),
   767 => (x"c8",x"49",x"bf",x"97"),
   768 => (x"dc",x"d4",x"c1",x"31"),
   769 => (x"73",x"4b",x"bf",x"97"),
   770 => (x"de",x"d4",x"c1",x"81"),
   771 => (x"d0",x"4b",x"bf",x"97"),
   772 => (x"c1",x"81",x"73",x"33"),
   773 => (x"bf",x"97",x"df",x"d4"),
   774 => (x"73",x"33",x"d8",x"4b"),
   775 => (x"ec",x"dc",x"c1",x"81"),
   776 => (x"e0",x"dc",x"c1",x"59"),
   777 => (x"dc",x"c1",x"91",x"bf"),
   778 => (x"c1",x"81",x"bf",x"cc"),
   779 => (x"c1",x"59",x"d4",x"dc"),
   780 => (x"bf",x"97",x"e5",x"d4"),
   781 => (x"c1",x"33",x"c8",x"4b"),
   782 => (x"bf",x"97",x"e4",x"d4"),
   783 => (x"c1",x"83",x"74",x"4c"),
   784 => (x"bf",x"97",x"e6",x"d4"),
   785 => (x"74",x"34",x"d0",x"4c"),
   786 => (x"e7",x"d4",x"c1",x"83"),
   787 => (x"cf",x"4c",x"bf",x"97"),
   788 => (x"74",x"34",x"d8",x"9c"),
   789 => (x"d8",x"dc",x"c1",x"83"),
   790 => (x"73",x"8b",x"c2",x"5b"),
   791 => (x"71",x"48",x"72",x"92"),
   792 => (x"dc",x"dc",x"c1",x"80"),
   793 => (x"87",x"cf",x"c1",x"58"),
   794 => (x"97",x"ca",x"d4",x"c1"),
   795 => (x"31",x"c8",x"49",x"bf"),
   796 => (x"97",x"c9",x"d4",x"c1"),
   797 => (x"81",x"72",x"4a",x"bf"),
   798 => (x"59",x"e8",x"dc",x"c1"),
   799 => (x"ff",x"c7",x"31",x"c5"),
   800 => (x"c1",x"29",x"c9",x"81"),
   801 => (x"c1",x"59",x"e0",x"dc"),
   802 => (x"bf",x"97",x"cf",x"d4"),
   803 => (x"c1",x"32",x"c8",x"4a"),
   804 => (x"bf",x"97",x"ce",x"d4"),
   805 => (x"c1",x"82",x"73",x"4b"),
   806 => (x"c1",x"5a",x"ec",x"dc"),
   807 => (x"92",x"bf",x"e0",x"dc"),
   808 => (x"bf",x"cc",x"dc",x"c1"),
   809 => (x"dc",x"dc",x"c1",x"82"),
   810 => (x"d4",x"dc",x"c1",x"5a"),
   811 => (x"72",x"78",x"c0",x"48"),
   812 => (x"c1",x"80",x"71",x"48"),
   813 => (x"c1",x"58",x"d4",x"dc"),
   814 => (x"87",x"ea",x"f3",x"48"),
   815 => (x"5c",x"5b",x"5e",x"0e"),
   816 => (x"c0",x"dc",x"c1",x"0e"),
   817 => (x"cf",x"c0",x"02",x"bf"),
   818 => (x"4a",x"66",x"cc",x"87"),
   819 => (x"cc",x"2a",x"b7",x"c7"),
   820 => (x"ff",x"c1",x"4b",x"66"),
   821 => (x"87",x"cc",x"c0",x"9b"),
   822 => (x"c8",x"4a",x"66",x"cc"),
   823 => (x"66",x"cc",x"2a",x"b7"),
   824 => (x"9b",x"ff",x"c3",x"4b"),
   825 => (x"1e",x"f8",x"d3",x"c1"),
   826 => (x"bf",x"cc",x"dc",x"c1"),
   827 => (x"71",x"81",x"72",x"49"),
   828 => (x"87",x"f5",x"e8",x"1e"),
   829 => (x"98",x"70",x"86",x"c8"),
   830 => (x"87",x"c5",x"c0",x"05"),
   831 => (x"ea",x"c0",x"48",x"c0"),
   832 => (x"c0",x"dc",x"c1",x"87"),
   833 => (x"d4",x"c0",x"02",x"bf"),
   834 => (x"c4",x"49",x"73",x"87"),
   835 => (x"d3",x"c1",x"91",x"b7"),
   836 => (x"4c",x"69",x"81",x"f8"),
   837 => (x"ff",x"ff",x"ff",x"cf"),
   838 => (x"cc",x"c0",x"9c",x"ff"),
   839 => (x"c2",x"49",x"73",x"87"),
   840 => (x"d3",x"c1",x"91",x"b7"),
   841 => (x"69",x"9f",x"81",x"f8"),
   842 => (x"f1",x"48",x"74",x"4c"),
   843 => (x"5e",x"0e",x"87",x"fa"),
   844 => (x"0e",x"5d",x"5c",x"5b"),
   845 => (x"4b",x"c0",x"86",x"f4"),
   846 => (x"dc",x"c1",x"48",x"76"),
   847 => (x"c4",x"78",x"bf",x"d4"),
   848 => (x"d8",x"dc",x"c1",x"80"),
   849 => (x"dc",x"c1",x"78",x"bf"),
   850 => (x"c0",x"02",x"bf",x"c0"),
   851 => (x"db",x"c1",x"87",x"ca"),
   852 => (x"c4",x"49",x"bf",x"f8"),
   853 => (x"87",x"c7",x"c0",x"31"),
   854 => (x"bf",x"dc",x"dc",x"c1"),
   855 => (x"cc",x"31",x"c4",x"49"),
   856 => (x"4d",x"c0",x"59",x"a6"),
   857 => (x"c0",x"48",x"66",x"c8"),
   858 => (x"f5",x"c2",x"06",x"a8"),
   859 => (x"cf",x"49",x"75",x"87"),
   860 => (x"05",x"99",x"71",x"99"),
   861 => (x"c1",x"87",x"db",x"c0"),
   862 => (x"c8",x"1e",x"f8",x"d3"),
   863 => (x"c1",x"48",x"49",x"66"),
   864 => (x"58",x"a6",x"cc",x"80"),
   865 => (x"e0",x"e6",x"1e",x"71"),
   866 => (x"c1",x"86",x"c8",x"87"),
   867 => (x"c0",x"4b",x"f8",x"d3"),
   868 => (x"e0",x"c0",x"87",x"c3"),
   869 => (x"49",x"6b",x"97",x"83"),
   870 => (x"c1",x"02",x"99",x"71"),
   871 => (x"6b",x"97",x"87",x"fb"),
   872 => (x"a9",x"e5",x"c3",x"49"),
   873 => (x"87",x"f1",x"c1",x"02"),
   874 => (x"81",x"cb",x"49",x"73"),
   875 => (x"d8",x"49",x"69",x"97"),
   876 => (x"05",x"99",x"71",x"99"),
   877 => (x"73",x"87",x"e2",x"c1"),
   878 => (x"d9",x"ca",x"ff",x"1e"),
   879 => (x"cb",x"86",x"c4",x"87"),
   880 => (x"66",x"e4",x"c0",x"1e"),
   881 => (x"ee",x"1e",x"73",x"1e"),
   882 => (x"86",x"cc",x"87",x"d2"),
   883 => (x"c1",x"05",x"98",x"70"),
   884 => (x"4a",x"73",x"87",x"c7"),
   885 => (x"66",x"dc",x"82",x"dc"),
   886 => (x"6a",x"81",x"c4",x"49"),
   887 => (x"da",x"4a",x"73",x"79"),
   888 => (x"49",x"66",x"dc",x"82"),
   889 => (x"6a",x"9f",x"81",x"c8"),
   890 => (x"71",x"79",x"70",x"48"),
   891 => (x"c0",x"dc",x"c1",x"4c"),
   892 => (x"d2",x"c0",x"02",x"bf"),
   893 => (x"d4",x"49",x"73",x"87"),
   894 => (x"49",x"69",x"9f",x"81"),
   895 => (x"99",x"ff",x"ff",x"c0"),
   896 => (x"32",x"d0",x"4a",x"71"),
   897 => (x"c0",x"87",x"c2",x"c0"),
   898 => (x"6c",x"48",x"72",x"4a"),
   899 => (x"dc",x"7c",x"70",x"80"),
   900 => (x"78",x"c0",x"48",x"66"),
   901 => (x"c0",x"c1",x"48",x"c1"),
   902 => (x"c8",x"85",x"c1",x"87"),
   903 => (x"fd",x"04",x"ad",x"66"),
   904 => (x"dc",x"c1",x"87",x"cb"),
   905 => (x"c0",x"02",x"bf",x"c0"),
   906 => (x"1e",x"6e",x"87",x"ed"),
   907 => (x"c4",x"87",x"cd",x"fa"),
   908 => (x"58",x"a6",x"c4",x"86"),
   909 => (x"ff",x"cf",x"49",x"6e"),
   910 => (x"99",x"f8",x"ff",x"ff"),
   911 => (x"d6",x"c0",x"02",x"a9"),
   912 => (x"c2",x"49",x"6e",x"87"),
   913 => (x"f8",x"db",x"c1",x"89"),
   914 => (x"dc",x"c1",x"91",x"bf"),
   915 => (x"71",x"48",x"bf",x"d0"),
   916 => (x"58",x"a6",x"c8",x"80"),
   917 => (x"c0",x"87",x"cb",x"fc"),
   918 => (x"ed",x"8e",x"f4",x"48"),
   919 => (x"5e",x"0e",x"87",x"c8"),
   920 => (x"66",x"c8",x"0e",x"5b"),
   921 => (x"81",x"c1",x"49",x"bf"),
   922 => (x"79",x"09",x"66",x"c8"),
   923 => (x"fc",x"db",x"c1",x"09"),
   924 => (x"99",x"71",x"99",x"bf"),
   925 => (x"87",x"d0",x"c0",x"05"),
   926 => (x"c8",x"4b",x"66",x"c8"),
   927 => (x"f8",x"1e",x"6b",x"83"),
   928 => (x"86",x"c4",x"87",x"fa"),
   929 => (x"7b",x"71",x"49",x"70"),
   930 => (x"dd",x"ec",x"48",x"c1"),
   931 => (x"0e",x"5e",x"0e",x"87"),
   932 => (x"bf",x"d0",x"dc",x"c1"),
   933 => (x"4a",x"66",x"c4",x"49"),
   934 => (x"4a",x"6a",x"82",x"c8"),
   935 => (x"db",x"c1",x"8a",x"c2"),
   936 => (x"72",x"92",x"bf",x"f8"),
   937 => (x"fc",x"db",x"c1",x"81"),
   938 => (x"66",x"c4",x"4a",x"bf"),
   939 => (x"81",x"72",x"9a",x"bf"),
   940 => (x"71",x"1e",x"66",x"c8"),
   941 => (x"87",x"f1",x"e1",x"1e"),
   942 => (x"98",x"70",x"86",x"c8"),
   943 => (x"87",x"c5",x"c0",x"05"),
   944 => (x"c2",x"c0",x"48",x"c0"),
   945 => (x"eb",x"48",x"c1",x"87"),
   946 => (x"5e",x"0e",x"87",x"e2"),
   947 => (x"cc",x"0e",x"5c",x"5b"),
   948 => (x"dc",x"c1",x"1e",x"66"),
   949 => (x"d5",x"f9",x"1e",x"f0"),
   950 => (x"70",x"86",x"c8",x"87"),
   951 => (x"d4",x"c1",x"02",x"98"),
   952 => (x"f4",x"dc",x"c1",x"87"),
   953 => (x"ff",x"c7",x"49",x"bf"),
   954 => (x"71",x"29",x"c9",x"81"),
   955 => (x"c0",x"4b",x"c0",x"4c"),
   956 => (x"ff",x"1e",x"cc",x"fd"),
   957 => (x"c4",x"87",x"df",x"c5"),
   958 => (x"ac",x"b7",x"c0",x"86"),
   959 => (x"87",x"c7",x"c1",x"06"),
   960 => (x"c1",x"1e",x"66",x"d0"),
   961 => (x"fe",x"1e",x"f0",x"dc"),
   962 => (x"86",x"c8",x"87",x"c3"),
   963 => (x"c0",x"05",x"98",x"70"),
   964 => (x"48",x"c0",x"87",x"c5"),
   965 => (x"c1",x"87",x"f2",x"c0"),
   966 => (x"fd",x"1e",x"f0",x"dc"),
   967 => (x"86",x"c4",x"87",x"c0"),
   968 => (x"c8",x"48",x"66",x"d0"),
   969 => (x"a6",x"d4",x"80",x"c0"),
   970 => (x"74",x"83",x"c1",x"58"),
   971 => (x"ff",x"04",x"ab",x"b7"),
   972 => (x"d2",x"c0",x"87",x"ce"),
   973 => (x"1e",x"66",x"cc",x"87"),
   974 => (x"1e",x"e5",x"fd",x"c0"),
   975 => (x"87",x"c7",x"c5",x"ff"),
   976 => (x"48",x"c0",x"86",x"c8"),
   977 => (x"c1",x"87",x"c2",x"c0"),
   978 => (x"87",x"dc",x"e9",x"48"),
   979 => (x"6e",x"65",x"70",x"4f"),
   980 => (x"66",x"20",x"64",x"65"),
   981 => (x"2c",x"65",x"6c",x"69"),
   982 => (x"61",x"6f",x"6c",x"20"),
   983 => (x"67",x"6e",x"69",x"64"),
   984 => (x"0a",x"2e",x"2e",x"2e"),
   985 => (x"6e",x"61",x"43",x"00"),
   986 => (x"6f",x"20",x"74",x"27"),
   987 => (x"20",x"6e",x"65",x"70"),
   988 => (x"00",x"0a",x"73",x"25"),
   989 => (x"64",x"61",x"65",x"52"),
   990 => (x"20",x"66",x"6f",x"20"),
   991 => (x"20",x"52",x"42",x"4d"),
   992 => (x"6c",x"69",x"61",x"66"),
   993 => (x"00",x"0a",x"64",x"65"),
   994 => (x"70",x"20",x"6f",x"4e"),
   995 => (x"69",x"74",x"72",x"61"),
   996 => (x"6e",x"6f",x"69",x"74"),
   997 => (x"67",x"69",x"73",x"20"),
   998 => (x"75",x"74",x"61",x"6e"),
   999 => (x"66",x"20",x"65",x"72"),
  1000 => (x"64",x"6e",x"75",x"6f"),
  1001 => (x"42",x"4d",x"00",x"0a"),
  1002 => (x"7a",x"69",x"73",x"52"),
  1003 => (x"25",x"20",x"3a",x"65"),
  1004 => (x"70",x"20",x"2c",x"64"),
  1005 => (x"69",x"74",x"72",x"61"),
  1006 => (x"6e",x"6f",x"69",x"74"),
  1007 => (x"65",x"7a",x"69",x"73"),
  1008 => (x"64",x"25",x"20",x"3a"),
  1009 => (x"66",x"6f",x"20",x"2c"),
  1010 => (x"74",x"65",x"73",x"66"),
  1011 => (x"20",x"66",x"6f",x"20"),
  1012 => (x"3a",x"67",x"69",x"73"),
  1013 => (x"2c",x"64",x"25",x"20"),
  1014 => (x"67",x"69",x"73",x"20"),
  1015 => (x"25",x"78",x"30",x"20"),
  1016 => (x"52",x"00",x"0a",x"78"),
  1017 => (x"69",x"64",x"61",x"65"),
  1018 => (x"62",x"20",x"67",x"6e"),
  1019 => (x"20",x"74",x"6f",x"6f"),
  1020 => (x"74",x"63",x"65",x"73"),
  1021 => (x"25",x"20",x"72",x"6f"),
  1022 => (x"52",x"00",x"0a",x"64"),
  1023 => (x"20",x"64",x"61",x"65"),
  1024 => (x"74",x"6f",x"6f",x"62"),
  1025 => (x"63",x"65",x"73",x"20"),
  1026 => (x"20",x"72",x"6f",x"74"),
  1027 => (x"6d",x"6f",x"72",x"66"),
  1028 => (x"72",x"69",x"66",x"20"),
  1029 => (x"70",x"20",x"74",x"73"),
  1030 => (x"69",x"74",x"72",x"61"),
  1031 => (x"6e",x"6f",x"69",x"74"),
  1032 => (x"6e",x"55",x"00",x"0a"),
  1033 => (x"70",x"70",x"75",x"73"),
  1034 => (x"65",x"74",x"72",x"6f"),
  1035 => (x"61",x"70",x"20",x"64"),
  1036 => (x"74",x"69",x"74",x"72"),
  1037 => (x"20",x"6e",x"6f",x"69"),
  1038 => (x"65",x"70",x"79",x"74"),
  1039 => (x"46",x"00",x"0d",x"21"),
  1040 => (x"32",x"33",x"54",x"41"),
  1041 => (x"00",x"20",x"20",x"20"),
  1042 => (x"64",x"61",x"65",x"52"),
  1043 => (x"20",x"67",x"6e",x"69"),
  1044 => (x"0a",x"52",x"42",x"4d"),
  1045 => (x"52",x"42",x"4d",x"00"),
  1046 => (x"63",x"75",x"73",x"20"),
  1047 => (x"73",x"73",x"65",x"63"),
  1048 => (x"6c",x"6c",x"75",x"66"),
  1049 => (x"65",x"72",x"20",x"79"),
  1050 => (x"00",x"0a",x"64",x"61"),
  1051 => (x"31",x"54",x"41",x"46"),
  1052 => (x"20",x"20",x"20",x"36"),
  1053 => (x"54",x"41",x"46",x"00"),
  1054 => (x"20",x"20",x"32",x"33"),
  1055 => (x"61",x"50",x"00",x"20"),
  1056 => (x"74",x"69",x"74",x"72"),
  1057 => (x"63",x"6e",x"6f",x"69"),
  1058 => (x"74",x"6e",x"75",x"6f"),
  1059 => (x"0a",x"64",x"25",x"20"),
  1060 => (x"6e",x"75",x"48",x"00"),
  1061 => (x"67",x"6e",x"69",x"74"),
  1062 => (x"72",x"6f",x"66",x"20"),
  1063 => (x"6c",x"69",x"66",x"20"),
  1064 => (x"73",x"79",x"73",x"65"),
  1065 => (x"0a",x"6d",x"65",x"74"),
  1066 => (x"54",x"41",x"46",x"00"),
  1067 => (x"20",x"20",x"32",x"33"),
  1068 => (x"41",x"46",x"00",x"20"),
  1069 => (x"20",x"36",x"31",x"54"),
  1070 => (x"43",x"00",x"20",x"20"),
  1071 => (x"74",x"73",x"75",x"6c"),
  1072 => (x"73",x"20",x"72",x"65"),
  1073 => (x"3a",x"65",x"7a",x"69"),
  1074 => (x"2c",x"64",x"25",x"20"),
  1075 => (x"75",x"6c",x"43",x"20"),
  1076 => (x"72",x"65",x"74",x"73"),
  1077 => (x"73",x"61",x"6d",x"20"),
  1078 => (x"25",x"20",x"2c",x"6b"),
  1079 => (x"0e",x"00",x"0a",x"64"),
  1080 => (x"66",x"c4",x"0e",x"5e"),
  1081 => (x"c3",x"29",x"d8",x"49"),
  1082 => (x"66",x"c4",x"99",x"ff"),
  1083 => (x"cf",x"2a",x"c8",x"4a"),
  1084 => (x"72",x"9a",x"c0",x"fc"),
  1085 => (x"4a",x"66",x"c4",x"b1"),
  1086 => (x"ff",x"c0",x"32",x"c8"),
  1087 => (x"9a",x"c0",x"c0",x"f0"),
  1088 => (x"66",x"c4",x"b1",x"72"),
  1089 => (x"ff",x"32",x"d8",x"4a"),
  1090 => (x"c0",x"c0",x"c0",x"c0"),
  1091 => (x"71",x"b1",x"72",x"9a"),
  1092 => (x"26",x"87",x"c6",x"48"),
  1093 => (x"26",x"4c",x"26",x"4d"),
  1094 => (x"0e",x"4f",x"26",x"4b"),
  1095 => (x"66",x"c4",x"0e",x"5e"),
  1096 => (x"c3",x"2a",x"c8",x"4a"),
  1097 => (x"ff",x"cf",x"9a",x"ff"),
  1098 => (x"66",x"c4",x"9a",x"ff"),
  1099 => (x"cf",x"31",x"c8",x"49"),
  1100 => (x"72",x"99",x"c0",x"fc"),
  1101 => (x"ff",x"ff",x"cf",x"b1"),
  1102 => (x"ff",x"48",x"71",x"99"),
  1103 => (x"5e",x"0e",x"87",x"db"),
  1104 => (x"49",x"66",x"c4",x"0e"),
  1105 => (x"ff",x"cf",x"29",x"d0"),
  1106 => (x"66",x"c4",x"99",x"ff"),
  1107 => (x"f0",x"32",x"d0",x"4a"),
  1108 => (x"72",x"9a",x"c0",x"c0"),
  1109 => (x"fe",x"48",x"71",x"b1"),
  1110 => (x"73",x"1e",x"87",x"ff"),
  1111 => (x"c0",x"c0",x"d0",x"1e"),
  1112 => (x"73",x"4b",x"c0",x"c0"),
  1113 => (x"c4",x"87",x"fe",x"0f"),
  1114 => (x"26",x"4d",x"26",x"87"),
  1115 => (x"26",x"4b",x"26",x"4c"),
  1116 => (x"66",x"c8",x"1e",x"4f"),
  1117 => (x"99",x"df",x"c3",x"49"),
  1118 => (x"c0",x"89",x"f7",x"c0"),
  1119 => (x"c3",x"03",x"a9",x"b7"),
  1120 => (x"81",x"e7",x"c0",x"87"),
  1121 => (x"c4",x"48",x"66",x"c4"),
  1122 => (x"58",x"a6",x"c8",x"30"),
  1123 => (x"71",x"48",x"66",x"c4"),
  1124 => (x"58",x"a6",x"c8",x"b0"),
  1125 => (x"ff",x"48",x"66",x"c4"),
  1126 => (x"5e",x"0e",x"87",x"d5"),
  1127 => (x"d0",x"0e",x"5c",x"5b"),
  1128 => (x"c0",x"c0",x"c0",x"c0"),
  1129 => (x"fc",x"dc",x"c1",x"4c"),
  1130 => (x"80",x"c1",x"48",x"bf"),
  1131 => (x"58",x"c0",x"dd",x"c1"),
  1132 => (x"49",x"66",x"cc",x"97"),
  1133 => (x"b9",x"81",x"c0",x"fe"),
  1134 => (x"05",x"a9",x"d3",x"c1"),
  1135 => (x"dc",x"c1",x"87",x"db"),
  1136 => (x"78",x"c0",x"48",x"fc"),
  1137 => (x"48",x"c0",x"dd",x"c1"),
  1138 => (x"dd",x"c1",x"78",x"c0"),
  1139 => (x"78",x"c0",x"48",x"c8"),
  1140 => (x"48",x"cc",x"dd",x"c1"),
  1141 => (x"fb",x"c6",x"78",x"c0"),
  1142 => (x"fc",x"dc",x"c1",x"87"),
  1143 => (x"a8",x"c1",x"48",x"bf"),
  1144 => (x"87",x"f8",x"c0",x"05"),
  1145 => (x"49",x"66",x"cc",x"97"),
  1146 => (x"b9",x"81",x"c0",x"fe"),
  1147 => (x"dd",x"c1",x"1e",x"71"),
  1148 => (x"fd",x"1e",x"bf",x"cc"),
  1149 => (x"86",x"c8",x"87",x"fb"),
  1150 => (x"58",x"d0",x"dd",x"c1"),
  1151 => (x"bf",x"cc",x"dd",x"c1"),
  1152 => (x"aa",x"b7",x"c3",x"4a"),
  1153 => (x"ca",x"87",x"c6",x"06"),
  1154 => (x"70",x"88",x"72",x"48"),
  1155 => (x"c1",x"49",x"72",x"4a"),
  1156 => (x"c1",x"48",x"71",x"81"),
  1157 => (x"c8",x"dd",x"c1",x"30"),
  1158 => (x"87",x"f8",x"c5",x"58"),
  1159 => (x"bf",x"cc",x"dd",x"c1"),
  1160 => (x"a8",x"b7",x"c9",x"48"),
  1161 => (x"87",x"ec",x"c5",x"01"),
  1162 => (x"bf",x"cc",x"dd",x"c1"),
  1163 => (x"a8",x"b7",x"c0",x"48"),
  1164 => (x"87",x"e0",x"c5",x"06"),
  1165 => (x"bf",x"fc",x"dc",x"c1"),
  1166 => (x"a8",x"b7",x"c3",x"48"),
  1167 => (x"97",x"87",x"db",x"01"),
  1168 => (x"fe",x"49",x"66",x"cc"),
  1169 => (x"71",x"b9",x"81",x"c0"),
  1170 => (x"c8",x"dd",x"c1",x"1e"),
  1171 => (x"e0",x"fc",x"1e",x"bf"),
  1172 => (x"c1",x"86",x"c8",x"87"),
  1173 => (x"c4",x"58",x"cc",x"dd"),
  1174 => (x"dd",x"c1",x"87",x"fa"),
  1175 => (x"c3",x"49",x"bf",x"c4"),
  1176 => (x"fc",x"dc",x"c1",x"81"),
  1177 => (x"04",x"a9",x"b7",x"bf"),
  1178 => (x"97",x"87",x"e1",x"c0"),
  1179 => (x"fe",x"49",x"66",x"cc"),
  1180 => (x"71",x"b9",x"81",x"c0"),
  1181 => (x"c0",x"dd",x"c1",x"1e"),
  1182 => (x"f4",x"fb",x"1e",x"bf"),
  1183 => (x"c1",x"86",x"c8",x"87"),
  1184 => (x"c1",x"58",x"c4",x"dd"),
  1185 => (x"c1",x"48",x"d0",x"dd"),
  1186 => (x"87",x"c8",x"c4",x"78"),
  1187 => (x"bf",x"cc",x"dd",x"c1"),
  1188 => (x"a8",x"b7",x"c0",x"48"),
  1189 => (x"87",x"db",x"c2",x"06"),
  1190 => (x"bf",x"cc",x"dd",x"c1"),
  1191 => (x"a8",x"b7",x"c3",x"48"),
  1192 => (x"87",x"cf",x"c2",x"01"),
  1193 => (x"bf",x"c8",x"dd",x"c1"),
  1194 => (x"81",x"31",x"c1",x"49"),
  1195 => (x"bf",x"fc",x"dc",x"c1"),
  1196 => (x"c1",x"04",x"a9",x"b7"),
  1197 => (x"cc",x"97",x"87",x"df"),
  1198 => (x"c0",x"fe",x"49",x"66"),
  1199 => (x"1e",x"71",x"b9",x"81"),
  1200 => (x"bf",x"d4",x"dd",x"c1"),
  1201 => (x"87",x"e9",x"fa",x"1e"),
  1202 => (x"dd",x"c1",x"86",x"c8"),
  1203 => (x"dd",x"c1",x"58",x"d8"),
  1204 => (x"c1",x"49",x"bf",x"d0"),
  1205 => (x"d4",x"dd",x"c1",x"89"),
  1206 => (x"a9",x"b7",x"c0",x"59"),
  1207 => (x"87",x"f4",x"c2",x"03"),
  1208 => (x"bf",x"c0",x"dd",x"c1"),
  1209 => (x"d4",x"dd",x"c1",x"49"),
  1210 => (x"c3",x"51",x"bf",x"97"),
  1211 => (x"dd",x"c1",x"98",x"ff"),
  1212 => (x"c1",x"49",x"bf",x"c0"),
  1213 => (x"c4",x"dd",x"c1",x"81"),
  1214 => (x"d8",x"dd",x"c1",x"59"),
  1215 => (x"06",x"a9",x"b7",x"bf"),
  1216 => (x"c1",x"87",x"c9",x"c0"),
  1217 => (x"c1",x"48",x"d8",x"dd"),
  1218 => (x"78",x"bf",x"c0",x"dd"),
  1219 => (x"48",x"d0",x"dd",x"c1"),
  1220 => (x"ff",x"c1",x"78",x"c1"),
  1221 => (x"d0",x"dd",x"c1",x"87"),
  1222 => (x"f7",x"c1",x"05",x"bf"),
  1223 => (x"d4",x"dd",x"c1",x"87"),
  1224 => (x"31",x"c4",x"49",x"bf"),
  1225 => (x"59",x"d8",x"dd",x"c1"),
  1226 => (x"bf",x"c0",x"dd",x"c1"),
  1227 => (x"09",x"79",x"97",x"09"),
  1228 => (x"c1",x"87",x"e1",x"c1"),
  1229 => (x"48",x"bf",x"cc",x"dd"),
  1230 => (x"04",x"a8",x"b7",x"c7"),
  1231 => (x"c0",x"87",x"d5",x"c1"),
  1232 => (x"48",x"f4",x"fe",x"4b"),
  1233 => (x"dd",x"c1",x"78",x"c1"),
  1234 => (x"74",x"1e",x"bf",x"d8"),
  1235 => (x"f1",x"d2",x"c1",x"1e"),
  1236 => (x"f2",x"f4",x"fe",x"1e"),
  1237 => (x"c1",x"86",x"cc",x"87"),
  1238 => (x"c1",x"5c",x"c4",x"dd"),
  1239 => (x"48",x"bf",x"c0",x"dd"),
  1240 => (x"bf",x"d8",x"dd",x"c1"),
  1241 => (x"c0",x"03",x"a8",x"b7"),
  1242 => (x"dd",x"c1",x"87",x"db"),
  1243 => (x"83",x"bf",x"bf",x"c0"),
  1244 => (x"bf",x"c0",x"dd",x"c1"),
  1245 => (x"c1",x"81",x"c4",x"49"),
  1246 => (x"c1",x"59",x"c4",x"dd"),
  1247 => (x"b7",x"bf",x"d8",x"dd"),
  1248 => (x"e5",x"ff",x"04",x"a9"),
  1249 => (x"c1",x"1e",x"73",x"87"),
  1250 => (x"fe",x"1e",x"d0",x"d3"),
  1251 => (x"c8",x"87",x"f8",x"f3"),
  1252 => (x"87",x"c6",x"f7",x"86"),
  1253 => (x"0e",x"87",x"d4",x"f7"),
  1254 => (x"5d",x"5c",x"5b",x"5e"),
  1255 => (x"f3",x"d1",x"c1",x"0e"),
  1256 => (x"f1",x"f2",x"fe",x"1e"),
  1257 => (x"ff",x"86",x"c4",x"87"),
  1258 => (x"70",x"87",x"fe",x"c3"),
  1259 => (x"cf",x"c0",x"02",x"98"),
  1260 => (x"f9",x"d7",x"ff",x"87"),
  1261 => (x"02",x"98",x"70",x"87"),
  1262 => (x"c1",x"87",x"c5",x"c0"),
  1263 => (x"87",x"c2",x"c0",x"49"),
  1264 => (x"4d",x"71",x"49",x"c0"),
  1265 => (x"1e",x"c9",x"d2",x"c1"),
  1266 => (x"87",x"ca",x"f2",x"fe"),
  1267 => (x"dd",x"c1",x"86",x"c4"),
  1268 => (x"78",x"c0",x"48",x"d8"),
  1269 => (x"fe",x"1e",x"ee",x"c0"),
  1270 => (x"c4",x"87",x"e1",x"f1"),
  1271 => (x"c8",x"f4",x"c3",x"86"),
  1272 => (x"c0",x"ff",x"4a",x"ff"),
  1273 => (x"49",x"74",x"4c",x"bf"),
  1274 => (x"02",x"99",x"c0",x"c8"),
  1275 => (x"74",x"87",x"cc",x"c1"),
  1276 => (x"9b",x"ff",x"c3",x"4b"),
  1277 => (x"c0",x"05",x"ab",x"db"),
  1278 => (x"9d",x"75",x"87",x"f5"),
  1279 => (x"87",x"e5",x"c0",x"02"),
  1280 => (x"c0",x"c0",x"c0",x"d0"),
  1281 => (x"d1",x"c1",x"1e",x"c0"),
  1282 => (x"fd",x"ea",x"1e",x"d7"),
  1283 => (x"70",x"86",x"c8",x"87"),
  1284 => (x"d0",x"c0",x"02",x"98"),
  1285 => (x"cb",x"d1",x"c1",x"87"),
  1286 => (x"f9",x"f0",x"fe",x"1e"),
  1287 => (x"f4",x"86",x"c4",x"87"),
  1288 => (x"ca",x"c0",x"87",x"f8"),
  1289 => (x"e3",x"d1",x"c1",x"87"),
  1290 => (x"e9",x"f0",x"fe",x"1e"),
  1291 => (x"73",x"86",x"c4",x"87"),
  1292 => (x"87",x"e6",x"f5",x"1e"),
  1293 => (x"f4",x"c3",x"86",x"c4"),
  1294 => (x"72",x"4a",x"c0",x"c9"),
  1295 => (x"71",x"8a",x"c1",x"49"),
  1296 => (x"dd",x"fe",x"05",x"99"),
  1297 => (x"87",x"cc",x"fe",x"87"),
  1298 => (x"42",x"87",x"de",x"f4"),
  1299 => (x"69",x"74",x"6f",x"6f"),
  1300 => (x"2e",x"2e",x"67",x"6e"),
  1301 => (x"42",x"00",x"0a",x"2e"),
  1302 => (x"38",x"54",x"4f",x"4f"),
  1303 => (x"42",x"20",x"32",x"33"),
  1304 => (x"53",x"00",x"4e",x"49"),
  1305 => (x"6f",x"62",x"20",x"44"),
  1306 => (x"66",x"20",x"74",x"6f"),
  1307 => (x"65",x"6c",x"69",x"61"),
  1308 => (x"49",x"00",x"0a",x"64"),
  1309 => (x"69",x"74",x"69",x"6e"),
  1310 => (x"7a",x"69",x"6c",x"61"),
  1311 => (x"20",x"67",x"6e",x"69"),
  1312 => (x"63",x"20",x"44",x"53"),
  1313 => (x"0a",x"64",x"72",x"61"),
  1314 => (x"32",x"53",x"52",x"00"),
  1315 => (x"62",x"20",x"32",x"33"),
  1316 => (x"20",x"74",x"6f",x"6f"),
  1317 => (x"72",x"70",x"20",x"2d"),
  1318 => (x"20",x"73",x"73",x"65"),
  1319 => (x"20",x"43",x"53",x"45"),
  1320 => (x"62",x"20",x"6f",x"74"),
  1321 => (x"20",x"74",x"6f",x"6f"),
  1322 => (x"6d",x"6f",x"72",x"66"),
  1323 => (x"2e",x"44",x"53",x"20"),
  1324 => (x"65",x"68",x"43",x"00"),
  1325 => (x"75",x"73",x"6b",x"63"),
  1326 => (x"6e",x"69",x"6d",x"6d"),
  1327 => (x"72",x"66",x"20",x"67"),
  1328 => (x"25",x"20",x"6d",x"6f"),
  1329 => (x"6f",x"74",x"20",x"64"),
  1330 => (x"2e",x"64",x"25",x"20"),
  1331 => (x"00",x"20",x"2e",x"2e"),
  1332 => (x"00",x"0a",x"64",x"25"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
