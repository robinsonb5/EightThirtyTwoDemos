
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"c9",x"01"),
     1 => (x"cf",x"03",x"87",x"cc"),
     2 => (x"87",x"fd",x"00",x"87"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"36",x"27",x"4f",x"00"),
     5 => (x"4f",x"00",x"00",x"00"),
     6 => (x"0e",x"1e",x"18",x"0e"),
     7 => (x"00",x"00",x"44",x"27"),
     8 => (x"48",x"26",x"0f",x"00"),
     9 => (x"08",x"26",x"80",x"ff"),
    10 => (x"c0",x"c0",x"c2",x"4f"),
    11 => (x"05",x"29",x"27",x"4e"),
    12 => (x"00",x"0f",x"00",x"00"),
    13 => (x"f0",x"c1",x"87",x"fd"),
    14 => (x"43",x"27",x"4e",x"c0"),
    15 => (x"0f",x"00",x"00",x"00"),
    16 => (x"4f",x"87",x"fd",x"00"),
    17 => (x"0e",x"1e",x"18",x"0e"),
    18 => (x"80",x"ff",x"48",x"26"),
    19 => (x"1e",x"4f",x"08",x"26"),
    20 => (x"ff",x"1e",x"1e",x"72"),
    21 => (x"48",x"6a",x"4a",x"c0"),
    22 => (x"c4",x"98",x"c0",x"c4"),
    23 => (x"02",x"6e",x"58",x"a6"),
    24 => (x"cc",x"87",x"f3",x"ff"),
    25 => (x"66",x"cc",x"7a",x"66"),
    26 => (x"4a",x"26",x"26",x"48"),
    27 => (x"5e",x"0e",x"4f",x"26"),
    28 => (x"5d",x"5c",x"5b",x"5a"),
    29 => (x"4d",x"66",x"d4",x"0e"),
    30 => (x"4b",x"15",x"4c",x"c0"),
    31 => (x"c0",x"02",x"9b",x"73"),
    32 => (x"4a",x"73",x"87",x"d6"),
    33 => (x"4f",x"27",x"1e",x"72"),
    34 => (x"0f",x"00",x"00",x"00"),
    35 => (x"84",x"c1",x"86",x"c4"),
    36 => (x"9b",x"73",x"4b",x"15"),
    37 => (x"87",x"ea",x"ff",x"05"),
    38 => (x"4d",x"26",x"48",x"74"),
    39 => (x"4b",x"26",x"4c",x"26"),
    40 => (x"4f",x"26",x"4a",x"26"),
    41 => (x"5b",x"5a",x"5e",x"0e"),
    42 => (x"1e",x"0e",x"5d",x"5c"),
    43 => (x"27",x"4d",x"66",x"d8"),
    44 => (x"00",x"00",x"16",x"40"),
    45 => (x"27",x"49",x"76",x"4b"),
    46 => (x"00",x"00",x"0e",x"68"),
    47 => (x"75",x"4c",x"c0",x"79"),
    48 => (x"a9",x"b7",x"c0",x"49"),
    49 => (x"87",x"ce",x"c0",x"03"),
    50 => (x"27",x"1e",x"ed",x"c0"),
    51 => (x"00",x"00",x"00",x"4f"),
    52 => (x"c0",x"86",x"c4",x"0f"),
    53 => (x"9d",x"75",x"8d",x"0d"),
    54 => (x"87",x"c6",x"c0",x"05"),
    55 => (x"c0",x"53",x"f0",x"c0"),
    56 => (x"9d",x"75",x"87",x"f6"),
    57 => (x"87",x"f0",x"c0",x"02"),
    58 => (x"1e",x"72",x"49",x"75"),
    59 => (x"4a",x"66",x"e4",x"c0"),
    60 => (x"00",x"04",x"c4",x"27"),
    61 => (x"4a",x"26",x"0f",x"00"),
    62 => (x"4a",x"72",x"4a",x"71"),
    63 => (x"53",x"12",x"82",x"6e"),
    64 => (x"1e",x"72",x"49",x"75"),
    65 => (x"4a",x"66",x"e4",x"c0"),
    66 => (x"00",x"04",x"c4",x"27"),
    67 => (x"4a",x"26",x"0f",x"00"),
    68 => (x"9d",x"75",x"4d",x"70"),
    69 => (x"87",x"d0",x"ff",x"05"),
    70 => (x"40",x"27",x"49",x"73"),
    71 => (x"b7",x"00",x"00",x"16"),
    72 => (x"e1",x"c0",x"02",x"a9"),
    73 => (x"dc",x"8b",x"c1",x"87"),
    74 => (x"97",x"49",x"bf",x"a6"),
    75 => (x"66",x"dc",x"51",x"6b"),
    76 => (x"c0",x"80",x"c1",x"48"),
    77 => (x"c1",x"58",x"a6",x"e0"),
    78 => (x"27",x"49",x"73",x"84"),
    79 => (x"00",x"00",x"16",x"40"),
    80 => (x"ff",x"05",x"a9",x"b7"),
    81 => (x"a6",x"dc",x"87",x"df"),
    82 => (x"51",x"c0",x"49",x"bf"),
    83 => (x"26",x"26",x"48",x"74"),
    84 => (x"26",x"4c",x"26",x"4d"),
    85 => (x"26",x"4a",x"26",x"4b"),
    86 => (x"5a",x"5e",x"0e",x"4f"),
    87 => (x"0e",x"5d",x"5c",x"5b"),
    88 => (x"76",x"4c",x"c0",x"1e"),
    89 => (x"dc",x"79",x"c0",x"49"),
    90 => (x"66",x"d8",x"4b",x"a6"),
    91 => (x"48",x"66",x"d8",x"4a"),
    92 => (x"a6",x"dc",x"80",x"c1"),
    93 => (x"d8",x"4d",x"12",x"58"),
    94 => (x"75",x"2d",x"b7",x"35"),
    95 => (x"d7",x"c4",x"02",x"9d"),
    96 => (x"c3",x"02",x"6e",x"87"),
    97 => (x"49",x"76",x"87",x"e1"),
    98 => (x"4a",x"75",x"79",x"c0"),
    99 => (x"e3",x"c1",x"49",x"75"),
   100 => (x"e5",x"c2",x"02",x"a9"),
   101 => (x"c1",x"49",x"72",x"87"),
   102 => (x"c0",x"02",x"a9",x"e4"),
   103 => (x"49",x"72",x"87",x"de"),
   104 => (x"02",x"a9",x"ec",x"c1"),
   105 => (x"72",x"87",x"cc",x"c2"),
   106 => (x"a9",x"f3",x"c1",x"49"),
   107 => (x"87",x"ea",x"c1",x"02"),
   108 => (x"f8",x"c1",x"49",x"72"),
   109 => (x"f2",x"c0",x"02",x"a9"),
   110 => (x"87",x"d3",x"c2",x"87"),
   111 => (x"90",x"27",x"1e",x"ca"),
   112 => (x"1e",x"00",x"00",x"16"),
   113 => (x"4a",x"73",x"83",x"c4"),
   114 => (x"1e",x"6a",x"8a",x"c4"),
   115 => (x"00",x"00",x"a4",x"27"),
   116 => (x"86",x"cc",x"0f",x"00"),
   117 => (x"4c",x"74",x"4a",x"70"),
   118 => (x"90",x"27",x"84",x"72"),
   119 => (x"1e",x"00",x"00",x"16"),
   120 => (x"00",x"00",x"6e",x"27"),
   121 => (x"86",x"c4",x"0f",x"00"),
   122 => (x"d0",x"87",x"d6",x"c2"),
   123 => (x"16",x"90",x"27",x"1e"),
   124 => (x"c4",x"1e",x"00",x"00"),
   125 => (x"c4",x"4a",x"73",x"83"),
   126 => (x"27",x"1e",x"6a",x"8a"),
   127 => (x"00",x"00",x"00",x"a4"),
   128 => (x"70",x"86",x"cc",x"0f"),
   129 => (x"72",x"4c",x"74",x"4a"),
   130 => (x"16",x"90",x"27",x"84"),
   131 => (x"27",x"1e",x"00",x"00"),
   132 => (x"00",x"00",x"00",x"6e"),
   133 => (x"c1",x"86",x"c4",x"0f"),
   134 => (x"83",x"c4",x"87",x"e7"),
   135 => (x"8a",x"c4",x"4a",x"73"),
   136 => (x"6e",x"27",x"1e",x"6a"),
   137 => (x"0f",x"00",x"00",x"00"),
   138 => (x"4a",x"70",x"86",x"c4"),
   139 => (x"84",x"72",x"4c",x"74"),
   140 => (x"76",x"87",x"ce",x"c1"),
   141 => (x"c1",x"79",x"c1",x"49"),
   142 => (x"83",x"c4",x"87",x"c7"),
   143 => (x"8a",x"c4",x"4a",x"73"),
   144 => (x"4f",x"27",x"1e",x"6a"),
   145 => (x"0f",x"00",x"00",x"00"),
   146 => (x"84",x"c1",x"86",x"c4"),
   147 => (x"c0",x"87",x"f2",x"c0"),
   148 => (x"4f",x"27",x"1e",x"e5"),
   149 => (x"0f",x"00",x"00",x"00"),
   150 => (x"1e",x"75",x"86",x"c4"),
   151 => (x"00",x"00",x"4f",x"27"),
   152 => (x"86",x"c4",x"0f",x"00"),
   153 => (x"75",x"87",x"da",x"c0"),
   154 => (x"a9",x"e5",x"c0",x"49"),
   155 => (x"87",x"c7",x"c0",x"05"),
   156 => (x"79",x"c1",x"49",x"76"),
   157 => (x"75",x"87",x"ca",x"c0"),
   158 => (x"00",x"4f",x"27",x"1e"),
   159 => (x"c4",x"0f",x"00",x"00"),
   160 => (x"4a",x"66",x"d8",x"86"),
   161 => (x"c1",x"48",x"66",x"d8"),
   162 => (x"58",x"a6",x"dc",x"80"),
   163 => (x"35",x"d8",x"4d",x"12"),
   164 => (x"9d",x"75",x"2d",x"b7"),
   165 => (x"87",x"e9",x"fb",x"05"),
   166 => (x"26",x"26",x"48",x"74"),
   167 => (x"26",x"4c",x"26",x"4d"),
   168 => (x"26",x"4a",x"26",x"4b"),
   169 => (x"5a",x"5e",x"0e",x"4f"),
   170 => (x"66",x"d0",x"0e",x"5b"),
   171 => (x"7b",x"66",x"cc",x"4b"),
   172 => (x"27",x"1e",x"66",x"cc"),
   173 => (x"00",x"00",x"04",x"b0"),
   174 => (x"70",x"86",x"c4",x"0f"),
   175 => (x"05",x"9a",x"72",x"4a"),
   176 => (x"c3",x"87",x"c2",x"c0"),
   177 => (x"4a",x"66",x"cc",x"7b"),
   178 => (x"c0",x"49",x"66",x"cc"),
   179 => (x"c0",x"02",x"a9",x"b7"),
   180 => (x"49",x"72",x"87",x"e7"),
   181 => (x"02",x"a9",x"b7",x"c1"),
   182 => (x"72",x"87",x"e3",x"c0"),
   183 => (x"a9",x"b7",x"c2",x"49"),
   184 => (x"87",x"f3",x"c0",x"02"),
   185 => (x"b7",x"c3",x"49",x"72"),
   186 => (x"f1",x"c0",x"02",x"a9"),
   187 => (x"c4",x"49",x"72",x"87"),
   188 => (x"c0",x"02",x"a9",x"b7"),
   189 => (x"e5",x"c0",x"87",x"e6"),
   190 => (x"c0",x"7b",x"c0",x"87"),
   191 => (x"3c",x"27",x"87",x"e0"),
   192 => (x"bf",x"00",x"00",x"18"),
   193 => (x"b7",x"e4",x"c1",x"49"),
   194 => (x"c5",x"c0",x"06",x"a9"),
   195 => (x"c0",x"7b",x"c0",x"87"),
   196 => (x"7b",x"c3",x"87",x"cc"),
   197 => (x"c1",x"87",x"c7",x"c0"),
   198 => (x"87",x"c2",x"c0",x"7b"),
   199 => (x"4b",x"26",x"7b",x"c2"),
   200 => (x"4f",x"26",x"4a",x"26"),
   201 => (x"c8",x"1e",x"72",x"1e"),
   202 => (x"82",x"c2",x"4a",x"66"),
   203 => (x"72",x"48",x"66",x"cc"),
   204 => (x"49",x"66",x"d0",x"80"),
   205 => (x"26",x"4a",x"26",x"58"),
   206 => (x"5a",x"5e",x"0e",x"4f"),
   207 => (x"0e",x"5d",x"5c",x"5b"),
   208 => (x"c5",x"4d",x"66",x"dc"),
   209 => (x"c4",x"4a",x"75",x"85"),
   210 => (x"d4",x"4a",x"72",x"92"),
   211 => (x"e0",x"c0",x"82",x"66"),
   212 => (x"4b",x"72",x"7a",x"66"),
   213 => (x"7b",x"6a",x"83",x"c4"),
   214 => (x"75",x"82",x"f8",x"c1"),
   215 => (x"75",x"4c",x"75",x"7a"),
   216 => (x"75",x"82",x"c1",x"4a"),
   217 => (x"a9",x"b7",x"72",x"49"),
   218 => (x"87",x"e3",x"c0",x"01"),
   219 => (x"c8",x"c3",x"4b",x"75"),
   220 => (x"d8",x"4b",x"73",x"93"),
   221 => (x"4a",x"74",x"83",x"66"),
   222 => (x"4a",x"72",x"92",x"c4"),
   223 => (x"7a",x"75",x"82",x"73"),
   224 => (x"4a",x"75",x"84",x"c1"),
   225 => (x"49",x"74",x"82",x"c1"),
   226 => (x"06",x"a9",x"b7",x"72"),
   227 => (x"75",x"87",x"dd",x"ff"),
   228 => (x"94",x"c8",x"c3",x"4c"),
   229 => (x"66",x"d8",x"4c",x"74"),
   230 => (x"c4",x"4a",x"75",x"84"),
   231 => (x"72",x"4b",x"74",x"92"),
   232 => (x"c1",x"48",x"6b",x"83"),
   233 => (x"66",x"d4",x"58",x"80"),
   234 => (x"c0",x"83",x"72",x"4b"),
   235 => (x"72",x"84",x"e0",x"fe"),
   236 => (x"6b",x"82",x"74",x"4a"),
   237 => (x"18",x"3c",x"27",x"7a"),
   238 => (x"c5",x"49",x"00",x"00"),
   239 => (x"26",x"4d",x"26",x"79"),
   240 => (x"26",x"4b",x"26",x"4c"),
   241 => (x"0e",x"4f",x"26",x"4a"),
   242 => (x"5c",x"5b",x"5a",x"5e"),
   243 => (x"66",x"d0",x"97",x"0e"),
   244 => (x"d8",x"4b",x"74",x"4c"),
   245 => (x"97",x"2b",x"b7",x"33"),
   246 => (x"d8",x"4a",x"66",x"d4"),
   247 => (x"73",x"2a",x"b7",x"32"),
   248 => (x"a9",x"b7",x"72",x"49"),
   249 => (x"87",x"c5",x"c0",x"02"),
   250 => (x"ca",x"c0",x"48",x"c0"),
   251 => (x"17",x"30",x"27",x"87"),
   252 => (x"74",x"49",x"00",x"00"),
   253 => (x"26",x"48",x"c1",x"51"),
   254 => (x"26",x"4b",x"26",x"4c"),
   255 => (x"0e",x"4f",x"26",x"4a"),
   256 => (x"0e",x"5b",x"5a",x"5e"),
   257 => (x"d4",x"4b",x"c2",x"1e"),
   258 => (x"82",x"c1",x"4a",x"66"),
   259 => (x"6a",x"97",x"82",x"73"),
   260 => (x"b7",x"32",x"d8",x"4a"),
   261 => (x"d4",x"1e",x"72",x"2a"),
   262 => (x"82",x"73",x"4a",x"66"),
   263 => (x"d8",x"4a",x"6a",x"97"),
   264 => (x"72",x"2a",x"b7",x"32"),
   265 => (x"03",x"c7",x"27",x"1e"),
   266 => (x"c8",x"0f",x"00",x"00"),
   267 => (x"72",x"4a",x"70",x"86"),
   268 => (x"c7",x"c0",x"05",x"9a"),
   269 => (x"c1",x"49",x"76",x"87"),
   270 => (x"83",x"c1",x"51",x"c1"),
   271 => (x"b7",x"c2",x"49",x"73"),
   272 => (x"c2",x"ff",x"06",x"a9"),
   273 => (x"4a",x"6e",x"97",x"87"),
   274 => (x"2a",x"b7",x"32",x"d8"),
   275 => (x"d7",x"c1",x"49",x"72"),
   276 => (x"c0",x"04",x"a9",x"b7"),
   277 => (x"6e",x"97",x"87",x"d3"),
   278 => (x"b7",x"32",x"d8",x"4a"),
   279 => (x"c1",x"49",x"72",x"2a"),
   280 => (x"03",x"a9",x"b7",x"da"),
   281 => (x"c7",x"87",x"c2",x"c0"),
   282 => (x"4a",x"6e",x"97",x"4b"),
   283 => (x"2a",x"b7",x"32",x"d8"),
   284 => (x"d2",x"c1",x"49",x"72"),
   285 => (x"c0",x"05",x"a9",x"b7"),
   286 => (x"48",x"c1",x"87",x"c5"),
   287 => (x"d4",x"87",x"ea",x"c0"),
   288 => (x"66",x"d4",x"1e",x"66"),
   289 => (x"05",x"0e",x"27",x"1e"),
   290 => (x"c8",x"0f",x"00",x"00"),
   291 => (x"72",x"4a",x"70",x"86"),
   292 => (x"a9",x"b7",x"c0",x"49"),
   293 => (x"87",x"cf",x"c0",x"06"),
   294 => (x"80",x"c7",x"48",x"73"),
   295 => (x"00",x"18",x"3c",x"27"),
   296 => (x"48",x"c1",x"58",x"00"),
   297 => (x"c0",x"87",x"c2",x"c0"),
   298 => (x"4b",x"26",x"26",x"48"),
   299 => (x"4f",x"26",x"4a",x"26"),
   300 => (x"49",x"66",x"c4",x"1e"),
   301 => (x"05",x"a9",x"b7",x"c2"),
   302 => (x"c1",x"87",x"c5",x"c0"),
   303 => (x"87",x"c2",x"c0",x"48"),
   304 => (x"4f",x"26",x"48",x"c0"),
   305 => (x"72",x"1e",x"73",x"1e"),
   306 => (x"87",x"d9",x"02",x"9a"),
   307 => (x"4b",x"c1",x"48",x"c0"),
   308 => (x"82",x"01",x"a9",x"72"),
   309 => (x"87",x"f8",x"83",x"73"),
   310 => (x"89",x"03",x"a9",x"72"),
   311 => (x"c1",x"07",x"80",x"73"),
   312 => (x"f3",x"05",x"2b",x"2a"),
   313 => (x"26",x"4b",x"26",x"87"),
   314 => (x"1e",x"75",x"1e",x"4f"),
   315 => (x"a1",x"71",x"4d",x"c0"),
   316 => (x"c1",x"b9",x"ff",x"04"),
   317 => (x"72",x"07",x"bd",x"81"),
   318 => (x"ba",x"ff",x"04",x"a2"),
   319 => (x"07",x"bd",x"82",x"c1"),
   320 => (x"9d",x"75",x"87",x"c2"),
   321 => (x"c1",x"b8",x"ff",x"05"),
   322 => (x"4d",x"25",x"07",x"80"),
   323 => (x"c4",x"1e",x"4f",x"26"),
   324 => (x"66",x"c8",x"49",x"66"),
   325 => (x"11",x"48",x"12",x"4a"),
   326 => (x"88",x"87",x"c4",x"02"),
   327 => (x"26",x"87",x"f6",x"02"),
   328 => (x"c8",x"ff",x"1e",x"4f"),
   329 => (x"26",x"48",x"68",x"48"),
   330 => (x"5a",x"5e",x"0e",x"4f"),
   331 => (x"0e",x"5d",x"5c",x"5b"),
   332 => (x"66",x"c4",x"8e",x"d0"),
   333 => (x"17",x"38",x"27",x"4c"),
   334 => (x"27",x"49",x"00",x"00"),
   335 => (x"00",x"00",x"17",x"40"),
   336 => (x"16",x"b8",x"27",x"79"),
   337 => (x"27",x"49",x"00",x"00"),
   338 => (x"00",x"00",x"17",x"00"),
   339 => (x"17",x"00",x"27",x"79"),
   340 => (x"27",x"49",x"00",x"00"),
   341 => (x"00",x"00",x"17",x"40"),
   342 => (x"17",x"04",x"27",x"79"),
   343 => (x"c0",x"49",x"00",x"00"),
   344 => (x"17",x"08",x"27",x"79"),
   345 => (x"c2",x"49",x"00",x"00"),
   346 => (x"17",x"0c",x"27",x"79"),
   347 => (x"c0",x"49",x"00",x"00"),
   348 => (x"10",x"27",x"79",x"e8"),
   349 => (x"49",x"00",x"00",x"17"),
   350 => (x"00",x"0f",x"f2",x"27"),
   351 => (x"1e",x"72",x"48",x"00"),
   352 => (x"10",x"4a",x"a1",x"df"),
   353 => (x"05",x"aa",x"71",x"51"),
   354 => (x"4a",x"26",x"87",x"f9"),
   355 => (x"00",x"16",x"c0",x"27"),
   356 => (x"11",x"27",x"49",x"00"),
   357 => (x"48",x"00",x"00",x"10"),
   358 => (x"a1",x"df",x"1e",x"72"),
   359 => (x"71",x"51",x"10",x"4a"),
   360 => (x"87",x"f9",x"05",x"aa"),
   361 => (x"ac",x"27",x"4a",x"26"),
   362 => (x"49",x"00",x"00",x"1e"),
   363 => (x"30",x"27",x"79",x"ca"),
   364 => (x"1e",x"00",x"00",x"10"),
   365 => (x"00",x"01",x"59",x"27"),
   366 => (x"86",x"c4",x"0f",x"00"),
   367 => (x"00",x"10",x"32",x"27"),
   368 => (x"59",x"27",x"1e",x"00"),
   369 => (x"0f",x"00",x"00",x"01"),
   370 => (x"62",x"27",x"86",x"c4"),
   371 => (x"1e",x"00",x"00",x"10"),
   372 => (x"00",x"01",x"59",x"27"),
   373 => (x"86",x"c4",x"0f",x"00"),
   374 => (x"00",x"16",x"34",x"27"),
   375 => (x"c0",x"02",x"bf",x"00"),
   376 => (x"79",x"27",x"87",x"df"),
   377 => (x"1e",x"00",x"00",x"0e"),
   378 => (x"00",x"01",x"59",x"27"),
   379 => (x"86",x"c4",x"0f",x"00"),
   380 => (x"00",x"0e",x"a5",x"27"),
   381 => (x"59",x"27",x"1e",x"00"),
   382 => (x"0f",x"00",x"00",x"01"),
   383 => (x"dc",x"c0",x"86",x"c4"),
   384 => (x"0e",x"a7",x"27",x"87"),
   385 => (x"27",x"1e",x"00",x"00"),
   386 => (x"00",x"00",x"01",x"59"),
   387 => (x"27",x"86",x"c4",x"0f"),
   388 => (x"00",x"00",x"0e",x"d6"),
   389 => (x"01",x"59",x"27",x"1e"),
   390 => (x"c4",x"0f",x"00",x"00"),
   391 => (x"16",x"38",x"27",x"86"),
   392 => (x"1e",x"bf",x"00",x"00"),
   393 => (x"00",x"10",x"64",x"27"),
   394 => (x"59",x"27",x"1e",x"00"),
   395 => (x"0f",x"00",x"00",x"01"),
   396 => (x"21",x"27",x"86",x"c8"),
   397 => (x"0f",x"00",x"00",x"05"),
   398 => (x"b4",x"27",x"86",x"c0"),
   399 => (x"58",x"00",x"00",x"16"),
   400 => (x"00",x"16",x"b4",x"27"),
   401 => (x"27",x"1e",x"bf",x"00"),
   402 => (x"00",x"00",x"10",x"91"),
   403 => (x"01",x"59",x"27",x"1e"),
   404 => (x"c8",x"0f",x"00",x"00"),
   405 => (x"05",x"21",x"27",x"86"),
   406 => (x"c0",x"0f",x"00",x"00"),
   407 => (x"16",x"b4",x"27",x"86"),
   408 => (x"c1",x"58",x"00",x"00"),
   409 => (x"16",x"38",x"27",x"4d"),
   410 => (x"49",x"bf",x"00",x"00"),
   411 => (x"06",x"a9",x"b7",x"c0"),
   412 => (x"27",x"87",x"d3",x"c6"),
   413 => (x"00",x"00",x"0e",x"53"),
   414 => (x"27",x"86",x"c0",x"0f"),
   415 => (x"00",x"00",x"0e",x"17"),
   416 => (x"76",x"86",x"c0",x"0f"),
   417 => (x"c3",x"79",x"c2",x"49"),
   418 => (x"16",x"e0",x"27",x"4c"),
   419 => (x"27",x"49",x"00",x"00"),
   420 => (x"00",x"00",x"0e",x"f7"),
   421 => (x"df",x"1e",x"72",x"48"),
   422 => (x"51",x"10",x"4a",x"a1"),
   423 => (x"f9",x"05",x"aa",x"71"),
   424 => (x"c8",x"4a",x"26",x"87"),
   425 => (x"79",x"c1",x"49",x"a6"),
   426 => (x"00",x"16",x"e0",x"27"),
   427 => (x"c0",x"27",x"1e",x"00"),
   428 => (x"1e",x"00",x"00",x"16"),
   429 => (x"00",x"03",x"ff",x"27"),
   430 => (x"86",x"c8",x"0f",x"00"),
   431 => (x"9a",x"72",x"4a",x"70"),
   432 => (x"87",x"c5",x"c0",x"05"),
   433 => (x"c2",x"c0",x"4a",x"c1"),
   434 => (x"27",x"4a",x"c0",x"87"),
   435 => (x"00",x"00",x"18",x"40"),
   436 => (x"6e",x"79",x"72",x"49"),
   437 => (x"a9",x"b7",x"74",x"49"),
   438 => (x"87",x"ed",x"c0",x"03"),
   439 => (x"92",x"c5",x"4a",x"6e"),
   440 => (x"88",x"74",x"48",x"72"),
   441 => (x"cc",x"58",x"a6",x"d0"),
   442 => (x"1e",x"72",x"4a",x"a6"),
   443 => (x"66",x"c8",x"1e",x"74"),
   444 => (x"03",x"24",x"27",x"1e"),
   445 => (x"cc",x"0f",x"00",x"00"),
   446 => (x"c1",x"48",x"6e",x"86"),
   447 => (x"58",x"a6",x"c4",x"80"),
   448 => (x"b7",x"74",x"49",x"6e"),
   449 => (x"d3",x"ff",x"04",x"a9"),
   450 => (x"1e",x"66",x"cc",x"87"),
   451 => (x"27",x"1e",x"66",x"c4"),
   452 => (x"00",x"00",x"18",x"50"),
   453 => (x"17",x"70",x"27",x"1e"),
   454 => (x"27",x"1e",x"00",x"00"),
   455 => (x"00",x"00",x"03",x"39"),
   456 => (x"27",x"86",x"d0",x"0f"),
   457 => (x"00",x"00",x"16",x"b8"),
   458 => (x"ff",x"27",x"1e",x"bf"),
   459 => (x"0f",x"00",x"00",x"0c"),
   460 => (x"a6",x"c4",x"86",x"c4"),
   461 => (x"51",x"c1",x"c1",x"49"),
   462 => (x"00",x"18",x"38",x"27"),
   463 => (x"4a",x"bf",x"97",x"00"),
   464 => (x"2a",x"b7",x"32",x"d8"),
   465 => (x"c1",x"c1",x"49",x"72"),
   466 => (x"c1",x"04",x"a9",x"b7"),
   467 => (x"c3",x"c1",x"87",x"fb"),
   468 => (x"66",x"c8",x"97",x"1e"),
   469 => (x"b7",x"32",x"d8",x"4a"),
   470 => (x"27",x"1e",x"72",x"2a"),
   471 => (x"00",x"00",x"03",x"c7"),
   472 => (x"70",x"86",x"c8",x"0f"),
   473 => (x"49",x"66",x"c8",x"4a"),
   474 => (x"05",x"a9",x"b7",x"72"),
   475 => (x"c8",x"87",x"f3",x"c0"),
   476 => (x"1e",x"72",x"4a",x"a6"),
   477 => (x"a5",x"27",x"1e",x"c0"),
   478 => (x"0f",x"00",x"00",x"02"),
   479 => (x"e0",x"27",x"86",x"c8"),
   480 => (x"49",x"00",x"00",x"16"),
   481 => (x"00",x"0e",x"d8",x"27"),
   482 => (x"1e",x"72",x"48",x"00"),
   483 => (x"10",x"4a",x"a1",x"df"),
   484 => (x"05",x"aa",x"71",x"51"),
   485 => (x"4a",x"26",x"87",x"f9"),
   486 => (x"3c",x"27",x"4c",x"75"),
   487 => (x"49",x"00",x"00",x"18"),
   488 => (x"c4",x"97",x"79",x"75"),
   489 => (x"80",x"c1",x"48",x"66"),
   490 => (x"50",x"08",x"a6",x"c4"),
   491 => (x"4b",x"66",x"c4",x"97"),
   492 => (x"2b",x"b7",x"33",x"d8"),
   493 => (x"00",x"18",x"38",x"27"),
   494 => (x"4a",x"bf",x"97",x"00"),
   495 => (x"2a",x"b7",x"32",x"d8"),
   496 => (x"b7",x"72",x"49",x"73"),
   497 => (x"c5",x"fe",x"06",x"a9"),
   498 => (x"74",x"94",x"6e",x"87"),
   499 => (x"d0",x"1e",x"72",x"49"),
   500 => (x"c4",x"27",x"4a",x"66"),
   501 => (x"0f",x"00",x"00",x"04"),
   502 => (x"48",x"70",x"4a",x"26"),
   503 => (x"74",x"58",x"a6",x"c4"),
   504 => (x"8a",x"66",x"cc",x"4a"),
   505 => (x"4c",x"72",x"92",x"c7"),
   506 => (x"4a",x"76",x"8c",x"6e"),
   507 => (x"9d",x"27",x"1e",x"72"),
   508 => (x"0f",x"00",x"00",x"0d"),
   509 => (x"85",x"c1",x"86",x"c4"),
   510 => (x"38",x"27",x"49",x"75"),
   511 => (x"bf",x"00",x"00",x"16"),
   512 => (x"f9",x"06",x"a9",x"b7"),
   513 => (x"21",x"27",x"87",x"ed"),
   514 => (x"0f",x"00",x"00",x"05"),
   515 => (x"34",x"27",x"86",x"c0"),
   516 => (x"58",x"00",x"00",x"17"),
   517 => (x"00",x"17",x"34",x"27"),
   518 => (x"27",x"1e",x"bf",x"00"),
   519 => (x"00",x"00",x"10",x"a1"),
   520 => (x"01",x"59",x"27",x"1e"),
   521 => (x"c8",x"0f",x"00",x"00"),
   522 => (x"10",x"af",x"27",x"86"),
   523 => (x"27",x"1e",x"00",x"00"),
   524 => (x"00",x"00",x"01",x"59"),
   525 => (x"27",x"86",x"c4",x"0f"),
   526 => (x"00",x"00",x"10",x"bf"),
   527 => (x"01",x"59",x"27",x"1e"),
   528 => (x"c4",x"0f",x"00",x"00"),
   529 => (x"10",x"c1",x"27",x"86"),
   530 => (x"27",x"1e",x"00",x"00"),
   531 => (x"00",x"00",x"01",x"59"),
   532 => (x"27",x"86",x"c4",x"0f"),
   533 => (x"00",x"00",x"10",x"f7"),
   534 => (x"01",x"59",x"27",x"1e"),
   535 => (x"c4",x"0f",x"00",x"00"),
   536 => (x"18",x"3c",x"27",x"86"),
   537 => (x"1e",x"bf",x"00",x"00"),
   538 => (x"00",x"10",x"f9",x"27"),
   539 => (x"59",x"27",x"1e",x"00"),
   540 => (x"0f",x"00",x"00",x"01"),
   541 => (x"1e",x"c5",x"86",x"c8"),
   542 => (x"00",x"11",x"12",x"27"),
   543 => (x"59",x"27",x"1e",x"00"),
   544 => (x"0f",x"00",x"00",x"01"),
   545 => (x"40",x"27",x"86",x"c8"),
   546 => (x"bf",x"00",x"00",x"18"),
   547 => (x"11",x"2b",x"27",x"1e"),
   548 => (x"27",x"1e",x"00",x"00"),
   549 => (x"00",x"00",x"01",x"59"),
   550 => (x"c1",x"86",x"c8",x"0f"),
   551 => (x"11",x"44",x"27",x"1e"),
   552 => (x"27",x"1e",x"00",x"00"),
   553 => (x"00",x"00",x"01",x"59"),
   554 => (x"27",x"86",x"c8",x"0f"),
   555 => (x"00",x"00",x"17",x"30"),
   556 => (x"d8",x"4a",x"bf",x"97"),
   557 => (x"72",x"2a",x"b7",x"32"),
   558 => (x"11",x"5d",x"27",x"1e"),
   559 => (x"27",x"1e",x"00",x"00"),
   560 => (x"00",x"00",x"01",x"59"),
   561 => (x"c1",x"86",x"c8",x"0f"),
   562 => (x"76",x"27",x"1e",x"c1"),
   563 => (x"1e",x"00",x"00",x"11"),
   564 => (x"00",x"01",x"59",x"27"),
   565 => (x"86",x"c8",x"0f",x"00"),
   566 => (x"00",x"18",x"38",x"27"),
   567 => (x"4a",x"bf",x"97",x"00"),
   568 => (x"2a",x"b7",x"32",x"d8"),
   569 => (x"8f",x"27",x"1e",x"72"),
   570 => (x"1e",x"00",x"00",x"11"),
   571 => (x"00",x"01",x"59",x"27"),
   572 => (x"86",x"c8",x"0f",x"00"),
   573 => (x"27",x"1e",x"c2",x"c1"),
   574 => (x"00",x"00",x"11",x"a8"),
   575 => (x"01",x"59",x"27",x"1e"),
   576 => (x"c8",x"0f",x"00",x"00"),
   577 => (x"17",x"90",x"27",x"86"),
   578 => (x"1e",x"bf",x"00",x"00"),
   579 => (x"00",x"11",x"c1",x"27"),
   580 => (x"59",x"27",x"1e",x"00"),
   581 => (x"0f",x"00",x"00",x"01"),
   582 => (x"1e",x"c7",x"86",x"c8"),
   583 => (x"00",x"11",x"da",x"27"),
   584 => (x"59",x"27",x"1e",x"00"),
   585 => (x"0f",x"00",x"00",x"01"),
   586 => (x"ac",x"27",x"86",x"c8"),
   587 => (x"bf",x"00",x"00",x"1e"),
   588 => (x"11",x"f3",x"27",x"1e"),
   589 => (x"27",x"1e",x"00",x"00"),
   590 => (x"00",x"00",x"01",x"59"),
   591 => (x"27",x"86",x"c8",x"0f"),
   592 => (x"00",x"00",x"12",x"0c"),
   593 => (x"01",x"59",x"27",x"1e"),
   594 => (x"c4",x"0f",x"00",x"00"),
   595 => (x"12",x"36",x"27",x"86"),
   596 => (x"27",x"1e",x"00",x"00"),
   597 => (x"00",x"00",x"01",x"59"),
   598 => (x"27",x"86",x"c4",x"0f"),
   599 => (x"00",x"00",x"16",x"b8"),
   600 => (x"42",x"27",x"1e",x"bf"),
   601 => (x"1e",x"00",x"00",x"12"),
   602 => (x"00",x"01",x"59",x"27"),
   603 => (x"86",x"c8",x"0f",x"00"),
   604 => (x"00",x"12",x"5b",x"27"),
   605 => (x"59",x"27",x"1e",x"00"),
   606 => (x"0f",x"00",x"00",x"01"),
   607 => (x"b8",x"27",x"86",x"c4"),
   608 => (x"bf",x"00",x"00",x"16"),
   609 => (x"6a",x"82",x"c4",x"4a"),
   610 => (x"12",x"8c",x"27",x"1e"),
   611 => (x"27",x"1e",x"00",x"00"),
   612 => (x"00",x"00",x"01",x"59"),
   613 => (x"c0",x"86",x"c8",x"0f"),
   614 => (x"12",x"a5",x"27",x"1e"),
   615 => (x"27",x"1e",x"00",x"00"),
   616 => (x"00",x"00",x"01",x"59"),
   617 => (x"27",x"86",x"c8",x"0f"),
   618 => (x"00",x"00",x"16",x"b8"),
   619 => (x"82",x"c8",x"4a",x"bf"),
   620 => (x"be",x"27",x"1e",x"6a"),
   621 => (x"1e",x"00",x"00",x"12"),
   622 => (x"00",x"01",x"59",x"27"),
   623 => (x"86",x"c8",x"0f",x"00"),
   624 => (x"d7",x"27",x"1e",x"c2"),
   625 => (x"1e",x"00",x"00",x"12"),
   626 => (x"00",x"01",x"59",x"27"),
   627 => (x"86",x"c8",x"0f",x"00"),
   628 => (x"00",x"16",x"b8",x"27"),
   629 => (x"cc",x"4a",x"bf",x"00"),
   630 => (x"27",x"1e",x"6a",x"82"),
   631 => (x"00",x"00",x"12",x"f0"),
   632 => (x"01",x"59",x"27",x"1e"),
   633 => (x"c8",x"0f",x"00",x"00"),
   634 => (x"27",x"1e",x"d1",x"86"),
   635 => (x"00",x"00",x"13",x"09"),
   636 => (x"01",x"59",x"27",x"1e"),
   637 => (x"c8",x"0f",x"00",x"00"),
   638 => (x"16",x"b8",x"27",x"86"),
   639 => (x"4a",x"bf",x"00",x"00"),
   640 => (x"1e",x"72",x"82",x"d0"),
   641 => (x"00",x"13",x"22",x"27"),
   642 => (x"59",x"27",x"1e",x"00"),
   643 => (x"0f",x"00",x"00",x"01"),
   644 => (x"3b",x"27",x"86",x"c8"),
   645 => (x"1e",x"00",x"00",x"13"),
   646 => (x"00",x"01",x"59",x"27"),
   647 => (x"86",x"c4",x"0f",x"00"),
   648 => (x"00",x"13",x"70",x"27"),
   649 => (x"59",x"27",x"1e",x"00"),
   650 => (x"0f",x"00",x"00",x"01"),
   651 => (x"38",x"27",x"86",x"c4"),
   652 => (x"bf",x"00",x"00",x"17"),
   653 => (x"13",x"81",x"27",x"1e"),
   654 => (x"27",x"1e",x"00",x"00"),
   655 => (x"00",x"00",x"01",x"59"),
   656 => (x"27",x"86",x"c8",x"0f"),
   657 => (x"00",x"00",x"13",x"9a"),
   658 => (x"01",x"59",x"27",x"1e"),
   659 => (x"c4",x"0f",x"00",x"00"),
   660 => (x"17",x"38",x"27",x"86"),
   661 => (x"4a",x"bf",x"00",x"00"),
   662 => (x"1e",x"6a",x"82",x"c4"),
   663 => (x"00",x"13",x"da",x"27"),
   664 => (x"59",x"27",x"1e",x"00"),
   665 => (x"0f",x"00",x"00",x"01"),
   666 => (x"1e",x"c0",x"86",x"c8"),
   667 => (x"00",x"13",x"f3",x"27"),
   668 => (x"59",x"27",x"1e",x"00"),
   669 => (x"0f",x"00",x"00",x"01"),
   670 => (x"38",x"27",x"86",x"c8"),
   671 => (x"bf",x"00",x"00",x"17"),
   672 => (x"6a",x"82",x"c8",x"4a"),
   673 => (x"14",x"0c",x"27",x"1e"),
   674 => (x"27",x"1e",x"00",x"00"),
   675 => (x"00",x"00",x"01",x"59"),
   676 => (x"c1",x"86",x"c8",x"0f"),
   677 => (x"14",x"25",x"27",x"1e"),
   678 => (x"27",x"1e",x"00",x"00"),
   679 => (x"00",x"00",x"01",x"59"),
   680 => (x"27",x"86",x"c8",x"0f"),
   681 => (x"00",x"00",x"17",x"38"),
   682 => (x"82",x"cc",x"4a",x"bf"),
   683 => (x"3e",x"27",x"1e",x"6a"),
   684 => (x"1e",x"00",x"00",x"14"),
   685 => (x"00",x"01",x"59",x"27"),
   686 => (x"86",x"c8",x"0f",x"00"),
   687 => (x"57",x"27",x"1e",x"d2"),
   688 => (x"1e",x"00",x"00",x"14"),
   689 => (x"00",x"01",x"59",x"27"),
   690 => (x"86",x"c8",x"0f",x"00"),
   691 => (x"00",x"17",x"38",x"27"),
   692 => (x"d0",x"4a",x"bf",x"00"),
   693 => (x"27",x"1e",x"72",x"82"),
   694 => (x"00",x"00",x"14",x"70"),
   695 => (x"01",x"59",x"27",x"1e"),
   696 => (x"c8",x"0f",x"00",x"00"),
   697 => (x"14",x"89",x"27",x"86"),
   698 => (x"27",x"1e",x"00",x"00"),
   699 => (x"00",x"00",x"01",x"59"),
   700 => (x"6e",x"86",x"c4",x"0f"),
   701 => (x"14",x"be",x"27",x"1e"),
   702 => (x"27",x"1e",x"00",x"00"),
   703 => (x"00",x"00",x"01",x"59"),
   704 => (x"c5",x"86",x"c8",x"0f"),
   705 => (x"14",x"d7",x"27",x"1e"),
   706 => (x"27",x"1e",x"00",x"00"),
   707 => (x"00",x"00",x"01",x"59"),
   708 => (x"74",x"86",x"c8",x"0f"),
   709 => (x"14",x"f0",x"27",x"1e"),
   710 => (x"27",x"1e",x"00",x"00"),
   711 => (x"00",x"00",x"01",x"59"),
   712 => (x"cd",x"86",x"c8",x"0f"),
   713 => (x"15",x"09",x"27",x"1e"),
   714 => (x"27",x"1e",x"00",x"00"),
   715 => (x"00",x"00",x"01",x"59"),
   716 => (x"cc",x"86",x"c8",x"0f"),
   717 => (x"22",x"27",x"1e",x"66"),
   718 => (x"1e",x"00",x"00",x"15"),
   719 => (x"00",x"01",x"59",x"27"),
   720 => (x"86",x"c8",x"0f",x"00"),
   721 => (x"3b",x"27",x"1e",x"c7"),
   722 => (x"1e",x"00",x"00",x"15"),
   723 => (x"00",x"01",x"59",x"27"),
   724 => (x"86",x"c8",x"0f",x"00"),
   725 => (x"27",x"1e",x"66",x"c8"),
   726 => (x"00",x"00",x"15",x"54"),
   727 => (x"01",x"59",x"27",x"1e"),
   728 => (x"c8",x"0f",x"00",x"00"),
   729 => (x"27",x"1e",x"c1",x"86"),
   730 => (x"00",x"00",x"15",x"6d"),
   731 => (x"01",x"59",x"27",x"1e"),
   732 => (x"c8",x"0f",x"00",x"00"),
   733 => (x"16",x"c0",x"27",x"86"),
   734 => (x"27",x"1e",x"00",x"00"),
   735 => (x"00",x"00",x"15",x"86"),
   736 => (x"01",x"59",x"27",x"1e"),
   737 => (x"c8",x"0f",x"00",x"00"),
   738 => (x"15",x"9f",x"27",x"86"),
   739 => (x"27",x"1e",x"00",x"00"),
   740 => (x"00",x"00",x"01",x"59"),
   741 => (x"27",x"86",x"c4",x"0f"),
   742 => (x"00",x"00",x"16",x"e0"),
   743 => (x"15",x"d4",x"27",x"1e"),
   744 => (x"27",x"1e",x"00",x"00"),
   745 => (x"00",x"00",x"01",x"59"),
   746 => (x"27",x"86",x"c8",x"0f"),
   747 => (x"00",x"00",x"15",x"ed"),
   748 => (x"01",x"59",x"27",x"1e"),
   749 => (x"c4",x"0f",x"00",x"00"),
   750 => (x"16",x"22",x"27",x"86"),
   751 => (x"27",x"1e",x"00",x"00"),
   752 => (x"00",x"00",x"01",x"59"),
   753 => (x"27",x"86",x"c4",x"0f"),
   754 => (x"00",x"00",x"17",x"34"),
   755 => (x"b4",x"27",x"4a",x"bf"),
   756 => (x"bf",x"00",x"00",x"16"),
   757 => (x"16",x"bc",x"27",x"8a"),
   758 => (x"72",x"49",x"00",x"00"),
   759 => (x"27",x"1e",x"72",x"79"),
   760 => (x"00",x"00",x"16",x"24"),
   761 => (x"01",x"59",x"27",x"1e"),
   762 => (x"c8",x"0f",x"00",x"00"),
   763 => (x"16",x"bc",x"27",x"86"),
   764 => (x"49",x"bf",x"00",x"00"),
   765 => (x"a9",x"b7",x"f8",x"c1"),
   766 => (x"87",x"ea",x"c0",x"03"),
   767 => (x"00",x"0f",x"16",x"27"),
   768 => (x"59",x"27",x"1e",x"00"),
   769 => (x"0f",x"00",x"00",x"01"),
   770 => (x"4c",x"27",x"86",x"c4"),
   771 => (x"1e",x"00",x"00",x"0f"),
   772 => (x"00",x"01",x"59",x"27"),
   773 => (x"86",x"c4",x"0f",x"00"),
   774 => (x"00",x"0f",x"6c",x"27"),
   775 => (x"59",x"27",x"1e",x"00"),
   776 => (x"0f",x"00",x"00",x"01"),
   777 => (x"bc",x"27",x"86",x"c4"),
   778 => (x"bf",x"00",x"00",x"16"),
   779 => (x"cf",x"4b",x"72",x"4a"),
   780 => (x"49",x"73",x"93",x"e8"),
   781 => (x"38",x"27",x"1e",x"72"),
   782 => (x"bf",x"00",x"00",x"16"),
   783 => (x"04",x"c4",x"27",x"4a"),
   784 => (x"26",x"0f",x"00",x"00"),
   785 => (x"27",x"48",x"70",x"4a"),
   786 => (x"00",x"00",x"17",x"3c"),
   787 => (x"16",x"38",x"27",x"58"),
   788 => (x"4b",x"bf",x"00",x"00"),
   789 => (x"e8",x"cf",x"4c",x"73"),
   790 => (x"72",x"49",x"74",x"94"),
   791 => (x"27",x"4a",x"72",x"1e"),
   792 => (x"00",x"00",x"04",x"c4"),
   793 => (x"70",x"4a",x"26",x"0f"),
   794 => (x"16",x"b0",x"27",x"48"),
   795 => (x"c8",x"58",x"00",x"00"),
   796 => (x"49",x"73",x"93",x"f9"),
   797 => (x"4a",x"72",x"1e",x"72"),
   798 => (x"00",x"04",x"c4",x"27"),
   799 => (x"4a",x"26",x"0f",x"00"),
   800 => (x"44",x"27",x"48",x"70"),
   801 => (x"58",x"00",x"00",x"18"),
   802 => (x"00",x"0f",x"6e",x"27"),
   803 => (x"59",x"27",x"1e",x"00"),
   804 => (x"0f",x"00",x"00",x"01"),
   805 => (x"3c",x"27",x"86",x"c4"),
   806 => (x"bf",x"00",x"00",x"17"),
   807 => (x"0f",x"9b",x"27",x"1e"),
   808 => (x"27",x"1e",x"00",x"00"),
   809 => (x"00",x"00",x"01",x"59"),
   810 => (x"27",x"86",x"c8",x"0f"),
   811 => (x"00",x"00",x"0f",x"a0"),
   812 => (x"01",x"59",x"27",x"1e"),
   813 => (x"c4",x"0f",x"00",x"00"),
   814 => (x"16",x"b0",x"27",x"86"),
   815 => (x"1e",x"bf",x"00",x"00"),
   816 => (x"00",x"0f",x"cd",x"27"),
   817 => (x"59",x"27",x"1e",x"00"),
   818 => (x"0f",x"00",x"00",x"01"),
   819 => (x"44",x"27",x"86",x"c8"),
   820 => (x"bf",x"00",x"00",x"18"),
   821 => (x"0f",x"d2",x"27",x"1e"),
   822 => (x"27",x"1e",x"00",x"00"),
   823 => (x"00",x"00",x"01",x"59"),
   824 => (x"27",x"86",x"c8",x"0f"),
   825 => (x"00",x"00",x"0f",x"f0"),
   826 => (x"01",x"59",x"27",x"1e"),
   827 => (x"c4",x"0f",x"00",x"00"),
   828 => (x"d0",x"48",x"c0",x"86"),
   829 => (x"26",x"4d",x"26",x"86"),
   830 => (x"26",x"4b",x"26",x"4c"),
   831 => (x"0e",x"4f",x"26",x"4a"),
   832 => (x"5c",x"5b",x"5a",x"5e"),
   833 => (x"a6",x"d4",x"0e",x"5d"),
   834 => (x"72",x"4a",x"bf",x"bf"),
   835 => (x"16",x"b8",x"27",x"4d"),
   836 => (x"48",x"bf",x"00",x"00"),
   837 => (x"f0",x"c0",x"1e",x"72"),
   838 => (x"52",x"10",x"49",x"a2"),
   839 => (x"f9",x"05",x"a9",x"72"),
   840 => (x"d4",x"4a",x"26",x"87"),
   841 => (x"84",x"cc",x"4c",x"66"),
   842 => (x"4b",x"72",x"7c",x"c5"),
   843 => (x"7b",x"6c",x"83",x"cc"),
   844 => (x"bf",x"bf",x"a6",x"d4"),
   845 => (x"27",x"1e",x"72",x"7a"),
   846 => (x"00",x"00",x"0d",x"df"),
   847 => (x"c4",x"86",x"c4",x"0f"),
   848 => (x"05",x"9a",x"6a",x"82"),
   849 => (x"75",x"87",x"f3",x"c0"),
   850 => (x"75",x"83",x"c8",x"4b"),
   851 => (x"c6",x"82",x"cc",x"4a"),
   852 => (x"d8",x"1e",x"73",x"7a"),
   853 => (x"83",x"c8",x"4b",x"66"),
   854 => (x"a5",x"27",x"1e",x"6b"),
   855 => (x"0f",x"00",x"00",x"02"),
   856 => (x"b8",x"27",x"86",x"c8"),
   857 => (x"bf",x"00",x"00",x"16"),
   858 => (x"ca",x"1e",x"72",x"7d"),
   859 => (x"27",x"1e",x"6a",x"1e"),
   860 => (x"00",x"00",x"03",x"24"),
   861 => (x"c0",x"86",x"cc",x"0f"),
   862 => (x"a6",x"d4",x"87",x"d9"),
   863 => (x"d4",x"4a",x"bf",x"bf"),
   864 => (x"48",x"49",x"bf",x"a6"),
   865 => (x"f0",x"c0",x"1e",x"72"),
   866 => (x"51",x"10",x"4a",x"a1"),
   867 => (x"f9",x"05",x"aa",x"71"),
   868 => (x"26",x"4a",x"26",x"87"),
   869 => (x"26",x"4c",x"26",x"4d"),
   870 => (x"26",x"4a",x"26",x"4b"),
   871 => (x"5a",x"5e",x"0e",x"4f"),
   872 => (x"d0",x"1e",x"0e",x"5b"),
   873 => (x"4b",x"bf",x"bf",x"a6"),
   874 => (x"30",x"27",x"83",x"ca"),
   875 => (x"97",x"00",x"00",x"17"),
   876 => (x"32",x"d8",x"4a",x"bf"),
   877 => (x"49",x"72",x"2a",x"b7"),
   878 => (x"a9",x"b7",x"c1",x"c1"),
   879 => (x"87",x"d3",x"c0",x"05"),
   880 => (x"48",x"73",x"8b",x"c1"),
   881 => (x"00",x"18",x"3c",x"27"),
   882 => (x"d0",x"88",x"bf",x"00"),
   883 => (x"76",x"58",x"49",x"66"),
   884 => (x"6e",x"79",x"c0",x"49"),
   885 => (x"87",x"d2",x"ff",x"05"),
   886 => (x"26",x"4b",x"26",x"26"),
   887 => (x"1e",x"4f",x"26",x"4a"),
   888 => (x"b8",x"27",x"1e",x"72"),
   889 => (x"bf",x"00",x"00",x"16"),
   890 => (x"87",x"cb",x"c0",x"02"),
   891 => (x"49",x"bf",x"a6",x"c8"),
   892 => (x"00",x"16",x"b8",x"27"),
   893 => (x"27",x"79",x"bf",x"00"),
   894 => (x"00",x"00",x"16",x"b8"),
   895 => (x"82",x"cc",x"4a",x"bf"),
   896 => (x"3c",x"27",x"1e",x"72"),
   897 => (x"bf",x"00",x"00",x"18"),
   898 => (x"27",x"1e",x"ca",x"1e"),
   899 => (x"00",x"00",x"03",x"24"),
   900 => (x"26",x"86",x"cc",x"0f"),
   901 => (x"1e",x"4f",x"26",x"4a"),
   902 => (x"30",x"27",x"1e",x"72"),
   903 => (x"97",x"00",x"00",x"17"),
   904 => (x"32",x"d8",x"4a",x"bf"),
   905 => (x"49",x"72",x"2a",x"b7"),
   906 => (x"a9",x"b7",x"c1",x"c1"),
   907 => (x"87",x"c5",x"c0",x"02"),
   908 => (x"c2",x"c0",x"4a",x"c0"),
   909 => (x"27",x"4a",x"c1",x"87"),
   910 => (x"00",x"00",x"18",x"40"),
   911 => (x"b0",x"72",x"48",x"bf"),
   912 => (x"00",x"18",x"40",x"27"),
   913 => (x"38",x"27",x"58",x"00"),
   914 => (x"49",x"00",x"00",x"18"),
   915 => (x"26",x"51",x"c2",x"c1"),
   916 => (x"1e",x"4f",x"26",x"4a"),
   917 => (x"00",x"17",x"30",x"27"),
   918 => (x"c1",x"c1",x"49",x"00"),
   919 => (x"18",x"40",x"27",x"51"),
   920 => (x"c0",x"49",x"00",x"00"),
   921 => (x"00",x"4f",x"26",x"79"),
   922 => (x"33",x"32",x"31",x"30"),
   923 => (x"37",x"36",x"35",x"34"),
   924 => (x"42",x"41",x"39",x"38"),
   925 => (x"46",x"45",x"44",x"43"),
   926 => (x"6f",x"72",x"50",x"00"),
   927 => (x"6d",x"61",x"72",x"67"),
   928 => (x"6d",x"6f",x"63",x"20"),
   929 => (x"65",x"6c",x"69",x"70"),
   930 => (x"69",x"77",x"20",x"64"),
   931 => (x"27",x"20",x"68",x"74"),
   932 => (x"69",x"67",x"65",x"72"),
   933 => (x"72",x"65",x"74",x"73"),
   934 => (x"74",x"61",x"20",x"27"),
   935 => (x"62",x"69",x"72",x"74"),
   936 => (x"0a",x"65",x"74",x"75"),
   937 => (x"50",x"00",x"0a",x"00"),
   938 => (x"72",x"67",x"6f",x"72"),
   939 => (x"63",x"20",x"6d",x"61"),
   940 => (x"69",x"70",x"6d",x"6f"),
   941 => (x"20",x"64",x"65",x"6c"),
   942 => (x"68",x"74",x"69",x"77"),
   943 => (x"20",x"74",x"75",x"6f"),
   944 => (x"67",x"65",x"72",x"27"),
   945 => (x"65",x"74",x"73",x"69"),
   946 => (x"61",x"20",x"27",x"72"),
   947 => (x"69",x"72",x"74",x"74"),
   948 => (x"65",x"74",x"75",x"62"),
   949 => (x"00",x"0a",x"00",x"0a"),
   950 => (x"59",x"52",x"48",x"44"),
   951 => (x"4e",x"4f",x"54",x"53"),
   952 => (x"52",x"50",x"20",x"45"),
   953 => (x"41",x"52",x"47",x"4f"),
   954 => (x"33",x"20",x"2c",x"4d"),
   955 => (x"20",x"44",x"52",x"27"),
   956 => (x"49",x"52",x"54",x"53"),
   957 => (x"44",x"00",x"47",x"4e"),
   958 => (x"53",x"59",x"52",x"48"),
   959 => (x"45",x"4e",x"4f",x"54"),
   960 => (x"4f",x"52",x"50",x"20"),
   961 => (x"4d",x"41",x"52",x"47"),
   962 => (x"27",x"32",x"20",x"2c"),
   963 => (x"53",x"20",x"44",x"4e"),
   964 => (x"4e",x"49",x"52",x"54"),
   965 => (x"65",x"4d",x"00",x"47"),
   966 => (x"72",x"75",x"73",x"61"),
   967 => (x"74",x"20",x"64",x"65"),
   968 => (x"20",x"65",x"6d",x"69"),
   969 => (x"20",x"6f",x"6f",x"74"),
   970 => (x"6c",x"61",x"6d",x"73"),
   971 => (x"6f",x"74",x"20",x"6c"),
   972 => (x"74",x"62",x"6f",x"20"),
   973 => (x"20",x"6e",x"69",x"61"),
   974 => (x"6e",x"61",x"65",x"6d"),
   975 => (x"66",x"67",x"6e",x"69"),
   976 => (x"72",x"20",x"6c",x"75"),
   977 => (x"6c",x"75",x"73",x"65"),
   978 => (x"00",x"0a",x"73",x"74"),
   979 => (x"61",x"65",x"6c",x"50"),
   980 => (x"69",x"20",x"65",x"73"),
   981 => (x"65",x"72",x"63",x"6e"),
   982 => (x"20",x"65",x"73",x"61"),
   983 => (x"62",x"6d",x"75",x"6e"),
   984 => (x"6f",x"20",x"72",x"65"),
   985 => (x"75",x"72",x"20",x"66"),
   986 => (x"00",x"0a",x"73",x"6e"),
   987 => (x"69",x"4d",x"00",x"0a"),
   988 => (x"73",x"6f",x"72",x"63"),
   989 => (x"6e",x"6f",x"63",x"65"),
   990 => (x"66",x"20",x"73",x"64"),
   991 => (x"6f",x"20",x"72",x"6f"),
   992 => (x"72",x"20",x"65",x"6e"),
   993 => (x"74",x"20",x"6e",x"75"),
   994 => (x"75",x"6f",x"72",x"68"),
   995 => (x"44",x"20",x"68",x"67"),
   996 => (x"73",x"79",x"72",x"68"),
   997 => (x"65",x"6e",x"6f",x"74"),
   998 => (x"25",x"00",x"20",x"3a"),
   999 => (x"00",x"0a",x"20",x"64"),
  1000 => (x"79",x"72",x"68",x"44"),
  1001 => (x"6e",x"6f",x"74",x"73"),
  1002 => (x"70",x"20",x"73",x"65"),
  1003 => (x"53",x"20",x"72",x"65"),
  1004 => (x"6e",x"6f",x"63",x"65"),
  1005 => (x"20",x"20",x"3a",x"64"),
  1006 => (x"20",x"20",x"20",x"20"),
  1007 => (x"20",x"20",x"20",x"20"),
  1008 => (x"20",x"20",x"20",x"20"),
  1009 => (x"20",x"20",x"20",x"20"),
  1010 => (x"20",x"20",x"20",x"20"),
  1011 => (x"20",x"64",x"25",x"00"),
  1012 => (x"41",x"56",x"00",x"0a"),
  1013 => (x"49",x"4d",x"20",x"58"),
  1014 => (x"72",x"20",x"53",x"50"),
  1015 => (x"6e",x"69",x"74",x"61"),
  1016 => (x"20",x"2a",x"20",x"67"),
  1017 => (x"30",x"30",x"30",x"31"),
  1018 => (x"25",x"20",x"3d",x"20"),
  1019 => (x"00",x"0a",x"20",x"64"),
  1020 => (x"48",x"44",x"00",x"0a"),
  1021 => (x"54",x"53",x"59",x"52"),
  1022 => (x"20",x"45",x"4e",x"4f"),
  1023 => (x"47",x"4f",x"52",x"50"),
  1024 => (x"2c",x"4d",x"41",x"52"),
  1025 => (x"4d",x"4f",x"53",x"20"),
  1026 => (x"54",x"53",x"20",x"45"),
  1027 => (x"47",x"4e",x"49",x"52"),
  1028 => (x"52",x"48",x"44",x"00"),
  1029 => (x"4f",x"54",x"53",x"59"),
  1030 => (x"50",x"20",x"45",x"4e"),
  1031 => (x"52",x"47",x"4f",x"52"),
  1032 => (x"20",x"2c",x"4d",x"41"),
  1033 => (x"54",x"53",x"27",x"31"),
  1034 => (x"52",x"54",x"53",x"20"),
  1035 => (x"00",x"47",x"4e",x"49"),
  1036 => (x"68",x"44",x"00",x"0a"),
  1037 => (x"74",x"73",x"79",x"72"),
  1038 => (x"20",x"65",x"6e",x"6f"),
  1039 => (x"63",x"6e",x"65",x"42"),
  1040 => (x"72",x"61",x"6d",x"68"),
  1041 => (x"56",x"20",x"2c",x"6b"),
  1042 => (x"69",x"73",x"72",x"65"),
  1043 => (x"32",x"20",x"6e",x"6f"),
  1044 => (x"28",x"20",x"31",x"2e"),
  1045 => (x"67",x"6e",x"61",x"4c"),
  1046 => (x"65",x"67",x"61",x"75"),
  1047 => (x"29",x"43",x"20",x"3a"),
  1048 => (x"00",x"0a",x"00",x"0a"),
  1049 => (x"63",x"65",x"78",x"45"),
  1050 => (x"6f",x"69",x"74",x"75"),
  1051 => (x"74",x"73",x"20",x"6e"),
  1052 => (x"73",x"74",x"72",x"61"),
  1053 => (x"64",x"25",x"20",x"2c"),
  1054 => (x"6e",x"75",x"72",x"20"),
  1055 => (x"68",x"74",x"20",x"73"),
  1056 => (x"67",x"75",x"6f",x"72"),
  1057 => (x"68",x"44",x"20",x"68"),
  1058 => (x"74",x"73",x"79",x"72"),
  1059 => (x"0a",x"65",x"6e",x"6f"),
  1060 => (x"67",x"65",x"42",x"00"),
  1061 => (x"74",x"20",x"6e",x"69"),
  1062 => (x"3a",x"65",x"6d",x"69"),
  1063 => (x"0a",x"64",x"25",x"20"),
  1064 => (x"64",x"6e",x"45",x"00"),
  1065 => (x"6d",x"69",x"74",x"20"),
  1066 => (x"25",x"20",x"3a",x"65"),
  1067 => (x"45",x"00",x"0a",x"64"),
  1068 => (x"75",x"63",x"65",x"78"),
  1069 => (x"6e",x"6f",x"69",x"74"),
  1070 => (x"64",x"6e",x"65",x"20"),
  1071 => (x"0a",x"00",x"0a",x"73"),
  1072 => (x"6e",x"69",x"46",x"00"),
  1073 => (x"76",x"20",x"6c",x"61"),
  1074 => (x"65",x"75",x"6c",x"61"),
  1075 => (x"66",x"6f",x"20",x"73"),
  1076 => (x"65",x"68",x"74",x"20"),
  1077 => (x"72",x"61",x"76",x"20"),
  1078 => (x"6c",x"62",x"61",x"69"),
  1079 => (x"75",x"20",x"73",x"65"),
  1080 => (x"20",x"64",x"65",x"73"),
  1081 => (x"74",x"20",x"6e",x"69"),
  1082 => (x"62",x"20",x"65",x"68"),
  1083 => (x"68",x"63",x"6e",x"65"),
  1084 => (x"6b",x"72",x"61",x"6d"),
  1085 => (x"0a",x"00",x"0a",x"3a"),
  1086 => (x"74",x"6e",x"49",x"00"),
  1087 => (x"6f",x"6c",x"47",x"5f"),
  1088 => (x"20",x"20",x"3a",x"62"),
  1089 => (x"20",x"20",x"20",x"20"),
  1090 => (x"20",x"20",x"20",x"20"),
  1091 => (x"64",x"25",x"20",x"20"),
  1092 => (x"20",x"20",x"00",x"0a"),
  1093 => (x"20",x"20",x"20",x"20"),
  1094 => (x"68",x"73",x"20",x"20"),
  1095 => (x"64",x"6c",x"75",x"6f"),
  1096 => (x"3a",x"65",x"62",x"20"),
  1097 => (x"25",x"20",x"20",x"20"),
  1098 => (x"42",x"00",x"0a",x"64"),
  1099 => (x"5f",x"6c",x"6f",x"6f"),
  1100 => (x"62",x"6f",x"6c",x"47"),
  1101 => (x"20",x"20",x"20",x"3a"),
  1102 => (x"20",x"20",x"20",x"20"),
  1103 => (x"20",x"20",x"20",x"20"),
  1104 => (x"00",x"0a",x"64",x"25"),
  1105 => (x"20",x"20",x"20",x"20"),
  1106 => (x"20",x"20",x"20",x"20"),
  1107 => (x"75",x"6f",x"68",x"73"),
  1108 => (x"62",x"20",x"64",x"6c"),
  1109 => (x"20",x"20",x"3a",x"65"),
  1110 => (x"0a",x"64",x"25",x"20"),
  1111 => (x"5f",x"68",x"43",x"00"),
  1112 => (x"6c",x"47",x"5f",x"31"),
  1113 => (x"20",x"3a",x"62",x"6f"),
  1114 => (x"20",x"20",x"20",x"20"),
  1115 => (x"20",x"20",x"20",x"20"),
  1116 => (x"63",x"25",x"20",x"20"),
  1117 => (x"20",x"20",x"00",x"0a"),
  1118 => (x"20",x"20",x"20",x"20"),
  1119 => (x"68",x"73",x"20",x"20"),
  1120 => (x"64",x"6c",x"75",x"6f"),
  1121 => (x"3a",x"65",x"62",x"20"),
  1122 => (x"25",x"20",x"20",x"20"),
  1123 => (x"43",x"00",x"0a",x"63"),
  1124 => (x"5f",x"32",x"5f",x"68"),
  1125 => (x"62",x"6f",x"6c",x"47"),
  1126 => (x"20",x"20",x"20",x"3a"),
  1127 => (x"20",x"20",x"20",x"20"),
  1128 => (x"20",x"20",x"20",x"20"),
  1129 => (x"00",x"0a",x"63",x"25"),
  1130 => (x"20",x"20",x"20",x"20"),
  1131 => (x"20",x"20",x"20",x"20"),
  1132 => (x"75",x"6f",x"68",x"73"),
  1133 => (x"62",x"20",x"64",x"6c"),
  1134 => (x"20",x"20",x"3a",x"65"),
  1135 => (x"0a",x"63",x"25",x"20"),
  1136 => (x"72",x"72",x"41",x"00"),
  1137 => (x"47",x"5f",x"31",x"5f"),
  1138 => (x"5b",x"62",x"6f",x"6c"),
  1139 => (x"20",x"3a",x"5d",x"38"),
  1140 => (x"20",x"20",x"20",x"20"),
  1141 => (x"64",x"25",x"20",x"20"),
  1142 => (x"20",x"20",x"00",x"0a"),
  1143 => (x"20",x"20",x"20",x"20"),
  1144 => (x"68",x"73",x"20",x"20"),
  1145 => (x"64",x"6c",x"75",x"6f"),
  1146 => (x"3a",x"65",x"62",x"20"),
  1147 => (x"25",x"20",x"20",x"20"),
  1148 => (x"41",x"00",x"0a",x"64"),
  1149 => (x"32",x"5f",x"72",x"72"),
  1150 => (x"6f",x"6c",x"47",x"5f"),
  1151 => (x"5d",x"38",x"5b",x"62"),
  1152 => (x"3a",x"5d",x"37",x"5b"),
  1153 => (x"20",x"20",x"20",x"20"),
  1154 => (x"00",x"0a",x"64",x"25"),
  1155 => (x"20",x"20",x"20",x"20"),
  1156 => (x"20",x"20",x"20",x"20"),
  1157 => (x"75",x"6f",x"68",x"73"),
  1158 => (x"62",x"20",x"64",x"6c"),
  1159 => (x"20",x"20",x"3a",x"65"),
  1160 => (x"6d",x"75",x"4e",x"20"),
  1161 => (x"5f",x"72",x"65",x"62"),
  1162 => (x"52",x"5f",x"66",x"4f"),
  1163 => (x"20",x"73",x"6e",x"75"),
  1164 => (x"30",x"31",x"20",x"2b"),
  1165 => (x"74",x"50",x"00",x"0a"),
  1166 => (x"6c",x"47",x"5f",x"72"),
  1167 => (x"3e",x"2d",x"62",x"6f"),
  1168 => (x"20",x"20",x"00",x"0a"),
  1169 => (x"5f",x"72",x"74",x"50"),
  1170 => (x"70",x"6d",x"6f",x"43"),
  1171 => (x"20",x"20",x"20",x"3a"),
  1172 => (x"20",x"20",x"20",x"20"),
  1173 => (x"25",x"20",x"20",x"20"),
  1174 => (x"20",x"00",x"0a",x"64"),
  1175 => (x"20",x"20",x"20",x"20"),
  1176 => (x"73",x"20",x"20",x"20"),
  1177 => (x"6c",x"75",x"6f",x"68"),
  1178 => (x"65",x"62",x"20",x"64"),
  1179 => (x"20",x"20",x"20",x"3a"),
  1180 => (x"70",x"6d",x"69",x"28"),
  1181 => (x"65",x"6d",x"65",x"6c"),
  1182 => (x"74",x"61",x"74",x"6e"),
  1183 => (x"2d",x"6e",x"6f",x"69"),
  1184 => (x"65",x"70",x"65",x"64"),
  1185 => (x"6e",x"65",x"64",x"6e"),
  1186 => (x"00",x"0a",x"29",x"74"),
  1187 => (x"69",x"44",x"20",x"20"),
  1188 => (x"3a",x"72",x"63",x"73"),
  1189 => (x"20",x"20",x"20",x"20"),
  1190 => (x"20",x"20",x"20",x"20"),
  1191 => (x"20",x"20",x"20",x"20"),
  1192 => (x"0a",x"64",x"25",x"20"),
  1193 => (x"20",x"20",x"20",x"00"),
  1194 => (x"20",x"20",x"20",x"20"),
  1195 => (x"6f",x"68",x"73",x"20"),
  1196 => (x"20",x"64",x"6c",x"75"),
  1197 => (x"20",x"3a",x"65",x"62"),
  1198 => (x"64",x"25",x"20",x"20"),
  1199 => (x"20",x"20",x"00",x"0a"),
  1200 => (x"6d",x"75",x"6e",x"45"),
  1201 => (x"6d",x"6f",x"43",x"5f"),
  1202 => (x"20",x"20",x"3a",x"70"),
  1203 => (x"20",x"20",x"20",x"20"),
  1204 => (x"25",x"20",x"20",x"20"),
  1205 => (x"20",x"00",x"0a",x"64"),
  1206 => (x"20",x"20",x"20",x"20"),
  1207 => (x"73",x"20",x"20",x"20"),
  1208 => (x"6c",x"75",x"6f",x"68"),
  1209 => (x"65",x"62",x"20",x"64"),
  1210 => (x"20",x"20",x"20",x"3a"),
  1211 => (x"00",x"0a",x"64",x"25"),
  1212 => (x"6e",x"49",x"20",x"20"),
  1213 => (x"6f",x"43",x"5f",x"74"),
  1214 => (x"20",x"3a",x"70",x"6d"),
  1215 => (x"20",x"20",x"20",x"20"),
  1216 => (x"20",x"20",x"20",x"20"),
  1217 => (x"0a",x"64",x"25",x"20"),
  1218 => (x"20",x"20",x"20",x"00"),
  1219 => (x"20",x"20",x"20",x"20"),
  1220 => (x"6f",x"68",x"73",x"20"),
  1221 => (x"20",x"64",x"6c",x"75"),
  1222 => (x"20",x"3a",x"65",x"62"),
  1223 => (x"64",x"25",x"20",x"20"),
  1224 => (x"20",x"20",x"00",x"0a"),
  1225 => (x"5f",x"72",x"74",x"53"),
  1226 => (x"70",x"6d",x"6f",x"43"),
  1227 => (x"20",x"20",x"20",x"3a"),
  1228 => (x"20",x"20",x"20",x"20"),
  1229 => (x"25",x"20",x"20",x"20"),
  1230 => (x"20",x"00",x"0a",x"73"),
  1231 => (x"20",x"20",x"20",x"20"),
  1232 => (x"73",x"20",x"20",x"20"),
  1233 => (x"6c",x"75",x"6f",x"68"),
  1234 => (x"65",x"62",x"20",x"64"),
  1235 => (x"20",x"20",x"20",x"3a"),
  1236 => (x"59",x"52",x"48",x"44"),
  1237 => (x"4e",x"4f",x"54",x"53"),
  1238 => (x"52",x"50",x"20",x"45"),
  1239 => (x"41",x"52",x"47",x"4f"),
  1240 => (x"53",x"20",x"2c",x"4d"),
  1241 => (x"20",x"45",x"4d",x"4f"),
  1242 => (x"49",x"52",x"54",x"53"),
  1243 => (x"00",x"0a",x"47",x"4e"),
  1244 => (x"74",x"78",x"65",x"4e"),
  1245 => (x"72",x"74",x"50",x"5f"),
  1246 => (x"6f",x"6c",x"47",x"5f"),
  1247 => (x"0a",x"3e",x"2d",x"62"),
  1248 => (x"50",x"20",x"20",x"00"),
  1249 => (x"43",x"5f",x"72",x"74"),
  1250 => (x"3a",x"70",x"6d",x"6f"),
  1251 => (x"20",x"20",x"20",x"20"),
  1252 => (x"20",x"20",x"20",x"20"),
  1253 => (x"64",x"25",x"20",x"20"),
  1254 => (x"20",x"20",x"00",x"0a"),
  1255 => (x"20",x"20",x"20",x"20"),
  1256 => (x"68",x"73",x"20",x"20"),
  1257 => (x"64",x"6c",x"75",x"6f"),
  1258 => (x"3a",x"65",x"62",x"20"),
  1259 => (x"28",x"20",x"20",x"20"),
  1260 => (x"6c",x"70",x"6d",x"69"),
  1261 => (x"6e",x"65",x"6d",x"65"),
  1262 => (x"69",x"74",x"61",x"74"),
  1263 => (x"64",x"2d",x"6e",x"6f"),
  1264 => (x"6e",x"65",x"70",x"65"),
  1265 => (x"74",x"6e",x"65",x"64"),
  1266 => (x"73",x"20",x"2c",x"29"),
  1267 => (x"20",x"65",x"6d",x"61"),
  1268 => (x"61",x"20",x"73",x"61"),
  1269 => (x"65",x"76",x"6f",x"62"),
  1270 => (x"20",x"20",x"00",x"0a"),
  1271 => (x"63",x"73",x"69",x"44"),
  1272 => (x"20",x"20",x"3a",x"72"),
  1273 => (x"20",x"20",x"20",x"20"),
  1274 => (x"20",x"20",x"20",x"20"),
  1275 => (x"25",x"20",x"20",x"20"),
  1276 => (x"20",x"00",x"0a",x"64"),
  1277 => (x"20",x"20",x"20",x"20"),
  1278 => (x"73",x"20",x"20",x"20"),
  1279 => (x"6c",x"75",x"6f",x"68"),
  1280 => (x"65",x"62",x"20",x"64"),
  1281 => (x"20",x"20",x"20",x"3a"),
  1282 => (x"00",x"0a",x"64",x"25"),
  1283 => (x"6e",x"45",x"20",x"20"),
  1284 => (x"43",x"5f",x"6d",x"75"),
  1285 => (x"3a",x"70",x"6d",x"6f"),
  1286 => (x"20",x"20",x"20",x"20"),
  1287 => (x"20",x"20",x"20",x"20"),
  1288 => (x"0a",x"64",x"25",x"20"),
  1289 => (x"20",x"20",x"20",x"00"),
  1290 => (x"20",x"20",x"20",x"20"),
  1291 => (x"6f",x"68",x"73",x"20"),
  1292 => (x"20",x"64",x"6c",x"75"),
  1293 => (x"20",x"3a",x"65",x"62"),
  1294 => (x"64",x"25",x"20",x"20"),
  1295 => (x"20",x"20",x"00",x"0a"),
  1296 => (x"5f",x"74",x"6e",x"49"),
  1297 => (x"70",x"6d",x"6f",x"43"),
  1298 => (x"20",x"20",x"20",x"3a"),
  1299 => (x"20",x"20",x"20",x"20"),
  1300 => (x"25",x"20",x"20",x"20"),
  1301 => (x"20",x"00",x"0a",x"64"),
  1302 => (x"20",x"20",x"20",x"20"),
  1303 => (x"73",x"20",x"20",x"20"),
  1304 => (x"6c",x"75",x"6f",x"68"),
  1305 => (x"65",x"62",x"20",x"64"),
  1306 => (x"20",x"20",x"20",x"3a"),
  1307 => (x"00",x"0a",x"64",x"25"),
  1308 => (x"74",x"53",x"20",x"20"),
  1309 => (x"6f",x"43",x"5f",x"72"),
  1310 => (x"20",x"3a",x"70",x"6d"),
  1311 => (x"20",x"20",x"20",x"20"),
  1312 => (x"20",x"20",x"20",x"20"),
  1313 => (x"0a",x"73",x"25",x"20"),
  1314 => (x"20",x"20",x"20",x"00"),
  1315 => (x"20",x"20",x"20",x"20"),
  1316 => (x"6f",x"68",x"73",x"20"),
  1317 => (x"20",x"64",x"6c",x"75"),
  1318 => (x"20",x"3a",x"65",x"62"),
  1319 => (x"48",x"44",x"20",x"20"),
  1320 => (x"54",x"53",x"59",x"52"),
  1321 => (x"20",x"45",x"4e",x"4f"),
  1322 => (x"47",x"4f",x"52",x"50"),
  1323 => (x"2c",x"4d",x"41",x"52"),
  1324 => (x"4d",x"4f",x"53",x"20"),
  1325 => (x"54",x"53",x"20",x"45"),
  1326 => (x"47",x"4e",x"49",x"52"),
  1327 => (x"6e",x"49",x"00",x"0a"),
  1328 => (x"5f",x"31",x"5f",x"74"),
  1329 => (x"3a",x"63",x"6f",x"4c"),
  1330 => (x"20",x"20",x"20",x"20"),
  1331 => (x"20",x"20",x"20",x"20"),
  1332 => (x"25",x"20",x"20",x"20"),
  1333 => (x"20",x"00",x"0a",x"64"),
  1334 => (x"20",x"20",x"20",x"20"),
  1335 => (x"73",x"20",x"20",x"20"),
  1336 => (x"6c",x"75",x"6f",x"68"),
  1337 => (x"65",x"62",x"20",x"64"),
  1338 => (x"20",x"20",x"20",x"3a"),
  1339 => (x"00",x"0a",x"64",x"25"),
  1340 => (x"5f",x"74",x"6e",x"49"),
  1341 => (x"6f",x"4c",x"5f",x"32"),
  1342 => (x"20",x"20",x"3a",x"63"),
  1343 => (x"20",x"20",x"20",x"20"),
  1344 => (x"20",x"20",x"20",x"20"),
  1345 => (x"0a",x"64",x"25",x"20"),
  1346 => (x"20",x"20",x"20",x"00"),
  1347 => (x"20",x"20",x"20",x"20"),
  1348 => (x"6f",x"68",x"73",x"20"),
  1349 => (x"20",x"64",x"6c",x"75"),
  1350 => (x"20",x"3a",x"65",x"62"),
  1351 => (x"64",x"25",x"20",x"20"),
  1352 => (x"6e",x"49",x"00",x"0a"),
  1353 => (x"5f",x"33",x"5f",x"74"),
  1354 => (x"3a",x"63",x"6f",x"4c"),
  1355 => (x"20",x"20",x"20",x"20"),
  1356 => (x"20",x"20",x"20",x"20"),
  1357 => (x"25",x"20",x"20",x"20"),
  1358 => (x"20",x"00",x"0a",x"64"),
  1359 => (x"20",x"20",x"20",x"20"),
  1360 => (x"73",x"20",x"20",x"20"),
  1361 => (x"6c",x"75",x"6f",x"68"),
  1362 => (x"65",x"62",x"20",x"64"),
  1363 => (x"20",x"20",x"20",x"3a"),
  1364 => (x"00",x"0a",x"64",x"25"),
  1365 => (x"6d",x"75",x"6e",x"45"),
  1366 => (x"63",x"6f",x"4c",x"5f"),
  1367 => (x"20",x"20",x"20",x"3a"),
  1368 => (x"20",x"20",x"20",x"20"),
  1369 => (x"20",x"20",x"20",x"20"),
  1370 => (x"0a",x"64",x"25",x"20"),
  1371 => (x"20",x"20",x"20",x"00"),
  1372 => (x"20",x"20",x"20",x"20"),
  1373 => (x"6f",x"68",x"73",x"20"),
  1374 => (x"20",x"64",x"6c",x"75"),
  1375 => (x"20",x"3a",x"65",x"62"),
  1376 => (x"64",x"25",x"20",x"20"),
  1377 => (x"74",x"53",x"00",x"0a"),
  1378 => (x"5f",x"31",x"5f",x"72"),
  1379 => (x"3a",x"63",x"6f",x"4c"),
  1380 => (x"20",x"20",x"20",x"20"),
  1381 => (x"20",x"20",x"20",x"20"),
  1382 => (x"25",x"20",x"20",x"20"),
  1383 => (x"20",x"00",x"0a",x"73"),
  1384 => (x"20",x"20",x"20",x"20"),
  1385 => (x"73",x"20",x"20",x"20"),
  1386 => (x"6c",x"75",x"6f",x"68"),
  1387 => (x"65",x"62",x"20",x"64"),
  1388 => (x"20",x"20",x"20",x"3a"),
  1389 => (x"59",x"52",x"48",x"44"),
  1390 => (x"4e",x"4f",x"54",x"53"),
  1391 => (x"52",x"50",x"20",x"45"),
  1392 => (x"41",x"52",x"47",x"4f"),
  1393 => (x"31",x"20",x"2c",x"4d"),
  1394 => (x"20",x"54",x"53",x"27"),
  1395 => (x"49",x"52",x"54",x"53"),
  1396 => (x"00",x"0a",x"47",x"4e"),
  1397 => (x"5f",x"72",x"74",x"53"),
  1398 => (x"6f",x"4c",x"5f",x"32"),
  1399 => (x"20",x"20",x"3a",x"63"),
  1400 => (x"20",x"20",x"20",x"20"),
  1401 => (x"20",x"20",x"20",x"20"),
  1402 => (x"0a",x"73",x"25",x"20"),
  1403 => (x"20",x"20",x"20",x"00"),
  1404 => (x"20",x"20",x"20",x"20"),
  1405 => (x"6f",x"68",x"73",x"20"),
  1406 => (x"20",x"64",x"6c",x"75"),
  1407 => (x"20",x"3a",x"65",x"62"),
  1408 => (x"48",x"44",x"20",x"20"),
  1409 => (x"54",x"53",x"59",x"52"),
  1410 => (x"20",x"45",x"4e",x"4f"),
  1411 => (x"47",x"4f",x"52",x"50"),
  1412 => (x"2c",x"4d",x"41",x"52"),
  1413 => (x"4e",x"27",x"32",x"20"),
  1414 => (x"54",x"53",x"20",x"44"),
  1415 => (x"47",x"4e",x"49",x"52"),
  1416 => (x"00",x"0a",x"00",x"0a"),
  1417 => (x"72",x"65",x"73",x"55"),
  1418 => (x"6d",x"69",x"74",x"20"),
  1419 => (x"25",x"20",x"3a",x"65"),
  1420 => (x"00",x"00",x"0a",x"64"),
  1421 => (x"00",x"00",x"00",x"00"),
  1422 => (x"00",x"00",x"61",x"a8"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
