
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"3b",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"38"),
    10 => (x"80",x"00",x"27",x"4f"),
    11 => (x"27",x"4e",x"00",x"00"),
    12 => (x"00",x"00",x"04",x"04"),
    13 => (x"87",x"fd",x"00",x"0f"),
    14 => (x"4f",x"87",x"fd",x"00"),
    15 => (x"ff",x"86",x"fc",x"1e"),
    16 => (x"48",x"69",x"49",x"c0"),
    17 => (x"c4",x"98",x"c0",x"c4"),
    18 => (x"02",x"6e",x"58",x"a6"),
    19 => (x"66",x"c8",x"87",x"f4"),
    20 => (x"8e",x"fc",x"48",x"79"),
    21 => (x"5e",x"0e",x"4f",x"26"),
    22 => (x"0e",x"5d",x"5c",x"5b"),
    23 => (x"c0",x"4b",x"66",x"d0"),
    24 => (x"c3",x"49",x"13",x"4c"),
    25 => (x"99",x"71",x"99",x"ff"),
    26 => (x"71",x"87",x"dd",x"02"),
    27 => (x"4a",x"c0",x"ff",x"4d"),
    28 => (x"c0",x"c4",x"49",x"6a"),
    29 => (x"02",x"99",x"71",x"99"),
    30 => (x"7a",x"75",x"87",x"f6"),
    31 => (x"49",x"13",x"84",x"c1"),
    32 => (x"71",x"99",x"ff",x"c3"),
    33 => (x"87",x"e3",x"05",x"99"),
    34 => (x"4d",x"26",x"48",x"74"),
    35 => (x"4b",x"26",x"4c",x"26"),
    36 => (x"5e",x"0e",x"4f",x"26"),
    37 => (x"0e",x"5d",x"5c",x"5b"),
    38 => (x"f4",x"c0",x"86",x"e4"),
    39 => (x"a6",x"c4",x"4d",x"66"),
    40 => (x"c4",x"78",x"c0",x"48"),
    41 => (x"c0",x"78",x"c0",x"80"),
    42 => (x"bf",x"97",x"66",x"ec"),
    43 => (x"83",x"c0",x"fe",x"4b"),
    44 => (x"66",x"ec",x"c0",x"bb"),
    45 => (x"c0",x"80",x"c1",x"48"),
    46 => (x"73",x"58",x"a6",x"f0"),
    47 => (x"f0",x"c7",x"02",x"9b"),
    48 => (x"02",x"66",x"c8",x"87"),
    49 => (x"d0",x"87",x"f9",x"c6"),
    50 => (x"78",x"c0",x"48",x"a6"),
    51 => (x"78",x"c0",x"80",x"f8"),
    52 => (x"02",x"ab",x"f0",x"c0"),
    53 => (x"c1",x"87",x"ea",x"c2"),
    54 => (x"c2",x"02",x"ab",x"e3"),
    55 => (x"e4",x"c1",x"87",x"eb"),
    56 => (x"e2",x"c0",x"02",x"ab"),
    57 => (x"ab",x"ec",x"c1",x"87"),
    58 => (x"87",x"d5",x"c2",x"02"),
    59 => (x"02",x"ab",x"f0",x"c1"),
    60 => (x"f3",x"c1",x"87",x"dd"),
    61 => (x"87",x"df",x"02",x"ab"),
    62 => (x"02",x"ab",x"f5",x"c1"),
    63 => (x"f8",x"c1",x"87",x"c9"),
    64 => (x"87",x"cb",x"02",x"ab"),
    65 => (x"d0",x"87",x"e6",x"c2"),
    66 => (x"78",x"ca",x"48",x"a6"),
    67 => (x"d0",x"87",x"fb",x"c2"),
    68 => (x"78",x"d0",x"48",x"a6"),
    69 => (x"c0",x"87",x"f3",x"c2"),
    70 => (x"c4",x"48",x"66",x"f0"),
    71 => (x"a6",x"f4",x"c0",x"80"),
    72 => (x"66",x"f0",x"c0",x"58"),
    73 => (x"76",x"89",x"c4",x"49"),
    74 => (x"d4",x"78",x"69",x"48"),
    75 => (x"6e",x"78",x"ff",x"80"),
    76 => (x"fe",x"48",x"bf",x"97"),
    77 => (x"dc",x"b8",x"80",x"c0"),
    78 => (x"48",x"6e",x"58",x"a6"),
    79 => (x"a6",x"c4",x"80",x"c1"),
    80 => (x"5b",x"a6",x"d0",x"58"),
    81 => (x"c0",x"02",x"66",x"d8"),
    82 => (x"66",x"d8",x"87",x"e8"),
    83 => (x"d4",x"4b",x"6e",x"4c"),
    84 => (x"80",x"c1",x"48",x"66"),
    85 => (x"c0",x"58",x"a6",x"d8"),
    86 => (x"74",x"1e",x"66",x"f8"),
    87 => (x"c8",x"0f",x"75",x"1e"),
    88 => (x"05",x"a8",x"74",x"86"),
    89 => (x"4c",x"13",x"87",x"cc"),
    90 => (x"bc",x"84",x"c0",x"fe"),
    91 => (x"ff",x"05",x"9c",x"74"),
    92 => (x"66",x"cc",x"87",x"dd"),
    93 => (x"48",x"66",x"d4",x"4b"),
    94 => (x"c8",x"80",x"66",x"c4"),
    95 => (x"c9",x"c1",x"58",x"a6"),
    96 => (x"48",x"a6",x"c8",x"87"),
    97 => (x"c1",x"c1",x"78",x"c1"),
    98 => (x"66",x"f8",x"c0",x"87"),
    99 => (x"66",x"f4",x"c0",x"1e"),
   100 => (x"c0",x"80",x"c4",x"48"),
   101 => (x"c0",x"58",x"a6",x"f8"),
   102 => (x"c4",x"49",x"66",x"f4"),
   103 => (x"75",x"1e",x"69",x"89"),
   104 => (x"c4",x"86",x"c8",x"0f"),
   105 => (x"80",x"c1",x"48",x"66"),
   106 => (x"dd",x"58",x"a6",x"c8"),
   107 => (x"66",x"f8",x"c0",x"87"),
   108 => (x"1e",x"e5",x"c0",x"1e"),
   109 => (x"86",x"c8",x"0f",x"75"),
   110 => (x"1e",x"66",x"f8",x"c0"),
   111 => (x"0f",x"75",x"1e",x"73"),
   112 => (x"66",x"c4",x"86",x"c8"),
   113 => (x"c8",x"80",x"c1",x"48"),
   114 => (x"66",x"d0",x"58",x"a6"),
   115 => (x"87",x"c7",x"c3",x"02"),
   116 => (x"48",x"66",x"f0",x"c0"),
   117 => (x"f4",x"c0",x"80",x"c4"),
   118 => (x"f0",x"c0",x"58",x"a6"),
   119 => (x"89",x"c4",x"49",x"66"),
   120 => (x"78",x"69",x"48",x"76"),
   121 => (x"05",x"ab",x"e4",x"c1"),
   122 => (x"48",x"6e",x"87",x"d8"),
   123 => (x"03",x"a8",x"b7",x"c0"),
   124 => (x"ed",x"c0",x"87",x"d0"),
   125 => (x"0f",x"fc",x"c0",x"1e"),
   126 => (x"48",x"6e",x"86",x"c4"),
   127 => (x"c4",x"88",x"08",x"c0"),
   128 => (x"4a",x"6e",x"58",x"a6"),
   129 => (x"4c",x"ea",x"d5",x"c1"),
   130 => (x"c0",x"48",x"a6",x"cc"),
   131 => (x"ce",x"05",x"6e",x"78"),
   132 => (x"eb",x"d5",x"c1",x"87"),
   133 => (x"ea",x"d5",x"c1",x"4c"),
   134 => (x"50",x"f0",x"c0",x"48"),
   135 => (x"6e",x"87",x"eb",x"c0"),
   136 => (x"87",x"e6",x"c0",x"02"),
   137 => (x"72",x"4b",x"66",x"d0"),
   138 => (x"73",x"49",x"72",x"1e"),
   139 => (x"87",x"d7",x"c5",x"4a"),
   140 => (x"f6",x"cd",x"4a",x"26"),
   141 => (x"71",x"54",x"11",x"81"),
   142 => (x"73",x"49",x"72",x"1e"),
   143 => (x"87",x"c7",x"c5",x"4a"),
   144 => (x"49",x"26",x"4a",x"70"),
   145 => (x"ff",x"05",x"9a",x"72"),
   146 => (x"d5",x"c1",x"87",x"dd"),
   147 => (x"c0",x"02",x"ac",x"ea"),
   148 => (x"f8",x"c0",x"87",x"e3"),
   149 => (x"8c",x"c1",x"1e",x"66"),
   150 => (x"fe",x"49",x"6c",x"97"),
   151 => (x"71",x"b9",x"81",x"c0"),
   152 => (x"c8",x"0f",x"75",x"1e"),
   153 => (x"48",x"66",x"cc",x"86"),
   154 => (x"a6",x"d0",x"80",x"c1"),
   155 => (x"ea",x"d5",x"c1",x"58"),
   156 => (x"dd",x"ff",x"05",x"ac"),
   157 => (x"48",x"66",x"cc",x"87"),
   158 => (x"c8",x"80",x"66",x"c4"),
   159 => (x"87",x"d7",x"58",x"a6"),
   160 => (x"05",x"ab",x"e5",x"c0"),
   161 => (x"a6",x"c8",x"87",x"c7"),
   162 => (x"ca",x"78",x"c1",x"48"),
   163 => (x"66",x"f8",x"c0",x"87"),
   164 => (x"75",x"1e",x"73",x"1e"),
   165 => (x"c0",x"86",x"c8",x"0f"),
   166 => (x"bf",x"97",x"66",x"ec"),
   167 => (x"83",x"c0",x"fe",x"4b"),
   168 => (x"66",x"ec",x"c0",x"bb"),
   169 => (x"c0",x"80",x"c1",x"48"),
   170 => (x"73",x"58",x"a6",x"f0"),
   171 => (x"d0",x"f8",x"05",x"9b"),
   172 => (x"48",x"66",x"c4",x"87"),
   173 => (x"4d",x"26",x"8e",x"e4"),
   174 => (x"4b",x"26",x"4c",x"26"),
   175 => (x"c0",x"1e",x"4f",x"26"),
   176 => (x"1e",x"fc",x"c0",x"1e"),
   177 => (x"d0",x"1e",x"66",x"d0"),
   178 => (x"d2",x"c2",x"1e",x"66"),
   179 => (x"26",x"86",x"d0",x"0f"),
   180 => (x"1e",x"c0",x"1e",x"4f"),
   181 => (x"d0",x"1e",x"fc",x"c0"),
   182 => (x"66",x"d0",x"1e",x"a6"),
   183 => (x"0f",x"d2",x"c2",x"1e"),
   184 => (x"4f",x"26",x"86",x"d0"),
   185 => (x"76",x"86",x"f8",x"1e"),
   186 => (x"78",x"66",x"cc",x"48"),
   187 => (x"78",x"ff",x"80",x"c4"),
   188 => (x"c7",x"cd",x"1e",x"76"),
   189 => (x"1e",x"a6",x"dc",x"1e"),
   190 => (x"c2",x"1e",x"66",x"dc"),
   191 => (x"86",x"d0",x"0f",x"d2"),
   192 => (x"4f",x"26",x"8e",x"f8"),
   193 => (x"76",x"86",x"f8",x"1e"),
   194 => (x"78",x"66",x"cc",x"48"),
   195 => (x"66",x"d0",x"80",x"c4"),
   196 => (x"cd",x"1e",x"76",x"78"),
   197 => (x"e0",x"c0",x"1e",x"c7"),
   198 => (x"e0",x"c0",x"1e",x"a6"),
   199 => (x"d2",x"c2",x"1e",x"66"),
   200 => (x"f8",x"86",x"d0",x"0f"),
   201 => (x"1e",x"4f",x"26",x"8e"),
   202 => (x"48",x"76",x"86",x"f8"),
   203 => (x"c4",x"78",x"66",x"cc"),
   204 => (x"76",x"78",x"ff",x"80"),
   205 => (x"1e",x"c7",x"cd",x"1e"),
   206 => (x"dc",x"1e",x"66",x"dc"),
   207 => (x"d2",x"c2",x"1e",x"66"),
   208 => (x"f8",x"86",x"d0",x"0f"),
   209 => (x"1e",x"4f",x"26",x"8e"),
   210 => (x"c4",x"4a",x"66",x"c8"),
   211 => (x"c0",x"02",x"6a",x"82"),
   212 => (x"48",x"6a",x"87",x"e0"),
   213 => (x"7a",x"70",x"88",x"c1"),
   214 => (x"49",x"bf",x"66",x"c8"),
   215 => (x"80",x"c1",x"48",x"71"),
   216 => (x"78",x"08",x"66",x"c8"),
   217 => (x"66",x"c4",x"97",x"08"),
   218 => (x"98",x"ff",x"c3",x"51"),
   219 => (x"c0",x"48",x"66",x"c4"),
   220 => (x"48",x"c0",x"87",x"c2"),
   221 => (x"31",x"30",x"4f",x"26"),
   222 => (x"35",x"34",x"33",x"32"),
   223 => (x"39",x"38",x"37",x"36"),
   224 => (x"44",x"43",x"42",x"41"),
   225 => (x"1e",x"00",x"46",x"45"),
   226 => (x"9a",x"72",x"1e",x"73"),
   227 => (x"87",x"e7",x"c0",x"02"),
   228 => (x"4b",x"c1",x"48",x"c0"),
   229 => (x"d1",x"06",x"a9",x"72"),
   230 => (x"06",x"82",x"72",x"87"),
   231 => (x"83",x"73",x"87",x"c9"),
   232 => (x"f4",x"01",x"a9",x"72"),
   233 => (x"c1",x"87",x"c3",x"87"),
   234 => (x"a9",x"72",x"3a",x"b2"),
   235 => (x"80",x"73",x"89",x"03"),
   236 => (x"2b",x"2a",x"c1",x"07"),
   237 => (x"26",x"87",x"f3",x"05"),
   238 => (x"1e",x"4f",x"26",x"4b"),
   239 => (x"4d",x"c4",x"1e",x"75"),
   240 => (x"04",x"a1",x"b7",x"71"),
   241 => (x"81",x"c1",x"b9",x"ff"),
   242 => (x"72",x"07",x"bd",x"c3"),
   243 => (x"ff",x"04",x"a2",x"b7"),
   244 => (x"c1",x"82",x"c1",x"ba"),
   245 => (x"ee",x"fe",x"07",x"bd"),
   246 => (x"04",x"2d",x"c1",x"87"),
   247 => (x"80",x"c1",x"b8",x"ff"),
   248 => (x"ff",x"04",x"2d",x"07"),
   249 => (x"07",x"81",x"c1",x"b9"),
   250 => (x"4f",x"26",x"4d",x"26"),
   251 => (x"12",x"1e",x"72",x"1e"),
   252 => (x"c4",x"02",x"11",x"48"),
   253 => (x"f6",x"02",x"88",x"87"),
   254 => (x"26",x"4a",x"26",x"87"),
   255 => (x"c8",x"ff",x"1e",x"4f"),
   256 => (x"4f",x"26",x"48",x"bf"),
   257 => (x"5c",x"5b",x"5e",x"0e"),
   258 => (x"dc",x"ff",x"0e",x"5d"),
   259 => (x"fe",x"d5",x"c1",x"86"),
   260 => (x"fc",x"f5",x"c3",x"48"),
   261 => (x"fa",x"d5",x"c1",x"78"),
   262 => (x"ec",x"f6",x"c3",x"48"),
   263 => (x"f5",x"c3",x"48",x"78"),
   264 => (x"f6",x"c3",x"78",x"fc"),
   265 => (x"78",x"c0",x"48",x"f0"),
   266 => (x"78",x"c2",x"80",x"c4"),
   267 => (x"48",x"f8",x"f6",x"c3"),
   268 => (x"71",x"78",x"e8",x"c0"),
   269 => (x"fc",x"f6",x"c3",x"1e"),
   270 => (x"ed",x"f5",x"c0",x"49"),
   271 => (x"20",x"41",x"20",x"48"),
   272 => (x"20",x"41",x"20",x"41"),
   273 => (x"20",x"41",x"20",x"41"),
   274 => (x"10",x"41",x"20",x"41"),
   275 => (x"10",x"51",x"10",x"51"),
   276 => (x"71",x"49",x"26",x"51"),
   277 => (x"dc",x"f7",x"c3",x"1e"),
   278 => (x"cc",x"f6",x"c0",x"49"),
   279 => (x"20",x"41",x"20",x"48"),
   280 => (x"20",x"41",x"20",x"41"),
   281 => (x"20",x"41",x"20",x"41"),
   282 => (x"10",x"41",x"20",x"41"),
   283 => (x"10",x"51",x"10",x"51"),
   284 => (x"c1",x"49",x"26",x"51"),
   285 => (x"ca",x"48",x"f0",x"f2"),
   286 => (x"eb",x"f6",x"c0",x"78"),
   287 => (x"0f",x"d1",x"cb",x"1e"),
   288 => (x"f6",x"c0",x"86",x"c4"),
   289 => (x"d1",x"cb",x"1e",x"ed"),
   290 => (x"c0",x"86",x"c4",x"0f"),
   291 => (x"cb",x"1e",x"dd",x"f7"),
   292 => (x"86",x"c4",x"0f",x"d1"),
   293 => (x"bf",x"ec",x"ef",x"c0"),
   294 => (x"c0",x"87",x"d4",x"02"),
   295 => (x"cb",x"1e",x"f4",x"ef"),
   296 => (x"86",x"c4",x"0f",x"d1"),
   297 => (x"1e",x"e0",x"f0",x"c0"),
   298 => (x"c4",x"0f",x"d1",x"cb"),
   299 => (x"c0",x"87",x"d2",x"86"),
   300 => (x"cb",x"1e",x"e2",x"f0"),
   301 => (x"86",x"c4",x"0f",x"d1"),
   302 => (x"1e",x"d1",x"f1",x"c0"),
   303 => (x"c4",x"0f",x"d1",x"cb"),
   304 => (x"f0",x"ef",x"c0",x"86"),
   305 => (x"f7",x"c0",x"1e",x"bf"),
   306 => (x"d1",x"cb",x"1e",x"df"),
   307 => (x"c3",x"86",x"c8",x"0f"),
   308 => (x"ff",x"48",x"e4",x"f5"),
   309 => (x"c8",x"78",x"bf",x"c8"),
   310 => (x"78",x"c1",x"48",x"a6"),
   311 => (x"bf",x"f0",x"ef",x"c0"),
   312 => (x"a8",x"b7",x"c0",x"48"),
   313 => (x"87",x"de",x"c9",x"06"),
   314 => (x"d4",x"48",x"a6",x"cc"),
   315 => (x"80",x"c8",x"58",x"a6"),
   316 => (x"dc",x"58",x"a6",x"dc"),
   317 => (x"a6",x"c8",x"48",x"a6"),
   318 => (x"ca",x"d6",x"c1",x"58"),
   319 => (x"50",x"c1",x"c1",x"48"),
   320 => (x"48",x"c6",x"d6",x"c1"),
   321 => (x"d6",x"c1",x"78",x"c0"),
   322 => (x"49",x"bf",x"97",x"ca"),
   323 => (x"b9",x"81",x"c0",x"fe"),
   324 => (x"02",x"a9",x"c1",x"c1"),
   325 => (x"76",x"87",x"c7",x"c0"),
   326 => (x"c0",x"78",x"c0",x"48"),
   327 => (x"48",x"76",x"87",x"c4"),
   328 => (x"d6",x"c1",x"78",x"c1"),
   329 => (x"6e",x"48",x"bf",x"c6"),
   330 => (x"ca",x"d6",x"c1",x"b0"),
   331 => (x"cb",x"d6",x"c1",x"58"),
   332 => (x"50",x"c2",x"c1",x"48"),
   333 => (x"c2",x"48",x"a6",x"dc"),
   334 => (x"c3",x"80",x"c4",x"78"),
   335 => (x"fb",x"f7",x"c3",x"78"),
   336 => (x"f2",x"f1",x"c0",x"49"),
   337 => (x"20",x"41",x"20",x"48"),
   338 => (x"20",x"41",x"20",x"41"),
   339 => (x"20",x"41",x"20",x"41"),
   340 => (x"10",x"41",x"20",x"41"),
   341 => (x"10",x"51",x"10",x"51"),
   342 => (x"48",x"a6",x"d4",x"51"),
   343 => (x"f7",x"c3",x"78",x"c1"),
   344 => (x"f7",x"c3",x"1e",x"fb"),
   345 => (x"d3",x"c1",x"1e",x"dc"),
   346 => (x"86",x"c8",x"0f",x"e6"),
   347 => (x"c0",x"05",x"98",x"70"),
   348 => (x"49",x"c1",x"87",x"c5"),
   349 => (x"c0",x"87",x"c2",x"c0"),
   350 => (x"ca",x"d6",x"c1",x"49"),
   351 => (x"48",x"66",x"dc",x"59"),
   352 => (x"03",x"a8",x"b7",x"c3"),
   353 => (x"dc",x"87",x"ef",x"c0"),
   354 => (x"b7",x"c5",x"49",x"66"),
   355 => (x"c3",x"48",x"71",x"91"),
   356 => (x"58",x"a6",x"d0",x"88"),
   357 => (x"c3",x"1e",x"66",x"d0"),
   358 => (x"66",x"e4",x"c0",x"1e"),
   359 => (x"fe",x"cf",x"c1",x"1e"),
   360 => (x"dc",x"86",x"cc",x"0f"),
   361 => (x"80",x"c1",x"48",x"66"),
   362 => (x"58",x"a6",x"e0",x"c0"),
   363 => (x"c3",x"48",x"66",x"dc"),
   364 => (x"ff",x"04",x"a8",x"b7"),
   365 => (x"66",x"cc",x"87",x"d1"),
   366 => (x"66",x"e0",x"c0",x"1e"),
   367 => (x"d4",x"d9",x"c1",x"1e"),
   368 => (x"cc",x"d6",x"c1",x"1e"),
   369 => (x"d0",x"d0",x"c1",x"1e"),
   370 => (x"c1",x"86",x"d0",x"0f"),
   371 => (x"4c",x"bf",x"fa",x"d5"),
   372 => (x"bf",x"fa",x"d5",x"c1"),
   373 => (x"1e",x"72",x"4b",x"bf"),
   374 => (x"d5",x"c1",x"49",x"73"),
   375 => (x"c0",x"48",x"bf",x"fa"),
   376 => (x"20",x"4a",x"a1",x"f0"),
   377 => (x"05",x"aa",x"71",x"41"),
   378 => (x"26",x"87",x"f8",x"ff"),
   379 => (x"c8",x"48",x"74",x"4a"),
   380 => (x"58",x"a6",x"c4",x"80"),
   381 => (x"81",x"cc",x"49",x"74"),
   382 => (x"4d",x"73",x"79",x"c5"),
   383 => (x"7d",x"69",x"85",x"cc"),
   384 => (x"1e",x"73",x"7b",x"6c"),
   385 => (x"0f",x"c2",x"ef",x"c0"),
   386 => (x"49",x"73",x"86",x"c4"),
   387 => (x"05",x"69",x"81",x"c4"),
   388 => (x"73",x"87",x"e7",x"c0"),
   389 => (x"c6",x"81",x"c8",x"49"),
   390 => (x"c4",x"1e",x"71",x"7d"),
   391 => (x"c1",x"1e",x"bf",x"66"),
   392 => (x"c8",x"0f",x"d0",x"ce"),
   393 => (x"fa",x"d5",x"c1",x"86"),
   394 => (x"75",x"7b",x"bf",x"bf"),
   395 => (x"6d",x"1e",x"ca",x"1e"),
   396 => (x"fe",x"cf",x"c1",x"1e"),
   397 => (x"c0",x"86",x"cc",x"0f"),
   398 => (x"49",x"6c",x"87",x"d9"),
   399 => (x"1e",x"72",x"1e",x"71"),
   400 => (x"c0",x"48",x"49",x"74"),
   401 => (x"20",x"4a",x"a1",x"f0"),
   402 => (x"05",x"aa",x"71",x"41"),
   403 => (x"26",x"87",x"f8",x"ff"),
   404 => (x"76",x"49",x"26",x"4a"),
   405 => (x"50",x"c1",x"c1",x"48"),
   406 => (x"97",x"cb",x"d6",x"c1"),
   407 => (x"c0",x"fe",x"49",x"bf"),
   408 => (x"c1",x"c1",x"b9",x"81"),
   409 => (x"c1",x"04",x"a9",x"b7"),
   410 => (x"6e",x"97",x"87",x"ed"),
   411 => (x"1e",x"c3",x"c1",x"4b"),
   412 => (x"c0",x"fe",x"49",x"73"),
   413 => (x"1e",x"71",x"b9",x"81"),
   414 => (x"0f",x"fb",x"d2",x"c1"),
   415 => (x"66",x"d4",x"86",x"c8"),
   416 => (x"f9",x"c0",x"05",x"a8"),
   417 => (x"1e",x"66",x"d8",x"87"),
   418 => (x"ce",x"c1",x"1e",x"c0"),
   419 => (x"86",x"c8",x"0f",x"d0"),
   420 => (x"f7",x"c3",x"1e",x"71"),
   421 => (x"f1",x"c0",x"49",x"fb"),
   422 => (x"41",x"20",x"48",x"d3"),
   423 => (x"41",x"20",x"41",x"20"),
   424 => (x"41",x"20",x"41",x"20"),
   425 => (x"41",x"20",x"41",x"20"),
   426 => (x"51",x"10",x"51",x"10"),
   427 => (x"49",x"26",x"51",x"10"),
   428 => (x"48",x"a6",x"e0",x"c0"),
   429 => (x"c1",x"78",x"66",x"c8"),
   430 => (x"c8",x"48",x"c2",x"d6"),
   431 => (x"83",x"c1",x"78",x"66"),
   432 => (x"c0",x"fe",x"4a",x"73"),
   433 => (x"d6",x"c1",x"ba",x"82"),
   434 => (x"49",x"bf",x"97",x"cb"),
   435 => (x"b9",x"81",x"c0",x"fe"),
   436 => (x"06",x"aa",x"b7",x"71"),
   437 => (x"c0",x"87",x"d6",x"fe"),
   438 => (x"dc",x"48",x"66",x"e0"),
   439 => (x"c0",x"90",x"b7",x"66"),
   440 => (x"71",x"58",x"a6",x"e4"),
   441 => (x"c0",x"1e",x"72",x"1e"),
   442 => (x"d4",x"49",x"66",x"e8"),
   443 => (x"ca",x"f3",x"4a",x"66"),
   444 => (x"26",x"4a",x"26",x"87"),
   445 => (x"a6",x"e0",x"c0",x"49"),
   446 => (x"66",x"e0",x"c0",x"58"),
   447 => (x"89",x"66",x"cc",x"49"),
   448 => (x"71",x"91",x"b7",x"c7"),
   449 => (x"88",x"66",x"dc",x"48"),
   450 => (x"58",x"a6",x"e4",x"c0"),
   451 => (x"4a",x"bf",x"66",x"c4"),
   452 => (x"d6",x"c1",x"82",x"ca"),
   453 => (x"49",x"bf",x"97",x"ca"),
   454 => (x"b9",x"81",x"c0",x"fe"),
   455 => (x"05",x"a9",x"c1",x"c1"),
   456 => (x"c1",x"87",x"ce",x"c0"),
   457 => (x"c1",x"48",x"72",x"8a"),
   458 => (x"88",x"bf",x"c2",x"d6"),
   459 => (x"78",x"08",x"66",x"c4"),
   460 => (x"48",x"66",x"c8",x"08"),
   461 => (x"a6",x"cc",x"80",x"c1"),
   462 => (x"48",x"66",x"c8",x"58"),
   463 => (x"bf",x"f0",x"ef",x"c0"),
   464 => (x"f6",x"06",x"a8",x"b7"),
   465 => (x"f5",x"c3",x"87",x"f3"),
   466 => (x"c8",x"ff",x"48",x"e8"),
   467 => (x"f8",x"c0",x"78",x"bf"),
   468 => (x"d1",x"cb",x"1e",x"cc"),
   469 => (x"c0",x"86",x"c4",x"0f"),
   470 => (x"cb",x"1e",x"dc",x"f8"),
   471 => (x"86",x"c4",x"0f",x"d1"),
   472 => (x"1e",x"de",x"f8",x"c0"),
   473 => (x"c4",x"0f",x"d1",x"cb"),
   474 => (x"d4",x"f9",x"c0",x"86"),
   475 => (x"0f",x"d1",x"cb",x"1e"),
   476 => (x"d6",x"c1",x"86",x"c4"),
   477 => (x"c0",x"1e",x"bf",x"c2"),
   478 => (x"cb",x"1e",x"d6",x"f9"),
   479 => (x"86",x"c8",x"0f",x"d1"),
   480 => (x"f9",x"c0",x"1e",x"c5"),
   481 => (x"d1",x"cb",x"1e",x"ef"),
   482 => (x"c1",x"86",x"c8",x"0f"),
   483 => (x"1e",x"bf",x"c6",x"d6"),
   484 => (x"1e",x"c8",x"fa",x"c0"),
   485 => (x"c8",x"0f",x"d1",x"cb"),
   486 => (x"c0",x"1e",x"c1",x"86"),
   487 => (x"cb",x"1e",x"e1",x"fa"),
   488 => (x"86",x"c8",x"0f",x"d1"),
   489 => (x"97",x"ca",x"d6",x"c1"),
   490 => (x"c0",x"fe",x"49",x"bf"),
   491 => (x"1e",x"71",x"b9",x"81"),
   492 => (x"1e",x"fa",x"fa",x"c0"),
   493 => (x"c8",x"0f",x"d1",x"cb"),
   494 => (x"1e",x"c1",x"c1",x"86"),
   495 => (x"1e",x"d3",x"fb",x"c0"),
   496 => (x"c8",x"0f",x"d1",x"cb"),
   497 => (x"cb",x"d6",x"c1",x"86"),
   498 => (x"fe",x"49",x"bf",x"97"),
   499 => (x"71",x"b9",x"81",x"c0"),
   500 => (x"ec",x"fb",x"c0",x"1e"),
   501 => (x"0f",x"d1",x"cb",x"1e"),
   502 => (x"c2",x"c1",x"86",x"c8"),
   503 => (x"c5",x"fc",x"c0",x"1e"),
   504 => (x"0f",x"d1",x"cb",x"1e"),
   505 => (x"d6",x"c1",x"86",x"c8"),
   506 => (x"c0",x"1e",x"bf",x"ec"),
   507 => (x"cb",x"1e",x"de",x"fc"),
   508 => (x"86",x"c8",x"0f",x"d1"),
   509 => (x"fc",x"c0",x"1e",x"c7"),
   510 => (x"d1",x"cb",x"1e",x"f7"),
   511 => (x"c1",x"86",x"c8",x"0f"),
   512 => (x"1e",x"bf",x"f0",x"f2"),
   513 => (x"1e",x"d0",x"fd",x"c0"),
   514 => (x"c8",x"0f",x"d1",x"cb"),
   515 => (x"e9",x"fd",x"c0",x"86"),
   516 => (x"0f",x"d1",x"cb",x"1e"),
   517 => (x"fe",x"c0",x"86",x"c4"),
   518 => (x"d1",x"cb",x"1e",x"d3"),
   519 => (x"c1",x"86",x"c4",x"0f"),
   520 => (x"bf",x"bf",x"fa",x"d5"),
   521 => (x"df",x"fe",x"c0",x"1e"),
   522 => (x"0f",x"d1",x"cb",x"1e"),
   523 => (x"fe",x"c0",x"86",x"c8"),
   524 => (x"d1",x"cb",x"1e",x"f8"),
   525 => (x"c1",x"86",x"c4",x"0f"),
   526 => (x"49",x"bf",x"fa",x"d5"),
   527 => (x"1e",x"69",x"81",x"c4"),
   528 => (x"1e",x"e9",x"ff",x"c0"),
   529 => (x"c8",x"0f",x"d1",x"cb"),
   530 => (x"c1",x"1e",x"c0",x"86"),
   531 => (x"cb",x"1e",x"c2",x"c0"),
   532 => (x"86",x"c8",x"0f",x"d1"),
   533 => (x"bf",x"fa",x"d5",x"c1"),
   534 => (x"69",x"81",x"c8",x"49"),
   535 => (x"db",x"c0",x"c1",x"1e"),
   536 => (x"0f",x"d1",x"cb",x"1e"),
   537 => (x"1e",x"c2",x"86",x"c8"),
   538 => (x"1e",x"f4",x"c0",x"c1"),
   539 => (x"c8",x"0f",x"d1",x"cb"),
   540 => (x"fa",x"d5",x"c1",x"86"),
   541 => (x"81",x"cc",x"49",x"bf"),
   542 => (x"c1",x"c1",x"1e",x"69"),
   543 => (x"d1",x"cb",x"1e",x"cd"),
   544 => (x"d1",x"86",x"c8",x"0f"),
   545 => (x"e6",x"c1",x"c1",x"1e"),
   546 => (x"0f",x"d1",x"cb",x"1e"),
   547 => (x"d5",x"c1",x"86",x"c8"),
   548 => (x"d0",x"49",x"bf",x"fa"),
   549 => (x"c1",x"1e",x"71",x"81"),
   550 => (x"cb",x"1e",x"ff",x"c1"),
   551 => (x"86",x"c8",x"0f",x"d1"),
   552 => (x"1e",x"d8",x"c2",x"c1"),
   553 => (x"c4",x"0f",x"d1",x"cb"),
   554 => (x"cd",x"c3",x"c1",x"86"),
   555 => (x"0f",x"d1",x"cb",x"1e"),
   556 => (x"d5",x"c1",x"86",x"c4"),
   557 => (x"1e",x"bf",x"bf",x"fe"),
   558 => (x"1e",x"de",x"c3",x"c1"),
   559 => (x"c8",x"0f",x"d1",x"cb"),
   560 => (x"f7",x"c3",x"c1",x"86"),
   561 => (x"0f",x"d1",x"cb",x"1e"),
   562 => (x"d5",x"c1",x"86",x"c4"),
   563 => (x"c4",x"49",x"bf",x"fe"),
   564 => (x"c1",x"1e",x"69",x"81"),
   565 => (x"cb",x"1e",x"f7",x"c4"),
   566 => (x"86",x"c8",x"0f",x"d1"),
   567 => (x"c5",x"c1",x"1e",x"c0"),
   568 => (x"d1",x"cb",x"1e",x"d0"),
   569 => (x"c1",x"86",x"c8",x"0f"),
   570 => (x"49",x"bf",x"fe",x"d5"),
   571 => (x"1e",x"69",x"81",x"c8"),
   572 => (x"1e",x"e9",x"c5",x"c1"),
   573 => (x"c8",x"0f",x"d1",x"cb"),
   574 => (x"c1",x"1e",x"c1",x"86"),
   575 => (x"cb",x"1e",x"c2",x"c6"),
   576 => (x"86",x"c8",x"0f",x"d1"),
   577 => (x"bf",x"fe",x"d5",x"c1"),
   578 => (x"69",x"81",x"cc",x"49"),
   579 => (x"db",x"c6",x"c1",x"1e"),
   580 => (x"0f",x"d1",x"cb",x"1e"),
   581 => (x"1e",x"d2",x"86",x"c8"),
   582 => (x"1e",x"f4",x"c6",x"c1"),
   583 => (x"c8",x"0f",x"d1",x"cb"),
   584 => (x"fe",x"d5",x"c1",x"86"),
   585 => (x"81",x"d0",x"49",x"bf"),
   586 => (x"c7",x"c1",x"1e",x"71"),
   587 => (x"d1",x"cb",x"1e",x"cd"),
   588 => (x"c1",x"86",x"c8",x"0f"),
   589 => (x"cb",x"1e",x"e6",x"c7"),
   590 => (x"86",x"c4",x"0f",x"d1"),
   591 => (x"c1",x"1e",x"66",x"dc"),
   592 => (x"cb",x"1e",x"db",x"c8"),
   593 => (x"86",x"c8",x"0f",x"d1"),
   594 => (x"c8",x"c1",x"1e",x"c5"),
   595 => (x"d1",x"cb",x"1e",x"f4"),
   596 => (x"c0",x"86",x"c8",x"0f"),
   597 => (x"c1",x"1e",x"66",x"e0"),
   598 => (x"cb",x"1e",x"cd",x"c9"),
   599 => (x"86",x"c8",x"0f",x"d1"),
   600 => (x"c9",x"c1",x"1e",x"cd"),
   601 => (x"d1",x"cb",x"1e",x"e6"),
   602 => (x"cc",x"86",x"c8",x"0f"),
   603 => (x"c9",x"c1",x"1e",x"66"),
   604 => (x"d1",x"cb",x"1e",x"ff"),
   605 => (x"c7",x"86",x"c8",x"0f"),
   606 => (x"d8",x"ca",x"c1",x"1e"),
   607 => (x"0f",x"d1",x"cb",x"1e"),
   608 => (x"66",x"d4",x"86",x"c8"),
   609 => (x"f1",x"ca",x"c1",x"1e"),
   610 => (x"0f",x"d1",x"cb",x"1e"),
   611 => (x"1e",x"c1",x"86",x"c8"),
   612 => (x"1e",x"ca",x"cb",x"c1"),
   613 => (x"c8",x"0f",x"d1",x"cb"),
   614 => (x"dc",x"f7",x"c3",x"86"),
   615 => (x"e3",x"cb",x"c1",x"1e"),
   616 => (x"0f",x"d1",x"cb",x"1e"),
   617 => (x"cb",x"c1",x"86",x"c8"),
   618 => (x"d1",x"cb",x"1e",x"fc"),
   619 => (x"c3",x"86",x"c4",x"0f"),
   620 => (x"c1",x"1e",x"fb",x"f7"),
   621 => (x"cb",x"1e",x"f1",x"cc"),
   622 => (x"86",x"c8",x"0f",x"d1"),
   623 => (x"1e",x"ca",x"cd",x"c1"),
   624 => (x"c4",x"0f",x"d1",x"cb"),
   625 => (x"ff",x"cd",x"c1",x"86"),
   626 => (x"0f",x"d1",x"cb",x"1e"),
   627 => (x"f5",x"c3",x"86",x"c4"),
   628 => (x"c3",x"49",x"bf",x"e8"),
   629 => (x"89",x"bf",x"e4",x"f5"),
   630 => (x"59",x"f0",x"f5",x"c3"),
   631 => (x"ce",x"c1",x"1e",x"71"),
   632 => (x"d1",x"cb",x"1e",x"c1"),
   633 => (x"c3",x"86",x"c8",x"0f"),
   634 => (x"48",x"bf",x"ec",x"f5"),
   635 => (x"a8",x"b7",x"f8",x"c1"),
   636 => (x"87",x"db",x"c0",x"03"),
   637 => (x"1e",x"d1",x"f2",x"c0"),
   638 => (x"c4",x"0f",x"d1",x"cb"),
   639 => (x"c7",x"f3",x"c0",x"86"),
   640 => (x"0f",x"d1",x"cb",x"1e"),
   641 => (x"f3",x"c0",x"86",x"c4"),
   642 => (x"d1",x"cb",x"1e",x"e7"),
   643 => (x"c3",x"86",x"c4",x"0f"),
   644 => (x"49",x"bf",x"ec",x"f5"),
   645 => (x"e8",x"cf",x"4a",x"71"),
   646 => (x"1e",x"71",x"92",x"b7"),
   647 => (x"49",x"72",x"1e",x"72"),
   648 => (x"bf",x"f0",x"ef",x"c0"),
   649 => (x"87",x"d3",x"e6",x"4a"),
   650 => (x"49",x"26",x"4a",x"26"),
   651 => (x"58",x"f4",x"f5",x"c3"),
   652 => (x"bf",x"f0",x"ef",x"c0"),
   653 => (x"cf",x"4b",x"72",x"4a"),
   654 => (x"71",x"93",x"b7",x"e8"),
   655 => (x"73",x"1e",x"72",x"1e"),
   656 => (x"f6",x"e5",x"4a",x"09"),
   657 => (x"26",x"4a",x"26",x"87"),
   658 => (x"f8",x"f5",x"c3",x"49"),
   659 => (x"b7",x"f9",x"c8",x"58"),
   660 => (x"72",x"1e",x"71",x"92"),
   661 => (x"4a",x"09",x"72",x"1e"),
   662 => (x"26",x"87",x"e0",x"e5"),
   663 => (x"c3",x"49",x"26",x"4a"),
   664 => (x"c0",x"58",x"fc",x"f5"),
   665 => (x"cb",x"1e",x"e9",x"f3"),
   666 => (x"86",x"c4",x"0f",x"d1"),
   667 => (x"bf",x"f0",x"f5",x"c3"),
   668 => (x"d6",x"f4",x"c0",x"1e"),
   669 => (x"0f",x"d1",x"cb",x"1e"),
   670 => (x"f4",x"c0",x"86",x"c8"),
   671 => (x"d1",x"cb",x"1e",x"db"),
   672 => (x"c3",x"86",x"c4",x"0f"),
   673 => (x"1e",x"bf",x"f4",x"f5"),
   674 => (x"1e",x"c8",x"f5",x"c0"),
   675 => (x"c8",x"0f",x"d1",x"cb"),
   676 => (x"f8",x"f5",x"c3",x"86"),
   677 => (x"f5",x"c0",x"1e",x"bf"),
   678 => (x"d1",x"cb",x"1e",x"cd"),
   679 => (x"c0",x"86",x"c8",x"0f"),
   680 => (x"cb",x"1e",x"eb",x"f5"),
   681 => (x"86",x"c4",x"0f",x"d1"),
   682 => (x"dc",x"ff",x"48",x"c0"),
   683 => (x"26",x"4d",x"26",x"8e"),
   684 => (x"26",x"4b",x"26",x"4c"),
   685 => (x"d6",x"c1",x"1e",x"4f"),
   686 => (x"c1",x"c1",x"48",x"ca"),
   687 => (x"c6",x"d6",x"c1",x"50"),
   688 => (x"26",x"78",x"c0",x"48"),
   689 => (x"d6",x"c1",x"1e",x"4f"),
   690 => (x"49",x"bf",x"97",x"ca"),
   691 => (x"b9",x"81",x"c0",x"fe"),
   692 => (x"02",x"a9",x"c1",x"c1"),
   693 => (x"c0",x"87",x"c5",x"c0"),
   694 => (x"87",x"c2",x"c0",x"49"),
   695 => (x"d6",x"c1",x"49",x"c1"),
   696 => (x"71",x"48",x"bf",x"c6"),
   697 => (x"ca",x"d6",x"c1",x"b0"),
   698 => (x"cb",x"d6",x"c1",x"58"),
   699 => (x"50",x"c2",x"c1",x"48"),
   700 => (x"5e",x"0e",x"4f",x"26"),
   701 => (x"0e",x"5d",x"5c",x"5b"),
   702 => (x"66",x"d4",x"86",x"fc"),
   703 => (x"73",x"4b",x"6d",x"4d"),
   704 => (x"fa",x"d5",x"c1",x"49"),
   705 => (x"f0",x"c0",x"48",x"bf"),
   706 => (x"41",x"20",x"4a",x"a1"),
   707 => (x"ff",x"05",x"aa",x"71"),
   708 => (x"48",x"75",x"87",x"f8"),
   709 => (x"a6",x"c4",x"80",x"c8"),
   710 => (x"cc",x"49",x"75",x"58"),
   711 => (x"73",x"79",x"c5",x"81"),
   712 => (x"c5",x"84",x"cc",x"4c"),
   713 => (x"c1",x"7b",x"6d",x"7c"),
   714 => (x"02",x"bf",x"fa",x"d5"),
   715 => (x"c1",x"87",x"c6",x"c0"),
   716 => (x"bf",x"bf",x"fa",x"d5"),
   717 => (x"fa",x"d5",x"c1",x"7b"),
   718 => (x"81",x"cc",x"49",x"bf"),
   719 => (x"d6",x"c1",x"1e",x"71"),
   720 => (x"ca",x"1e",x"bf",x"c2"),
   721 => (x"fe",x"cf",x"c1",x"1e"),
   722 => (x"73",x"86",x"cc",x"0f"),
   723 => (x"69",x"81",x"c4",x"49"),
   724 => (x"87",x"e7",x"c0",x"05"),
   725 => (x"81",x"c8",x"49",x"73"),
   726 => (x"1e",x"71",x"7c",x"c6"),
   727 => (x"1e",x"bf",x"66",x"c4"),
   728 => (x"0f",x"d0",x"ce",x"c1"),
   729 => (x"d5",x"c1",x"86",x"c8"),
   730 => (x"7b",x"bf",x"bf",x"fa"),
   731 => (x"1e",x"ca",x"1e",x"74"),
   732 => (x"cf",x"c1",x"1e",x"6c"),
   733 => (x"86",x"cc",x"0f",x"fe"),
   734 => (x"6d",x"87",x"d5",x"c0"),
   735 => (x"75",x"1e",x"71",x"49"),
   736 => (x"f0",x"c0",x"48",x"49"),
   737 => (x"41",x"20",x"4a",x"a1"),
   738 => (x"ff",x"05",x"aa",x"71"),
   739 => (x"49",x"26",x"87",x"f8"),
   740 => (x"4d",x"26",x"8e",x"fc"),
   741 => (x"4b",x"26",x"4c",x"26"),
   742 => (x"c4",x"1e",x"4f",x"26"),
   743 => (x"ca",x"4a",x"bf",x"66"),
   744 => (x"ca",x"d6",x"c1",x"82"),
   745 => (x"fe",x"49",x"bf",x"97"),
   746 => (x"c1",x"b9",x"81",x"c0"),
   747 => (x"c0",x"05",x"a9",x"c1"),
   748 => (x"8a",x"c1",x"87",x"ce"),
   749 => (x"d6",x"c1",x"48",x"72"),
   750 => (x"c4",x"88",x"bf",x"c2"),
   751 => (x"08",x"78",x"08",x"66"),
   752 => (x"c1",x"1e",x"4f",x"26"),
   753 => (x"02",x"bf",x"fa",x"d5"),
   754 => (x"c4",x"87",x"c9",x"c0"),
   755 => (x"d5",x"c1",x"48",x"66"),
   756 => (x"78",x"bf",x"bf",x"fa"),
   757 => (x"bf",x"fa",x"d5",x"c1"),
   758 => (x"71",x"81",x"cc",x"49"),
   759 => (x"c2",x"d6",x"c1",x"1e"),
   760 => (x"1e",x"ca",x"1e",x"bf"),
   761 => (x"0f",x"fe",x"cf",x"c1"),
   762 => (x"4f",x"26",x"86",x"cc"),
   763 => (x"00",x"00",x"00",x"00"),
   764 => (x"00",x"00",x"61",x"a8"),
   765 => (x"67",x"6f",x"72",x"50"),
   766 => (x"20",x"6d",x"61",x"72"),
   767 => (x"70",x"6d",x"6f",x"63"),
   768 => (x"64",x"65",x"6c",x"69"),
   769 => (x"74",x"69",x"77",x"20"),
   770 => (x"72",x"27",x"20",x"68"),
   771 => (x"73",x"69",x"67",x"65"),
   772 => (x"27",x"72",x"65",x"74"),
   773 => (x"74",x"74",x"61",x"20"),
   774 => (x"75",x"62",x"69",x"72"),
   775 => (x"00",x"0a",x"65",x"74"),
   776 => (x"72",x"50",x"00",x"0a"),
   777 => (x"61",x"72",x"67",x"6f"),
   778 => (x"6f",x"63",x"20",x"6d"),
   779 => (x"6c",x"69",x"70",x"6d"),
   780 => (x"77",x"20",x"64",x"65"),
   781 => (x"6f",x"68",x"74",x"69"),
   782 => (x"27",x"20",x"74",x"75"),
   783 => (x"69",x"67",x"65",x"72"),
   784 => (x"72",x"65",x"74",x"73"),
   785 => (x"74",x"61",x"20",x"27"),
   786 => (x"62",x"69",x"72",x"74"),
   787 => (x"0a",x"65",x"74",x"75"),
   788 => (x"44",x"00",x"0a",x"00"),
   789 => (x"53",x"59",x"52",x"48"),
   790 => (x"45",x"4e",x"4f",x"54"),
   791 => (x"4f",x"52",x"50",x"20"),
   792 => (x"4d",x"41",x"52",x"47"),
   793 => (x"27",x"33",x"20",x"2c"),
   794 => (x"53",x"20",x"44",x"52"),
   795 => (x"4e",x"49",x"52",x"54"),
   796 => (x"48",x"44",x"00",x"47"),
   797 => (x"54",x"53",x"59",x"52"),
   798 => (x"20",x"45",x"4e",x"4f"),
   799 => (x"47",x"4f",x"52",x"50"),
   800 => (x"2c",x"4d",x"41",x"52"),
   801 => (x"4e",x"27",x"32",x"20"),
   802 => (x"54",x"53",x"20",x"44"),
   803 => (x"47",x"4e",x"49",x"52"),
   804 => (x"61",x"65",x"4d",x"00"),
   805 => (x"65",x"72",x"75",x"73"),
   806 => (x"69",x"74",x"20",x"64"),
   807 => (x"74",x"20",x"65",x"6d"),
   808 => (x"73",x"20",x"6f",x"6f"),
   809 => (x"6c",x"6c",x"61",x"6d"),
   810 => (x"20",x"6f",x"74",x"20"),
   811 => (x"61",x"74",x"62",x"6f"),
   812 => (x"6d",x"20",x"6e",x"69"),
   813 => (x"69",x"6e",x"61",x"65"),
   814 => (x"75",x"66",x"67",x"6e"),
   815 => (x"65",x"72",x"20",x"6c"),
   816 => (x"74",x"6c",x"75",x"73"),
   817 => (x"50",x"00",x"0a",x"73"),
   818 => (x"73",x"61",x"65",x"6c"),
   819 => (x"6e",x"69",x"20",x"65"),
   820 => (x"61",x"65",x"72",x"63"),
   821 => (x"6e",x"20",x"65",x"73"),
   822 => (x"65",x"62",x"6d",x"75"),
   823 => (x"66",x"6f",x"20",x"72"),
   824 => (x"6e",x"75",x"72",x"20"),
   825 => (x"0a",x"00",x"0a",x"73"),
   826 => (x"63",x"69",x"4d",x"00"),
   827 => (x"65",x"73",x"6f",x"72"),
   828 => (x"64",x"6e",x"6f",x"63"),
   829 => (x"6f",x"66",x"20",x"73"),
   830 => (x"6e",x"6f",x"20",x"72"),
   831 => (x"75",x"72",x"20",x"65"),
   832 => (x"68",x"74",x"20",x"6e"),
   833 => (x"67",x"75",x"6f",x"72"),
   834 => (x"68",x"44",x"20",x"68"),
   835 => (x"74",x"73",x"79",x"72"),
   836 => (x"3a",x"65",x"6e",x"6f"),
   837 => (x"64",x"25",x"00",x"20"),
   838 => (x"44",x"00",x"0a",x"20"),
   839 => (x"73",x"79",x"72",x"68"),
   840 => (x"65",x"6e",x"6f",x"74"),
   841 => (x"65",x"70",x"20",x"73"),
   842 => (x"65",x"53",x"20",x"72"),
   843 => (x"64",x"6e",x"6f",x"63"),
   844 => (x"20",x"20",x"20",x"3a"),
   845 => (x"20",x"20",x"20",x"20"),
   846 => (x"20",x"20",x"20",x"20"),
   847 => (x"20",x"20",x"20",x"20"),
   848 => (x"20",x"20",x"20",x"20"),
   849 => (x"00",x"20",x"20",x"20"),
   850 => (x"0a",x"20",x"64",x"25"),
   851 => (x"58",x"41",x"56",x"00"),
   852 => (x"50",x"49",x"4d",x"20"),
   853 => (x"61",x"72",x"20",x"53"),
   854 => (x"67",x"6e",x"69",x"74"),
   855 => (x"31",x"20",x"2a",x"20"),
   856 => (x"20",x"30",x"30",x"30"),
   857 => (x"64",x"25",x"20",x"3d"),
   858 => (x"0a",x"00",x"0a",x"20"),
   859 => (x"52",x"48",x"44",x"00"),
   860 => (x"4f",x"54",x"53",x"59"),
   861 => (x"50",x"20",x"45",x"4e"),
   862 => (x"52",x"47",x"4f",x"52"),
   863 => (x"20",x"2c",x"4d",x"41"),
   864 => (x"45",x"4d",x"4f",x"53"),
   865 => (x"52",x"54",x"53",x"20"),
   866 => (x"00",x"47",x"4e",x"49"),
   867 => (x"59",x"52",x"48",x"44"),
   868 => (x"4e",x"4f",x"54",x"53"),
   869 => (x"52",x"50",x"20",x"45"),
   870 => (x"41",x"52",x"47",x"4f"),
   871 => (x"31",x"20",x"2c",x"4d"),
   872 => (x"20",x"54",x"53",x"27"),
   873 => (x"49",x"52",x"54",x"53"),
   874 => (x"0a",x"00",x"47",x"4e"),
   875 => (x"72",x"68",x"44",x"00"),
   876 => (x"6f",x"74",x"73",x"79"),
   877 => (x"42",x"20",x"65",x"6e"),
   878 => (x"68",x"63",x"6e",x"65"),
   879 => (x"6b",x"72",x"61",x"6d"),
   880 => (x"65",x"56",x"20",x"2c"),
   881 => (x"6f",x"69",x"73",x"72"),
   882 => (x"2e",x"32",x"20",x"6e"),
   883 => (x"4c",x"28",x"20",x"31"),
   884 => (x"75",x"67",x"6e",x"61"),
   885 => (x"3a",x"65",x"67",x"61"),
   886 => (x"0a",x"29",x"43",x"20"),
   887 => (x"45",x"00",x"0a",x"00"),
   888 => (x"75",x"63",x"65",x"78"),
   889 => (x"6e",x"6f",x"69",x"74"),
   890 => (x"61",x"74",x"73",x"20"),
   891 => (x"2c",x"73",x"74",x"72"),
   892 => (x"20",x"64",x"25",x"20"),
   893 => (x"73",x"6e",x"75",x"72"),
   894 => (x"72",x"68",x"74",x"20"),
   895 => (x"68",x"67",x"75",x"6f"),
   896 => (x"72",x"68",x"44",x"20"),
   897 => (x"6f",x"74",x"73",x"79"),
   898 => (x"00",x"0a",x"65",x"6e"),
   899 => (x"63",x"65",x"78",x"45"),
   900 => (x"6f",x"69",x"74",x"75"),
   901 => (x"6e",x"65",x"20",x"6e"),
   902 => (x"00",x"0a",x"73",x"64"),
   903 => (x"69",x"46",x"00",x"0a"),
   904 => (x"20",x"6c",x"61",x"6e"),
   905 => (x"75",x"6c",x"61",x"76"),
   906 => (x"6f",x"20",x"73",x"65"),
   907 => (x"68",x"74",x"20",x"66"),
   908 => (x"61",x"76",x"20",x"65"),
   909 => (x"62",x"61",x"69",x"72"),
   910 => (x"20",x"73",x"65",x"6c"),
   911 => (x"64",x"65",x"73",x"75"),
   912 => (x"20",x"6e",x"69",x"20"),
   913 => (x"20",x"65",x"68",x"74"),
   914 => (x"63",x"6e",x"65",x"62"),
   915 => (x"72",x"61",x"6d",x"68"),
   916 => (x"00",x"0a",x"3a",x"6b"),
   917 => (x"6e",x"49",x"00",x"0a"),
   918 => (x"6c",x"47",x"5f",x"74"),
   919 => (x"20",x"3a",x"62",x"6f"),
   920 => (x"20",x"20",x"20",x"20"),
   921 => (x"20",x"20",x"20",x"20"),
   922 => (x"25",x"20",x"20",x"20"),
   923 => (x"20",x"00",x"0a",x"64"),
   924 => (x"20",x"20",x"20",x"20"),
   925 => (x"73",x"20",x"20",x"20"),
   926 => (x"6c",x"75",x"6f",x"68"),
   927 => (x"65",x"62",x"20",x"64"),
   928 => (x"20",x"20",x"20",x"3a"),
   929 => (x"00",x"0a",x"64",x"25"),
   930 => (x"6c",x"6f",x"6f",x"42"),
   931 => (x"6f",x"6c",x"47",x"5f"),
   932 => (x"20",x"20",x"3a",x"62"),
   933 => (x"20",x"20",x"20",x"20"),
   934 => (x"20",x"20",x"20",x"20"),
   935 => (x"0a",x"64",x"25",x"20"),
   936 => (x"20",x"20",x"20",x"00"),
   937 => (x"20",x"20",x"20",x"20"),
   938 => (x"6f",x"68",x"73",x"20"),
   939 => (x"20",x"64",x"6c",x"75"),
   940 => (x"20",x"3a",x"65",x"62"),
   941 => (x"64",x"25",x"20",x"20"),
   942 => (x"68",x"43",x"00",x"0a"),
   943 => (x"47",x"5f",x"31",x"5f"),
   944 => (x"3a",x"62",x"6f",x"6c"),
   945 => (x"20",x"20",x"20",x"20"),
   946 => (x"20",x"20",x"20",x"20"),
   947 => (x"25",x"20",x"20",x"20"),
   948 => (x"20",x"00",x"0a",x"63"),
   949 => (x"20",x"20",x"20",x"20"),
   950 => (x"73",x"20",x"20",x"20"),
   951 => (x"6c",x"75",x"6f",x"68"),
   952 => (x"65",x"62",x"20",x"64"),
   953 => (x"20",x"20",x"20",x"3a"),
   954 => (x"00",x"0a",x"63",x"25"),
   955 => (x"32",x"5f",x"68",x"43"),
   956 => (x"6f",x"6c",x"47",x"5f"),
   957 => (x"20",x"20",x"3a",x"62"),
   958 => (x"20",x"20",x"20",x"20"),
   959 => (x"20",x"20",x"20",x"20"),
   960 => (x"0a",x"63",x"25",x"20"),
   961 => (x"20",x"20",x"20",x"00"),
   962 => (x"20",x"20",x"20",x"20"),
   963 => (x"6f",x"68",x"73",x"20"),
   964 => (x"20",x"64",x"6c",x"75"),
   965 => (x"20",x"3a",x"65",x"62"),
   966 => (x"63",x"25",x"20",x"20"),
   967 => (x"72",x"41",x"00",x"0a"),
   968 => (x"5f",x"31",x"5f",x"72"),
   969 => (x"62",x"6f",x"6c",x"47"),
   970 => (x"3a",x"5d",x"38",x"5b"),
   971 => (x"20",x"20",x"20",x"20"),
   972 => (x"25",x"20",x"20",x"20"),
   973 => (x"20",x"00",x"0a",x"64"),
   974 => (x"20",x"20",x"20",x"20"),
   975 => (x"73",x"20",x"20",x"20"),
   976 => (x"6c",x"75",x"6f",x"68"),
   977 => (x"65",x"62",x"20",x"64"),
   978 => (x"20",x"20",x"20",x"3a"),
   979 => (x"00",x"0a",x"64",x"25"),
   980 => (x"5f",x"72",x"72",x"41"),
   981 => (x"6c",x"47",x"5f",x"32"),
   982 => (x"38",x"5b",x"62",x"6f"),
   983 => (x"5d",x"37",x"5b",x"5d"),
   984 => (x"20",x"20",x"20",x"3a"),
   985 => (x"0a",x"64",x"25",x"20"),
   986 => (x"20",x"20",x"20",x"00"),
   987 => (x"20",x"20",x"20",x"20"),
   988 => (x"6f",x"68",x"73",x"20"),
   989 => (x"20",x"64",x"6c",x"75"),
   990 => (x"20",x"3a",x"65",x"62"),
   991 => (x"75",x"4e",x"20",x"20"),
   992 => (x"72",x"65",x"62",x"6d"),
   993 => (x"5f",x"66",x"4f",x"5f"),
   994 => (x"73",x"6e",x"75",x"52"),
   995 => (x"31",x"20",x"2b",x"20"),
   996 => (x"50",x"00",x"0a",x"30"),
   997 => (x"47",x"5f",x"72",x"74"),
   998 => (x"2d",x"62",x"6f",x"6c"),
   999 => (x"20",x"00",x"0a",x"3e"),
  1000 => (x"72",x"74",x"50",x"20"),
  1001 => (x"6d",x"6f",x"43",x"5f"),
  1002 => (x"20",x"20",x"3a",x"70"),
  1003 => (x"20",x"20",x"20",x"20"),
  1004 => (x"20",x"20",x"20",x"20"),
  1005 => (x"00",x"0a",x"64",x"25"),
  1006 => (x"20",x"20",x"20",x"20"),
  1007 => (x"20",x"20",x"20",x"20"),
  1008 => (x"75",x"6f",x"68",x"73"),
  1009 => (x"62",x"20",x"64",x"6c"),
  1010 => (x"20",x"20",x"3a",x"65"),
  1011 => (x"6d",x"69",x"28",x"20"),
  1012 => (x"6d",x"65",x"6c",x"70"),
  1013 => (x"61",x"74",x"6e",x"65"),
  1014 => (x"6e",x"6f",x"69",x"74"),
  1015 => (x"70",x"65",x"64",x"2d"),
  1016 => (x"65",x"64",x"6e",x"65"),
  1017 => (x"0a",x"29",x"74",x"6e"),
  1018 => (x"44",x"20",x"20",x"00"),
  1019 => (x"72",x"63",x"73",x"69"),
  1020 => (x"20",x"20",x"20",x"3a"),
  1021 => (x"20",x"20",x"20",x"20"),
  1022 => (x"20",x"20",x"20",x"20"),
  1023 => (x"64",x"25",x"20",x"20"),
  1024 => (x"20",x"20",x"00",x"0a"),
  1025 => (x"20",x"20",x"20",x"20"),
  1026 => (x"68",x"73",x"20",x"20"),
  1027 => (x"64",x"6c",x"75",x"6f"),
  1028 => (x"3a",x"65",x"62",x"20"),
  1029 => (x"25",x"20",x"20",x"20"),
  1030 => (x"20",x"00",x"0a",x"64"),
  1031 => (x"75",x"6e",x"45",x"20"),
  1032 => (x"6f",x"43",x"5f",x"6d"),
  1033 => (x"20",x"3a",x"70",x"6d"),
  1034 => (x"20",x"20",x"20",x"20"),
  1035 => (x"20",x"20",x"20",x"20"),
  1036 => (x"00",x"0a",x"64",x"25"),
  1037 => (x"20",x"20",x"20",x"20"),
  1038 => (x"20",x"20",x"20",x"20"),
  1039 => (x"75",x"6f",x"68",x"73"),
  1040 => (x"62",x"20",x"64",x"6c"),
  1041 => (x"20",x"20",x"3a",x"65"),
  1042 => (x"0a",x"64",x"25",x"20"),
  1043 => (x"49",x"20",x"20",x"00"),
  1044 => (x"43",x"5f",x"74",x"6e"),
  1045 => (x"3a",x"70",x"6d",x"6f"),
  1046 => (x"20",x"20",x"20",x"20"),
  1047 => (x"20",x"20",x"20",x"20"),
  1048 => (x"64",x"25",x"20",x"20"),
  1049 => (x"20",x"20",x"00",x"0a"),
  1050 => (x"20",x"20",x"20",x"20"),
  1051 => (x"68",x"73",x"20",x"20"),
  1052 => (x"64",x"6c",x"75",x"6f"),
  1053 => (x"3a",x"65",x"62",x"20"),
  1054 => (x"25",x"20",x"20",x"20"),
  1055 => (x"20",x"00",x"0a",x"64"),
  1056 => (x"72",x"74",x"53",x"20"),
  1057 => (x"6d",x"6f",x"43",x"5f"),
  1058 => (x"20",x"20",x"3a",x"70"),
  1059 => (x"20",x"20",x"20",x"20"),
  1060 => (x"20",x"20",x"20",x"20"),
  1061 => (x"00",x"0a",x"73",x"25"),
  1062 => (x"20",x"20",x"20",x"20"),
  1063 => (x"20",x"20",x"20",x"20"),
  1064 => (x"75",x"6f",x"68",x"73"),
  1065 => (x"62",x"20",x"64",x"6c"),
  1066 => (x"20",x"20",x"3a",x"65"),
  1067 => (x"52",x"48",x"44",x"20"),
  1068 => (x"4f",x"54",x"53",x"59"),
  1069 => (x"50",x"20",x"45",x"4e"),
  1070 => (x"52",x"47",x"4f",x"52"),
  1071 => (x"20",x"2c",x"4d",x"41"),
  1072 => (x"45",x"4d",x"4f",x"53"),
  1073 => (x"52",x"54",x"53",x"20"),
  1074 => (x"0a",x"47",x"4e",x"49"),
  1075 => (x"78",x"65",x"4e",x"00"),
  1076 => (x"74",x"50",x"5f",x"74"),
  1077 => (x"6c",x"47",x"5f",x"72"),
  1078 => (x"3e",x"2d",x"62",x"6f"),
  1079 => (x"20",x"20",x"00",x"0a"),
  1080 => (x"5f",x"72",x"74",x"50"),
  1081 => (x"70",x"6d",x"6f",x"43"),
  1082 => (x"20",x"20",x"20",x"3a"),
  1083 => (x"20",x"20",x"20",x"20"),
  1084 => (x"25",x"20",x"20",x"20"),
  1085 => (x"20",x"00",x"0a",x"64"),
  1086 => (x"20",x"20",x"20",x"20"),
  1087 => (x"73",x"20",x"20",x"20"),
  1088 => (x"6c",x"75",x"6f",x"68"),
  1089 => (x"65",x"62",x"20",x"64"),
  1090 => (x"20",x"20",x"20",x"3a"),
  1091 => (x"70",x"6d",x"69",x"28"),
  1092 => (x"65",x"6d",x"65",x"6c"),
  1093 => (x"74",x"61",x"74",x"6e"),
  1094 => (x"2d",x"6e",x"6f",x"69"),
  1095 => (x"65",x"70",x"65",x"64"),
  1096 => (x"6e",x"65",x"64",x"6e"),
  1097 => (x"20",x"2c",x"29",x"74"),
  1098 => (x"65",x"6d",x"61",x"73"),
  1099 => (x"20",x"73",x"61",x"20"),
  1100 => (x"76",x"6f",x"62",x"61"),
  1101 => (x"20",x"00",x"0a",x"65"),
  1102 => (x"73",x"69",x"44",x"20"),
  1103 => (x"20",x"3a",x"72",x"63"),
  1104 => (x"20",x"20",x"20",x"20"),
  1105 => (x"20",x"20",x"20",x"20"),
  1106 => (x"20",x"20",x"20",x"20"),
  1107 => (x"00",x"0a",x"64",x"25"),
  1108 => (x"20",x"20",x"20",x"20"),
  1109 => (x"20",x"20",x"20",x"20"),
  1110 => (x"75",x"6f",x"68",x"73"),
  1111 => (x"62",x"20",x"64",x"6c"),
  1112 => (x"20",x"20",x"3a",x"65"),
  1113 => (x"0a",x"64",x"25",x"20"),
  1114 => (x"45",x"20",x"20",x"00"),
  1115 => (x"5f",x"6d",x"75",x"6e"),
  1116 => (x"70",x"6d",x"6f",x"43"),
  1117 => (x"20",x"20",x"20",x"3a"),
  1118 => (x"20",x"20",x"20",x"20"),
  1119 => (x"64",x"25",x"20",x"20"),
  1120 => (x"20",x"20",x"00",x"0a"),
  1121 => (x"20",x"20",x"20",x"20"),
  1122 => (x"68",x"73",x"20",x"20"),
  1123 => (x"64",x"6c",x"75",x"6f"),
  1124 => (x"3a",x"65",x"62",x"20"),
  1125 => (x"25",x"20",x"20",x"20"),
  1126 => (x"20",x"00",x"0a",x"64"),
  1127 => (x"74",x"6e",x"49",x"20"),
  1128 => (x"6d",x"6f",x"43",x"5f"),
  1129 => (x"20",x"20",x"3a",x"70"),
  1130 => (x"20",x"20",x"20",x"20"),
  1131 => (x"20",x"20",x"20",x"20"),
  1132 => (x"00",x"0a",x"64",x"25"),
  1133 => (x"20",x"20",x"20",x"20"),
  1134 => (x"20",x"20",x"20",x"20"),
  1135 => (x"75",x"6f",x"68",x"73"),
  1136 => (x"62",x"20",x"64",x"6c"),
  1137 => (x"20",x"20",x"3a",x"65"),
  1138 => (x"0a",x"64",x"25",x"20"),
  1139 => (x"53",x"20",x"20",x"00"),
  1140 => (x"43",x"5f",x"72",x"74"),
  1141 => (x"3a",x"70",x"6d",x"6f"),
  1142 => (x"20",x"20",x"20",x"20"),
  1143 => (x"20",x"20",x"20",x"20"),
  1144 => (x"73",x"25",x"20",x"20"),
  1145 => (x"20",x"20",x"00",x"0a"),
  1146 => (x"20",x"20",x"20",x"20"),
  1147 => (x"68",x"73",x"20",x"20"),
  1148 => (x"64",x"6c",x"75",x"6f"),
  1149 => (x"3a",x"65",x"62",x"20"),
  1150 => (x"44",x"20",x"20",x"20"),
  1151 => (x"53",x"59",x"52",x"48"),
  1152 => (x"45",x"4e",x"4f",x"54"),
  1153 => (x"4f",x"52",x"50",x"20"),
  1154 => (x"4d",x"41",x"52",x"47"),
  1155 => (x"4f",x"53",x"20",x"2c"),
  1156 => (x"53",x"20",x"45",x"4d"),
  1157 => (x"4e",x"49",x"52",x"54"),
  1158 => (x"49",x"00",x"0a",x"47"),
  1159 => (x"31",x"5f",x"74",x"6e"),
  1160 => (x"63",x"6f",x"4c",x"5f"),
  1161 => (x"20",x"20",x"20",x"3a"),
  1162 => (x"20",x"20",x"20",x"20"),
  1163 => (x"20",x"20",x"20",x"20"),
  1164 => (x"00",x"0a",x"64",x"25"),
  1165 => (x"20",x"20",x"20",x"20"),
  1166 => (x"20",x"20",x"20",x"20"),
  1167 => (x"75",x"6f",x"68",x"73"),
  1168 => (x"62",x"20",x"64",x"6c"),
  1169 => (x"20",x"20",x"3a",x"65"),
  1170 => (x"0a",x"64",x"25",x"20"),
  1171 => (x"74",x"6e",x"49",x"00"),
  1172 => (x"4c",x"5f",x"32",x"5f"),
  1173 => (x"20",x"3a",x"63",x"6f"),
  1174 => (x"20",x"20",x"20",x"20"),
  1175 => (x"20",x"20",x"20",x"20"),
  1176 => (x"64",x"25",x"20",x"20"),
  1177 => (x"20",x"20",x"00",x"0a"),
  1178 => (x"20",x"20",x"20",x"20"),
  1179 => (x"68",x"73",x"20",x"20"),
  1180 => (x"64",x"6c",x"75",x"6f"),
  1181 => (x"3a",x"65",x"62",x"20"),
  1182 => (x"25",x"20",x"20",x"20"),
  1183 => (x"49",x"00",x"0a",x"64"),
  1184 => (x"33",x"5f",x"74",x"6e"),
  1185 => (x"63",x"6f",x"4c",x"5f"),
  1186 => (x"20",x"20",x"20",x"3a"),
  1187 => (x"20",x"20",x"20",x"20"),
  1188 => (x"20",x"20",x"20",x"20"),
  1189 => (x"00",x"0a",x"64",x"25"),
  1190 => (x"20",x"20",x"20",x"20"),
  1191 => (x"20",x"20",x"20",x"20"),
  1192 => (x"75",x"6f",x"68",x"73"),
  1193 => (x"62",x"20",x"64",x"6c"),
  1194 => (x"20",x"20",x"3a",x"65"),
  1195 => (x"0a",x"64",x"25",x"20"),
  1196 => (x"75",x"6e",x"45",x"00"),
  1197 => (x"6f",x"4c",x"5f",x"6d"),
  1198 => (x"20",x"20",x"3a",x"63"),
  1199 => (x"20",x"20",x"20",x"20"),
  1200 => (x"20",x"20",x"20",x"20"),
  1201 => (x"64",x"25",x"20",x"20"),
  1202 => (x"20",x"20",x"00",x"0a"),
  1203 => (x"20",x"20",x"20",x"20"),
  1204 => (x"68",x"73",x"20",x"20"),
  1205 => (x"64",x"6c",x"75",x"6f"),
  1206 => (x"3a",x"65",x"62",x"20"),
  1207 => (x"25",x"20",x"20",x"20"),
  1208 => (x"53",x"00",x"0a",x"64"),
  1209 => (x"31",x"5f",x"72",x"74"),
  1210 => (x"63",x"6f",x"4c",x"5f"),
  1211 => (x"20",x"20",x"20",x"3a"),
  1212 => (x"20",x"20",x"20",x"20"),
  1213 => (x"20",x"20",x"20",x"20"),
  1214 => (x"00",x"0a",x"73",x"25"),
  1215 => (x"20",x"20",x"20",x"20"),
  1216 => (x"20",x"20",x"20",x"20"),
  1217 => (x"75",x"6f",x"68",x"73"),
  1218 => (x"62",x"20",x"64",x"6c"),
  1219 => (x"20",x"20",x"3a",x"65"),
  1220 => (x"52",x"48",x"44",x"20"),
  1221 => (x"4f",x"54",x"53",x"59"),
  1222 => (x"50",x"20",x"45",x"4e"),
  1223 => (x"52",x"47",x"4f",x"52"),
  1224 => (x"20",x"2c",x"4d",x"41"),
  1225 => (x"54",x"53",x"27",x"31"),
  1226 => (x"52",x"54",x"53",x"20"),
  1227 => (x"0a",x"47",x"4e",x"49"),
  1228 => (x"72",x"74",x"53",x"00"),
  1229 => (x"4c",x"5f",x"32",x"5f"),
  1230 => (x"20",x"3a",x"63",x"6f"),
  1231 => (x"20",x"20",x"20",x"20"),
  1232 => (x"20",x"20",x"20",x"20"),
  1233 => (x"73",x"25",x"20",x"20"),
  1234 => (x"20",x"20",x"00",x"0a"),
  1235 => (x"20",x"20",x"20",x"20"),
  1236 => (x"68",x"73",x"20",x"20"),
  1237 => (x"64",x"6c",x"75",x"6f"),
  1238 => (x"3a",x"65",x"62",x"20"),
  1239 => (x"44",x"20",x"20",x"20"),
  1240 => (x"53",x"59",x"52",x"48"),
  1241 => (x"45",x"4e",x"4f",x"54"),
  1242 => (x"4f",x"52",x"50",x"20"),
  1243 => (x"4d",x"41",x"52",x"47"),
  1244 => (x"27",x"32",x"20",x"2c"),
  1245 => (x"53",x"20",x"44",x"4e"),
  1246 => (x"4e",x"49",x"52",x"54"),
  1247 => (x"0a",x"00",x"0a",x"47"),
  1248 => (x"65",x"73",x"55",x"00"),
  1249 => (x"69",x"74",x"20",x"72"),
  1250 => (x"20",x"3a",x"65",x"6d"),
  1251 => (x"00",x"0a",x"64",x"25"),
  1252 => (x"0e",x"5b",x"5e",x"0e"),
  1253 => (x"cc",x"4b",x"66",x"c8"),
  1254 => (x"79",x"73",x"49",x"66"),
  1255 => (x"c4",x"05",x"ab",x"c2"),
  1256 => (x"c2",x"4a",x"c1",x"87"),
  1257 => (x"72",x"4a",x"c0",x"87"),
  1258 => (x"87",x"c2",x"05",x"9a"),
  1259 => (x"ab",x"c0",x"79",x"c3"),
  1260 => (x"c1",x"87",x"d8",x"02"),
  1261 => (x"87",x"d7",x"02",x"ab"),
  1262 => (x"c0",x"02",x"ab",x"c2"),
  1263 => (x"ab",x"c3",x"87",x"e5"),
  1264 => (x"87",x"e5",x"c0",x"02"),
  1265 => (x"de",x"02",x"ab",x"c4"),
  1266 => (x"c0",x"87",x"de",x"87"),
  1267 => (x"c1",x"87",x"da",x"79"),
  1268 => (x"48",x"bf",x"c2",x"d6"),
  1269 => (x"a8",x"b7",x"e4",x"c1"),
  1270 => (x"c0",x"87",x"c4",x"06"),
  1271 => (x"c3",x"87",x"ca",x"79"),
  1272 => (x"c1",x"87",x"c6",x"79"),
  1273 => (x"c2",x"87",x"c2",x"79"),
  1274 => (x"26",x"4b",x"26",x"79"),
  1275 => (x"66",x"c4",x"1e",x"4f"),
  1276 => (x"05",x"a8",x"c2",x"48"),
  1277 => (x"48",x"c1",x"87",x"c4"),
  1278 => (x"48",x"c0",x"87",x"c2"),
  1279 => (x"c4",x"1e",x"4f",x"26"),
  1280 => (x"81",x"c2",x"49",x"66"),
  1281 => (x"71",x"48",x"66",x"c8"),
  1282 => (x"08",x"66",x"cc",x"80"),
  1283 => (x"4f",x"26",x"08",x"78"),
  1284 => (x"5c",x"5b",x"5e",x"0e"),
  1285 => (x"86",x"f4",x"0e",x"5d"),
  1286 => (x"4c",x"66",x"e4",x"c0"),
  1287 => (x"48",x"74",x"84",x"c5"),
  1288 => (x"c8",x"90",x"b7",x"c4"),
  1289 => (x"66",x"dc",x"58",x"a6"),
  1290 => (x"80",x"66",x"c4",x"48"),
  1291 => (x"6e",x"58",x"a6",x"c4"),
  1292 => (x"66",x"e8",x"c0",x"48"),
  1293 => (x"c1",x"48",x"74",x"78"),
  1294 => (x"58",x"a6",x"cc",x"80"),
  1295 => (x"c4",x"49",x"66",x"c8"),
  1296 => (x"66",x"dc",x"91",x"b7"),
  1297 => (x"66",x"e8",x"c0",x"81"),
  1298 => (x"de",x"49",x"74",x"79"),
  1299 => (x"91",x"b7",x"c4",x"81"),
  1300 => (x"74",x"81",x"66",x"dc"),
  1301 => (x"b7",x"66",x"c8",x"79"),
  1302 => (x"e3",x"c0",x"01",x"ac"),
  1303 => (x"c3",x"49",x"74",x"87"),
  1304 => (x"c0",x"91",x"b7",x"c8"),
  1305 => (x"c4",x"81",x"66",x"e0"),
  1306 => (x"c4",x"4a",x"71",x"4d"),
  1307 => (x"66",x"c8",x"82",x"66"),
  1308 => (x"c1",x"8b",x"74",x"4b"),
  1309 => (x"75",x"7a",x"74",x"83"),
  1310 => (x"73",x"8b",x"c1",x"82"),
  1311 => (x"87",x"f5",x"01",x"9b"),
  1312 => (x"c8",x"c3",x"4a",x"74"),
  1313 => (x"e0",x"c0",x"92",x"b7"),
  1314 => (x"49",x"74",x"82",x"66"),
  1315 => (x"b7",x"c4",x"89",x"c1"),
  1316 => (x"69",x"81",x"72",x"91"),
  1317 => (x"70",x"80",x"c1",x"48"),
  1318 => (x"d4",x"49",x"74",x"79"),
  1319 => (x"b7",x"c8",x"c3",x"81"),
  1320 => (x"66",x"e0",x"c0",x"91"),
  1321 => (x"81",x"66",x"c4",x"81"),
  1322 => (x"c1",x"79",x"bf",x"6e"),
  1323 => (x"c5",x"48",x"c2",x"d6"),
  1324 => (x"26",x"8e",x"f4",x"78"),
  1325 => (x"26",x"4c",x"26",x"4d"),
  1326 => (x"0e",x"4f",x"26",x"4b"),
  1327 => (x"97",x"0e",x"5b",x"5e"),
  1328 => (x"73",x"4b",x"66",x"c8"),
  1329 => (x"82",x"c0",x"fe",x"4a"),
  1330 => (x"66",x"cc",x"97",x"ba"),
  1331 => (x"81",x"c0",x"fe",x"49"),
  1332 => (x"aa",x"b7",x"71",x"b9"),
  1333 => (x"c0",x"87",x"c4",x"02"),
  1334 => (x"c1",x"87",x"c7",x"48"),
  1335 => (x"5b",x"97",x"ce",x"d6"),
  1336 => (x"4b",x"26",x"48",x"c1"),
  1337 => (x"5e",x"0e",x"4f",x"26"),
  1338 => (x"0e",x"5d",x"5c",x"5b"),
  1339 => (x"4d",x"c2",x"86",x"f8"),
  1340 => (x"c1",x"49",x"66",x"dc"),
  1341 => (x"4c",x"66",x"d8",x"81"),
  1342 => (x"4b",x"71",x"84",x"c2"),
  1343 => (x"49",x"13",x"83",x"c2"),
  1344 => (x"b9",x"81",x"c0",x"fe"),
  1345 => (x"14",x"99",x"ff",x"c3"),
  1346 => (x"82",x"c0",x"fe",x"4a"),
  1347 => (x"97",x"a6",x"c4",x"ba"),
  1348 => (x"4a",x"6e",x"97",x"5a"),
  1349 => (x"ba",x"82",x"c0",x"fe"),
  1350 => (x"b9",x"81",x"c0",x"fe"),
  1351 => (x"02",x"aa",x"b7",x"71"),
  1352 => (x"a6",x"c4",x"87",x"c7"),
  1353 => (x"cc",x"78",x"c0",x"48"),
  1354 => (x"ca",x"d6",x"c1",x"87"),
  1355 => (x"50",x"6e",x"97",x"48"),
  1356 => (x"c1",x"48",x"a6",x"c4"),
  1357 => (x"05",x"66",x"c4",x"78"),
  1358 => (x"85",x"c1",x"87",x"c2"),
  1359 => (x"06",x"ad",x"b7",x"c2"),
  1360 => (x"d8",x"87",x"fb",x"fe"),
  1361 => (x"66",x"dc",x"4a",x"66"),
  1362 => (x"0f",x"ec",x"cf",x"49"),
  1363 => (x"06",x"a8",x"b7",x"c0"),
  1364 => (x"48",x"75",x"87",x"cc"),
  1365 => (x"d6",x"c1",x"80",x"c7"),
  1366 => (x"48",x"c1",x"58",x"c6"),
  1367 => (x"48",x"c0",x"87",x"c2"),
  1368 => (x"4d",x"26",x"8e",x"f8"),
  1369 => (x"4b",x"26",x"4c",x"26"),
  1370 => (x"4b",x"26",x"4f",x"26"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
