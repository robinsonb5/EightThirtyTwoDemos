
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"d7",x"01"),
     1 => (x"58",x"0e",x"87",x"da"),
     2 => (x"27",x"0e",x"59",x"5e"),
     3 => (x"00",x"00",x"00",x"41"),
     4 => (x"26",x"49",x"26",x"0f"),
     5 => (x"26",x"80",x"ff",x"48"),
     6 => (x"26",x"27",x"4f",x"08"),
     7 => (x"4f",x"00",x"00",x"00"),
     8 => (x"00",x"00",x"33",x"27"),
     9 => (x"c0",x"c2",x"4f",x"00"),
    10 => (x"6b",x"27",x"4e",x"c0"),
    11 => (x"0f",x"00",x"00",x"16"),
    12 => (x"c1",x"87",x"fd",x"00"),
    13 => (x"27",x"4e",x"c0",x"f0"),
    14 => (x"00",x"00",x"00",x"40"),
    15 => (x"87",x"fd",x"00",x"0f"),
    16 => (x"72",x"1e",x"4f",x"4f"),
    17 => (x"c0",x"ff",x"1e",x"1e"),
    18 => (x"c4",x"48",x"6a",x"4a"),
    19 => (x"a6",x"c4",x"98",x"c0"),
    20 => (x"ff",x"02",x"6e",x"58"),
    21 => (x"66",x"cc",x"87",x"f3"),
    22 => (x"48",x"66",x"cc",x"7a"),
    23 => (x"26",x"4a",x"26",x"26"),
    24 => (x"5a",x"5e",x"0e",x"4f"),
    25 => (x"0e",x"5d",x"5c",x"5b"),
    26 => (x"c0",x"4b",x"66",x"d4"),
    27 => (x"74",x"4c",x"13",x"4d"),
    28 => (x"d9",x"c0",x"02",x"9c"),
    29 => (x"c3",x"4a",x"74",x"87"),
    30 => (x"1e",x"72",x"9a",x"ff"),
    31 => (x"00",x"00",x"42",x"27"),
    32 => (x"86",x"c4",x"0f",x"00"),
    33 => (x"4c",x"13",x"85",x"c1"),
    34 => (x"ff",x"05",x"9c",x"74"),
    35 => (x"48",x"75",x"87",x"e7"),
    36 => (x"4c",x"26",x"4d",x"26"),
    37 => (x"4a",x"26",x"4b",x"26"),
    38 => (x"5e",x"0e",x"4f",x"26"),
    39 => (x"5d",x"5c",x"5b",x"5a"),
    40 => (x"c0",x"8e",x"d0",x"0e"),
    41 => (x"49",x"a6",x"c4",x"4c"),
    42 => (x"e8",x"c0",x"79",x"c0"),
    43 => (x"e4",x"c0",x"4b",x"a6"),
    44 => (x"e4",x"c0",x"4a",x"66"),
    45 => (x"80",x"c1",x"48",x"66"),
    46 => (x"58",x"a6",x"e8",x"c0"),
    47 => (x"c0",x"c1",x"48",x"12"),
    48 => (x"90",x"c0",x"c0",x"c0"),
    49 => (x"90",x"b7",x"c0",x"c4"),
    50 => (x"58",x"a6",x"c4",x"48"),
    51 => (x"c2",x"c5",x"02",x"6e"),
    52 => (x"02",x"66",x"c4",x"87"),
    53 => (x"c4",x"87",x"fe",x"c3"),
    54 => (x"79",x"c0",x"49",x"a6"),
    55 => (x"49",x"6e",x"4a",x"6e"),
    56 => (x"02",x"a9",x"f0",x"c0"),
    57 => (x"c1",x"87",x"c4",x"c3"),
    58 => (x"c3",x"02",x"aa",x"e3"),
    59 => (x"e4",x"c1",x"87",x"c5"),
    60 => (x"e3",x"c0",x"02",x"aa"),
    61 => (x"aa",x"ec",x"c1",x"87"),
    62 => (x"87",x"ef",x"c2",x"02"),
    63 => (x"02",x"aa",x"f0",x"c1"),
    64 => (x"c1",x"87",x"d5",x"c0"),
    65 => (x"c2",x"02",x"aa",x"f3"),
    66 => (x"f5",x"c1",x"87",x"c8"),
    67 => (x"c7",x"c0",x"02",x"aa"),
    68 => (x"aa",x"f8",x"c1",x"87"),
    69 => (x"87",x"f0",x"c2",x"05"),
    70 => (x"4a",x"73",x"83",x"c4"),
    71 => (x"49",x"76",x"8a",x"c4"),
    72 => (x"02",x"6e",x"79",x"6a"),
    73 => (x"c8",x"87",x"db",x"c1"),
    74 => (x"79",x"c0",x"49",x"a6"),
    75 => (x"c0",x"49",x"a6",x"cc"),
    76 => (x"dc",x"4a",x"6e",x"79"),
    77 => (x"4d",x"72",x"2a",x"b7"),
    78 => (x"48",x"6e",x"9d",x"cf"),
    79 => (x"a6",x"c4",x"30",x"c4"),
    80 => (x"02",x"9d",x"75",x"58"),
    81 => (x"c8",x"87",x"c5",x"c0"),
    82 => (x"79",x"c1",x"49",x"a6"),
    83 => (x"c0",x"06",x"ad",x"c9"),
    84 => (x"f7",x"c0",x"87",x"c6"),
    85 => (x"87",x"c3",x"c0",x"85"),
    86 => (x"c8",x"85",x"f0",x"c0"),
    87 => (x"cc",x"c0",x"02",x"66"),
    88 => (x"27",x"1e",x"75",x"87"),
    89 => (x"00",x"00",x"00",x"42"),
    90 => (x"c1",x"86",x"c4",x"0f"),
    91 => (x"48",x"66",x"cc",x"84"),
    92 => (x"a6",x"d0",x"80",x"c1"),
    93 => (x"49",x"66",x"cc",x"58"),
    94 => (x"04",x"a9",x"b7",x"c8"),
    95 => (x"c1",x"87",x"f2",x"fe"),
    96 => (x"f0",x"c0",x"87",x"ee"),
    97 => (x"00",x"42",x"27",x"1e"),
    98 => (x"c4",x"0f",x"00",x"00"),
    99 => (x"c1",x"84",x"c1",x"86"),
   100 => (x"83",x"c4",x"87",x"de"),
   101 => (x"8a",x"c4",x"4a",x"73"),
   102 => (x"61",x"27",x"1e",x"6a"),
   103 => (x"0f",x"00",x"00",x"00"),
   104 => (x"4a",x"70",x"86",x"c4"),
   105 => (x"84",x"72",x"4c",x"74"),
   106 => (x"c4",x"87",x"c5",x"c1"),
   107 => (x"79",x"c1",x"49",x"a6"),
   108 => (x"c4",x"87",x"fd",x"c0"),
   109 => (x"c4",x"4a",x"73",x"83"),
   110 => (x"27",x"1e",x"6a",x"8a"),
   111 => (x"00",x"00",x"00",x"42"),
   112 => (x"c1",x"86",x"c4",x"0f"),
   113 => (x"87",x"e8",x"c0",x"84"),
   114 => (x"42",x"27",x"1e",x"6e"),
   115 => (x"0f",x"00",x"00",x"00"),
   116 => (x"db",x"c0",x"86",x"c4"),
   117 => (x"c0",x"49",x"6e",x"87"),
   118 => (x"c0",x"05",x"a9",x"e5"),
   119 => (x"a6",x"c4",x"87",x"c8"),
   120 => (x"c0",x"79",x"c1",x"49"),
   121 => (x"1e",x"6e",x"87",x"ca"),
   122 => (x"00",x"00",x"42",x"27"),
   123 => (x"86",x"c4",x"0f",x"00"),
   124 => (x"4a",x"66",x"e4",x"c0"),
   125 => (x"48",x"66",x"e4",x"c0"),
   126 => (x"e8",x"c0",x"80",x"c1"),
   127 => (x"48",x"12",x"58",x"a6"),
   128 => (x"c0",x"c0",x"c0",x"c1"),
   129 => (x"c0",x"c4",x"90",x"c0"),
   130 => (x"c4",x"48",x"90",x"b7"),
   131 => (x"05",x"6e",x"58",x"a6"),
   132 => (x"74",x"87",x"fe",x"fa"),
   133 => (x"26",x"86",x"d0",x"48"),
   134 => (x"26",x"4c",x"26",x"4d"),
   135 => (x"26",x"4a",x"26",x"4b"),
   136 => (x"00",x"00",x"00",x"4f"),
   137 => (x"1e",x"75",x"1e",x"00"),
   138 => (x"c3",x"4d",x"d4",x"ff"),
   139 => (x"6d",x"7d",x"49",x"ff"),
   140 => (x"71",x"38",x"c8",x"48"),
   141 => (x"c8",x"b0",x"6d",x"7d"),
   142 => (x"6d",x"7d",x"71",x"38"),
   143 => (x"71",x"38",x"c8",x"b0"),
   144 => (x"c8",x"b0",x"6d",x"7d"),
   145 => (x"26",x"4d",x"26",x"38"),
   146 => (x"1e",x"75",x"1e",x"4f"),
   147 => (x"c3",x"4d",x"d4",x"ff"),
   148 => (x"6d",x"7d",x"49",x"ff"),
   149 => (x"71",x"30",x"c8",x"48"),
   150 => (x"c8",x"b0",x"6d",x"7d"),
   151 => (x"6d",x"7d",x"71",x"30"),
   152 => (x"71",x"30",x"c8",x"b0"),
   153 => (x"26",x"b0",x"6d",x"7d"),
   154 => (x"1e",x"4f",x"26",x"4d"),
   155 => (x"d4",x"ff",x"1e",x"75"),
   156 => (x"49",x"66",x"cc",x"4d"),
   157 => (x"7d",x"48",x"66",x"c8"),
   158 => (x"02",x"67",x"e6",x"fe"),
   159 => (x"d8",x"07",x"31",x"c9"),
   160 => (x"09",x"7d",x"09",x"39"),
   161 => (x"09",x"7d",x"09",x"39"),
   162 => (x"09",x"7d",x"09",x"39"),
   163 => (x"d0",x"7d",x"09",x"39"),
   164 => (x"c9",x"7d",x"70",x"38"),
   165 => (x"c3",x"49",x"c0",x"f1"),
   166 => (x"08",x"6d",x"48",x"ff"),
   167 => (x"87",x"c7",x"05",x"a8"),
   168 => (x"89",x"c1",x"7d",x"08"),
   169 => (x"26",x"87",x"f3",x"05"),
   170 => (x"1e",x"4f",x"26",x"4d"),
   171 => (x"c3",x"49",x"d4",x"ff"),
   172 => (x"79",x"ff",x"48",x"c8"),
   173 => (x"87",x"fa",x"05",x"80"),
   174 => (x"5e",x"0e",x"4f",x"26"),
   175 => (x"5d",x"5c",x"5b",x"5a"),
   176 => (x"f0",x"ff",x"c0",x"0e"),
   177 => (x"c1",x"4d",x"f7",x"c1"),
   178 => (x"c0",x"c0",x"c0",x"c0"),
   179 => (x"ab",x"27",x"4b",x"c0"),
   180 => (x"0f",x"00",x"00",x"02"),
   181 => (x"4c",x"df",x"f8",x"c4"),
   182 => (x"1e",x"75",x"1e",x"c0"),
   183 => (x"00",x"02",x"6b",x"27"),
   184 => (x"86",x"c8",x"0f",x"00"),
   185 => (x"b7",x"c1",x"4a",x"70"),
   186 => (x"ef",x"c0",x"05",x"aa"),
   187 => (x"49",x"d4",x"ff",x"87"),
   188 => (x"73",x"79",x"ff",x"c3"),
   189 => (x"f0",x"e1",x"c0",x"1e"),
   190 => (x"27",x"1e",x"e9",x"c1"),
   191 => (x"00",x"00",x"02",x"6b"),
   192 => (x"70",x"86",x"c8",x"0f"),
   193 => (x"05",x"9a",x"72",x"4a"),
   194 => (x"ff",x"87",x"cb",x"c0"),
   195 => (x"ff",x"c3",x"49",x"d4"),
   196 => (x"c0",x"48",x"c1",x"79"),
   197 => (x"ab",x"27",x"87",x"d0"),
   198 => (x"0f",x"00",x"00",x"02"),
   199 => (x"9c",x"74",x"8c",x"c1"),
   200 => (x"87",x"f4",x"fe",x"05"),
   201 => (x"4d",x"26",x"48",x"c0"),
   202 => (x"4b",x"26",x"4c",x"26"),
   203 => (x"4f",x"26",x"4a",x"26"),
   204 => (x"5b",x"5a",x"5e",x"0e"),
   205 => (x"ff",x"c0",x"0e",x"5c"),
   206 => (x"4c",x"c1",x"c1",x"f0"),
   207 => (x"c3",x"49",x"d4",x"ff"),
   208 => (x"bc",x"27",x"79",x"ff"),
   209 => (x"1e",x"00",x"00",x"17"),
   210 => (x"00",x"00",x"61",x"27"),
   211 => (x"86",x"c4",x"0f",x"00"),
   212 => (x"1e",x"c0",x"4b",x"d3"),
   213 => (x"6b",x"27",x"1e",x"74"),
   214 => (x"0f",x"00",x"00",x"02"),
   215 => (x"4a",x"70",x"86",x"c8"),
   216 => (x"c0",x"05",x"9a",x"72"),
   217 => (x"d4",x"ff",x"87",x"cb"),
   218 => (x"79",x"ff",x"c3",x"49"),
   219 => (x"d0",x"c0",x"48",x"c1"),
   220 => (x"02",x"ab",x"27",x"87"),
   221 => (x"c1",x"0f",x"00",x"00"),
   222 => (x"05",x"9b",x"73",x"8b"),
   223 => (x"c0",x"87",x"d3",x"ff"),
   224 => (x"26",x"4c",x"26",x"48"),
   225 => (x"26",x"4a",x"26",x"4b"),
   226 => (x"5a",x"5e",x"0e",x"4f"),
   227 => (x"0e",x"5d",x"5c",x"5b"),
   228 => (x"4d",x"ff",x"c3",x"1e"),
   229 => (x"27",x"4c",x"d4",x"ff"),
   230 => (x"00",x"00",x"02",x"ab"),
   231 => (x"1e",x"ea",x"c6",x"0f"),
   232 => (x"c1",x"f0",x"e1",x"c0"),
   233 => (x"6b",x"27",x"1e",x"c8"),
   234 => (x"0f",x"00",x"00",x"02"),
   235 => (x"4a",x"70",x"86",x"c8"),
   236 => (x"e8",x"27",x"1e",x"72"),
   237 => (x"1e",x"00",x"00",x"04"),
   238 => (x"00",x"00",x"9a",x"27"),
   239 => (x"86",x"c8",x"0f",x"00"),
   240 => (x"02",x"aa",x"b7",x"c1"),
   241 => (x"27",x"87",x"cb",x"c0"),
   242 => (x"00",x"00",x"03",x"30"),
   243 => (x"c3",x"48",x"c0",x"0f"),
   244 => (x"49",x"27",x"87",x"c9"),
   245 => (x"0f",x"00",x"00",x"02"),
   246 => (x"ff",x"cf",x"4a",x"70"),
   247 => (x"ea",x"c6",x"9a",x"ff"),
   248 => (x"c0",x"02",x"aa",x"b7"),
   249 => (x"30",x"27",x"87",x"cb"),
   250 => (x"0f",x"00",x"00",x"03"),
   251 => (x"ea",x"c2",x"48",x"c0"),
   252 => (x"76",x"7c",x"75",x"87"),
   253 => (x"79",x"f1",x"c0",x"49"),
   254 => (x"00",x"02",x"ba",x"27"),
   255 => (x"4a",x"70",x"0f",x"00"),
   256 => (x"c1",x"02",x"9a",x"72"),
   257 => (x"1e",x"c0",x"87",x"eb"),
   258 => (x"c1",x"f0",x"ff",x"c0"),
   259 => (x"6b",x"27",x"1e",x"fa"),
   260 => (x"0f",x"00",x"00",x"02"),
   261 => (x"4b",x"70",x"86",x"c8"),
   262 => (x"c1",x"05",x"9b",x"73"),
   263 => (x"1e",x"73",x"87",x"c3"),
   264 => (x"00",x"04",x"a6",x"27"),
   265 => (x"9a",x"27",x"1e",x"00"),
   266 => (x"0f",x"00",x"00",x"00"),
   267 => (x"7c",x"75",x"86",x"c8"),
   268 => (x"9b",x"75",x"4b",x"6c"),
   269 => (x"b2",x"27",x"1e",x"73"),
   270 => (x"1e",x"00",x"00",x"04"),
   271 => (x"00",x"00",x"9a",x"27"),
   272 => (x"86",x"c8",x"0f",x"00"),
   273 => (x"7c",x"75",x"7c",x"75"),
   274 => (x"7c",x"75",x"7c",x"75"),
   275 => (x"c0",x"c1",x"4a",x"73"),
   276 => (x"02",x"9a",x"72",x"9a"),
   277 => (x"c1",x"87",x"c5",x"c0"),
   278 => (x"87",x"ff",x"c0",x"48"),
   279 => (x"fa",x"c0",x"48",x"c0"),
   280 => (x"27",x"1e",x"73",x"87"),
   281 => (x"00",x"00",x"04",x"c0"),
   282 => (x"00",x"9a",x"27",x"1e"),
   283 => (x"c8",x"0f",x"00",x"00"),
   284 => (x"c2",x"49",x"6e",x"86"),
   285 => (x"c0",x"05",x"a9",x"b7"),
   286 => (x"cc",x"27",x"87",x"d3"),
   287 => (x"1e",x"00",x"00",x"04"),
   288 => (x"00",x"00",x"9a",x"27"),
   289 => (x"86",x"c4",x"0f",x"00"),
   290 => (x"ce",x"c0",x"48",x"c0"),
   291 => (x"c1",x"48",x"6e",x"87"),
   292 => (x"58",x"a6",x"c4",x"88"),
   293 => (x"df",x"fd",x"05",x"6e"),
   294 => (x"26",x"48",x"c0",x"87"),
   295 => (x"4c",x"26",x"4d",x"26"),
   296 => (x"4a",x"26",x"4b",x"26"),
   297 => (x"4d",x"43",x"4f",x"26"),
   298 => (x"20",x"38",x"35",x"44"),
   299 => (x"20",x"0a",x"64",x"25"),
   300 => (x"4d",x"43",x"00",x"20"),
   301 => (x"5f",x"38",x"35",x"44"),
   302 => (x"64",x"25",x"20",x"32"),
   303 => (x"00",x"20",x"20",x"0a"),
   304 => (x"35",x"44",x"4d",x"43"),
   305 => (x"64",x"25",x"20",x"38"),
   306 => (x"00",x"20",x"20",x"0a"),
   307 => (x"43",x"48",x"44",x"53"),
   308 => (x"69",x"6e",x"49",x"20"),
   309 => (x"6c",x"61",x"69",x"74"),
   310 => (x"74",x"61",x"7a",x"69"),
   311 => (x"20",x"6e",x"6f",x"69"),
   312 => (x"6f",x"72",x"72",x"65"),
   313 => (x"00",x"0a",x"21",x"72"),
   314 => (x"5f",x"64",x"6d",x"63"),
   315 => (x"38",x"44",x"4d",x"43"),
   316 => (x"73",x"65",x"72",x"20"),
   317 => (x"73",x"6e",x"6f",x"70"),
   318 => (x"25",x"20",x"3a",x"65"),
   319 => (x"0e",x"00",x"0a",x"64"),
   320 => (x"5c",x"5b",x"5a",x"5e"),
   321 => (x"ff",x"1e",x"0e",x"5d"),
   322 => (x"c0",x"c8",x"4c",x"d0"),
   323 => (x"21",x"27",x"4b",x"c0"),
   324 => (x"49",x"00",x"00",x"02"),
   325 => (x"1c",x"27",x"79",x"c1"),
   326 => (x"1e",x"00",x"00",x"06"),
   327 => (x"00",x"00",x"61",x"27"),
   328 => (x"86",x"c4",x"0f",x"00"),
   329 => (x"48",x"6c",x"4d",x"c7"),
   330 => (x"a6",x"c4",x"98",x"73"),
   331 => (x"c0",x"02",x"6e",x"58"),
   332 => (x"48",x"6c",x"87",x"cc"),
   333 => (x"a6",x"c4",x"98",x"73"),
   334 => (x"ff",x"05",x"6e",x"58"),
   335 => (x"7c",x"c0",x"87",x"f4"),
   336 => (x"00",x"02",x"ab",x"27"),
   337 => (x"48",x"6c",x"0f",x"00"),
   338 => (x"a6",x"c4",x"98",x"73"),
   339 => (x"c0",x"02",x"6e",x"58"),
   340 => (x"48",x"6c",x"87",x"cc"),
   341 => (x"a6",x"c4",x"98",x"73"),
   342 => (x"ff",x"05",x"6e",x"58"),
   343 => (x"7c",x"c1",x"87",x"f4"),
   344 => (x"e5",x"c0",x"1e",x"c0"),
   345 => (x"1e",x"c0",x"c1",x"d0"),
   346 => (x"00",x"02",x"6b",x"27"),
   347 => (x"86",x"c8",x"0f",x"00"),
   348 => (x"b7",x"c1",x"4a",x"70"),
   349 => (x"c2",x"c0",x"05",x"aa"),
   350 => (x"c2",x"4d",x"c1",x"87"),
   351 => (x"c0",x"05",x"ad",x"b7"),
   352 => (x"17",x"27",x"87",x"d3"),
   353 => (x"1e",x"00",x"00",x"06"),
   354 => (x"00",x"00",x"61",x"27"),
   355 => (x"86",x"c4",x"0f",x"00"),
   356 => (x"f7",x"c1",x"48",x"c0"),
   357 => (x"75",x"8d",x"c1",x"87"),
   358 => (x"c9",x"fe",x"05",x"9d"),
   359 => (x"03",x"89",x"27",x"87"),
   360 => (x"27",x"0f",x"00",x"00"),
   361 => (x"00",x"00",x"02",x"25"),
   362 => (x"02",x"21",x"27",x"58"),
   363 => (x"05",x"bf",x"00",x"00"),
   364 => (x"c1",x"87",x"d0",x"c0"),
   365 => (x"f0",x"ff",x"c0",x"1e"),
   366 => (x"27",x"1e",x"d0",x"c1"),
   367 => (x"00",x"00",x"02",x"6b"),
   368 => (x"ff",x"86",x"c8",x"0f"),
   369 => (x"ff",x"c3",x"49",x"d4"),
   370 => (x"08",x"b2",x"27",x"79"),
   371 => (x"27",x"0f",x"00",x"00"),
   372 => (x"00",x"00",x"19",x"58"),
   373 => (x"19",x"54",x"27",x"58"),
   374 => (x"1e",x"bf",x"00",x"00"),
   375 => (x"00",x"06",x"20",x"27"),
   376 => (x"9a",x"27",x"1e",x"00"),
   377 => (x"0f",x"00",x"00",x"00"),
   378 => (x"48",x"6c",x"86",x"c8"),
   379 => (x"a6",x"c4",x"98",x"73"),
   380 => (x"c0",x"02",x"6e",x"58"),
   381 => (x"48",x"6c",x"87",x"cc"),
   382 => (x"a6",x"c4",x"98",x"73"),
   383 => (x"ff",x"05",x"6e",x"58"),
   384 => (x"7c",x"c0",x"87",x"f4"),
   385 => (x"c3",x"49",x"d4",x"ff"),
   386 => (x"48",x"c1",x"79",x"ff"),
   387 => (x"26",x"4d",x"26",x"26"),
   388 => (x"26",x"4b",x"26",x"4c"),
   389 => (x"49",x"4f",x"26",x"4a"),
   390 => (x"00",x"52",x"52",x"45"),
   391 => (x"00",x"49",x"50",x"53"),
   392 => (x"63",x"20",x"44",x"53"),
   393 => (x"20",x"64",x"72",x"61"),
   394 => (x"65",x"7a",x"69",x"73"),
   395 => (x"20",x"73",x"69",x"20"),
   396 => (x"00",x"0a",x"64",x"25"),
   397 => (x"5b",x"5a",x"5e",x"0e"),
   398 => (x"1e",x"0e",x"5d",x"5c"),
   399 => (x"ff",x"4d",x"ff",x"c3"),
   400 => (x"7c",x"75",x"4c",x"d4"),
   401 => (x"48",x"bf",x"d0",x"ff"),
   402 => (x"98",x"c0",x"c0",x"c8"),
   403 => (x"6e",x"58",x"a6",x"c4"),
   404 => (x"87",x"d2",x"c0",x"02"),
   405 => (x"4a",x"c0",x"c0",x"c8"),
   406 => (x"48",x"bf",x"d0",x"ff"),
   407 => (x"a6",x"c4",x"98",x"72"),
   408 => (x"ff",x"05",x"6e",x"58"),
   409 => (x"d0",x"ff",x"87",x"f2"),
   410 => (x"79",x"c1",x"c4",x"49"),
   411 => (x"66",x"d8",x"7c",x"75"),
   412 => (x"f0",x"ff",x"c0",x"1e"),
   413 => (x"27",x"1e",x"d8",x"c1"),
   414 => (x"00",x"00",x"02",x"6b"),
   415 => (x"70",x"86",x"c8",x"0f"),
   416 => (x"02",x"9a",x"72",x"4a"),
   417 => (x"27",x"87",x"d3",x"c0"),
   418 => (x"00",x"00",x"07",x"3c"),
   419 => (x"00",x"61",x"27",x"1e"),
   420 => (x"c4",x"0f",x"00",x"00"),
   421 => (x"c2",x"48",x"c1",x"86"),
   422 => (x"7c",x"75",x"87",x"d7"),
   423 => (x"76",x"7c",x"fe",x"c3"),
   424 => (x"dc",x"79",x"c0",x"49"),
   425 => (x"72",x"4a",x"bf",x"66"),
   426 => (x"2b",x"b7",x"d8",x"4b"),
   427 => (x"98",x"75",x"48",x"73"),
   428 => (x"4b",x"72",x"7c",x"70"),
   429 => (x"73",x"2b",x"b7",x"d0"),
   430 => (x"70",x"98",x"75",x"48"),
   431 => (x"c8",x"4b",x"72",x"7c"),
   432 => (x"48",x"73",x"2b",x"b7"),
   433 => (x"7c",x"70",x"98",x"75"),
   434 => (x"98",x"75",x"48",x"72"),
   435 => (x"66",x"dc",x"7c",x"70"),
   436 => (x"c0",x"80",x"c4",x"48"),
   437 => (x"6e",x"58",x"a6",x"e0"),
   438 => (x"c4",x"80",x"c1",x"48"),
   439 => (x"49",x"6e",x"58",x"a6"),
   440 => (x"a9",x"b7",x"c0",x"c2"),
   441 => (x"87",x"fb",x"fe",x"04"),
   442 => (x"7c",x"75",x"7c",x"75"),
   443 => (x"da",x"d8",x"7c",x"75"),
   444 => (x"7c",x"75",x"4b",x"e0"),
   445 => (x"9a",x"75",x"4a",x"6c"),
   446 => (x"c0",x"05",x"9a",x"72"),
   447 => (x"8b",x"c1",x"87",x"c8"),
   448 => (x"ff",x"05",x"9b",x"73"),
   449 => (x"7c",x"75",x"87",x"ec"),
   450 => (x"48",x"bf",x"d0",x"ff"),
   451 => (x"98",x"c0",x"c0",x"c8"),
   452 => (x"6e",x"58",x"a6",x"c4"),
   453 => (x"87",x"d2",x"c0",x"02"),
   454 => (x"4a",x"c0",x"c0",x"c8"),
   455 => (x"48",x"bf",x"d0",x"ff"),
   456 => (x"a6",x"c4",x"98",x"72"),
   457 => (x"ff",x"05",x"6e",x"58"),
   458 => (x"d0",x"ff",x"87",x"f2"),
   459 => (x"c0",x"79",x"c0",x"49"),
   460 => (x"4d",x"26",x"26",x"48"),
   461 => (x"4b",x"26",x"4c",x"26"),
   462 => (x"4f",x"26",x"4a",x"26"),
   463 => (x"74",x"69",x"72",x"57"),
   464 => (x"61",x"66",x"20",x"65"),
   465 => (x"64",x"65",x"6c",x"69"),
   466 => (x"5e",x"0e",x"00",x"0a"),
   467 => (x"5d",x"5c",x"5b",x"5a"),
   468 => (x"66",x"d8",x"1e",x"0e"),
   469 => (x"4b",x"66",x"dc",x"4c"),
   470 => (x"79",x"c0",x"49",x"76"),
   471 => (x"df",x"cd",x"ee",x"c5"),
   472 => (x"49",x"d4",x"ff",x"4d"),
   473 => (x"ff",x"79",x"ff",x"c3"),
   474 => (x"c3",x"4a",x"bf",x"d4"),
   475 => (x"fe",x"c3",x"9a",x"ff"),
   476 => (x"c1",x"05",x"aa",x"b7"),
   477 => (x"50",x"27",x"87",x"e5"),
   478 => (x"49",x"00",x"00",x"19"),
   479 => (x"b7",x"c4",x"79",x"c0"),
   480 => (x"e4",x"c0",x"04",x"ab"),
   481 => (x"02",x"25",x"27",x"87"),
   482 => (x"70",x"0f",x"00",x"00"),
   483 => (x"c4",x"7c",x"72",x"4a"),
   484 => (x"19",x"50",x"27",x"84"),
   485 => (x"48",x"bf",x"00",x"00"),
   486 => (x"54",x"27",x"80",x"72"),
   487 => (x"58",x"00",x"00",x"19"),
   488 => (x"b7",x"c4",x"8b",x"c4"),
   489 => (x"dc",x"ff",x"03",x"ab"),
   490 => (x"ab",x"b7",x"c0",x"87"),
   491 => (x"87",x"e5",x"c0",x"06"),
   492 => (x"c3",x"4d",x"d4",x"ff"),
   493 => (x"4a",x"6d",x"7d",x"ff"),
   494 => (x"c1",x"7c",x"97",x"72"),
   495 => (x"19",x"50",x"27",x"84"),
   496 => (x"48",x"bf",x"00",x"00"),
   497 => (x"54",x"27",x"80",x"72"),
   498 => (x"58",x"00",x"00",x"19"),
   499 => (x"b7",x"c0",x"8b",x"c1"),
   500 => (x"de",x"ff",x"01",x"ab"),
   501 => (x"76",x"4d",x"c1",x"87"),
   502 => (x"c1",x"79",x"c1",x"49"),
   503 => (x"05",x"9d",x"75",x"8d"),
   504 => (x"ff",x"87",x"fe",x"fd"),
   505 => (x"ff",x"c3",x"49",x"d4"),
   506 => (x"26",x"48",x"6e",x"79"),
   507 => (x"4c",x"26",x"4d",x"26"),
   508 => (x"4a",x"26",x"4b",x"26"),
   509 => (x"5e",x"0e",x"4f",x"26"),
   510 => (x"5d",x"5c",x"5b",x"5a"),
   511 => (x"d0",x"ff",x"1e",x"0e"),
   512 => (x"c0",x"c0",x"c8",x"4b"),
   513 => (x"ff",x"4c",x"c0",x"4a"),
   514 => (x"ff",x"c3",x"49",x"d4"),
   515 => (x"72",x"48",x"6b",x"79"),
   516 => (x"58",x"a6",x"c4",x"98"),
   517 => (x"cc",x"c0",x"02",x"6e"),
   518 => (x"72",x"48",x"6b",x"87"),
   519 => (x"58",x"a6",x"c4",x"98"),
   520 => (x"f4",x"ff",x"05",x"6e"),
   521 => (x"7b",x"c1",x"c4",x"87"),
   522 => (x"c3",x"49",x"d4",x"ff"),
   523 => (x"66",x"d8",x"79",x"ff"),
   524 => (x"f0",x"ff",x"c0",x"1e"),
   525 => (x"27",x"1e",x"d1",x"c1"),
   526 => (x"00",x"00",x"02",x"6b"),
   527 => (x"70",x"86",x"c8",x"0f"),
   528 => (x"02",x"9d",x"75",x"4d"),
   529 => (x"75",x"87",x"d6",x"c0"),
   530 => (x"1e",x"66",x"dc",x"1e"),
   531 => (x"00",x"08",x"92",x"27"),
   532 => (x"9a",x"27",x"1e",x"00"),
   533 => (x"0f",x"00",x"00",x"00"),
   534 => (x"e8",x"c0",x"86",x"cc"),
   535 => (x"1e",x"c0",x"c8",x"87"),
   536 => (x"1e",x"66",x"e0",x"c0"),
   537 => (x"c8",x"87",x"e3",x"fb"),
   538 => (x"6b",x"4c",x"70",x"86"),
   539 => (x"c4",x"98",x"72",x"48"),
   540 => (x"02",x"6e",x"58",x"a6"),
   541 => (x"6b",x"87",x"cc",x"c0"),
   542 => (x"c4",x"98",x"72",x"48"),
   543 => (x"05",x"6e",x"58",x"a6"),
   544 => (x"c0",x"87",x"f4",x"ff"),
   545 => (x"26",x"48",x"74",x"7b"),
   546 => (x"4c",x"26",x"4d",x"26"),
   547 => (x"4a",x"26",x"4b",x"26"),
   548 => (x"65",x"52",x"4f",x"26"),
   549 => (x"63",x"20",x"64",x"61"),
   550 => (x"61",x"6d",x"6d",x"6f"),
   551 => (x"66",x"20",x"64",x"6e"),
   552 => (x"65",x"6c",x"69",x"61"),
   553 => (x"74",x"61",x"20",x"64"),
   554 => (x"20",x"64",x"25",x"20"),
   555 => (x"29",x"64",x"25",x"28"),
   556 => (x"5e",x"0e",x"00",x"0a"),
   557 => (x"5d",x"5c",x"5b",x"5a"),
   558 => (x"1e",x"c0",x"1e",x"0e"),
   559 => (x"c1",x"f0",x"ff",x"c0"),
   560 => (x"6b",x"27",x"1e",x"c9"),
   561 => (x"0f",x"00",x"00",x"02"),
   562 => (x"1e",x"d2",x"86",x"c8"),
   563 => (x"00",x"19",x"60",x"27"),
   564 => (x"f5",x"f9",x"1e",x"00"),
   565 => (x"c0",x"86",x"c8",x"87"),
   566 => (x"d2",x"85",x"c1",x"4d"),
   567 => (x"ff",x"04",x"ad",x"b7"),
   568 => (x"60",x"27",x"87",x"f7"),
   569 => (x"97",x"00",x"00",x"19"),
   570 => (x"c0",x"c3",x"4a",x"bf"),
   571 => (x"b7",x"c0",x"c1",x"9a"),
   572 => (x"f2",x"c0",x"05",x"aa"),
   573 => (x"19",x"67",x"27",x"87"),
   574 => (x"bf",x"97",x"00",x"00"),
   575 => (x"27",x"32",x"d0",x"4a"),
   576 => (x"00",x"00",x"19",x"68"),
   577 => (x"c8",x"4b",x"bf",x"97"),
   578 => (x"73",x"4a",x"72",x"33"),
   579 => (x"19",x"69",x"27",x"b2"),
   580 => (x"bf",x"97",x"00",x"00"),
   581 => (x"73",x"4a",x"72",x"4b"),
   582 => (x"ff",x"ff",x"cf",x"b2"),
   583 => (x"4d",x"72",x"9a",x"ff"),
   584 => (x"35",x"ca",x"85",x"c1"),
   585 => (x"27",x"87",x"cb",x"c3"),
   586 => (x"00",x"00",x"19",x"69"),
   587 => (x"c1",x"4a",x"bf",x"97"),
   588 => (x"27",x"9a",x"c6",x"32"),
   589 => (x"00",x"00",x"19",x"6a"),
   590 => (x"c7",x"4b",x"bf",x"97"),
   591 => (x"4a",x"72",x"2b",x"b7"),
   592 => (x"65",x"27",x"b2",x"73"),
   593 => (x"97",x"00",x"00",x"19"),
   594 => (x"48",x"73",x"4b",x"bf"),
   595 => (x"a6",x"c4",x"98",x"cf"),
   596 => (x"19",x"66",x"27",x"58"),
   597 => (x"bf",x"97",x"00",x"00"),
   598 => (x"ca",x"9b",x"c3",x"4b"),
   599 => (x"19",x"67",x"27",x"33"),
   600 => (x"bf",x"97",x"00",x"00"),
   601 => (x"73",x"34",x"c2",x"4c"),
   602 => (x"27",x"b3",x"74",x"4b"),
   603 => (x"00",x"00",x"19",x"68"),
   604 => (x"c3",x"4c",x"bf",x"97"),
   605 => (x"b7",x"c6",x"9c",x"c0"),
   606 => (x"74",x"4b",x"73",x"2c"),
   607 => (x"c4",x"1e",x"73",x"b3"),
   608 => (x"1e",x"72",x"1e",x"66"),
   609 => (x"00",x"09",x"ff",x"27"),
   610 => (x"9a",x"27",x"1e",x"00"),
   611 => (x"0f",x"00",x"00",x"00"),
   612 => (x"82",x"c2",x"86",x"d0"),
   613 => (x"30",x"72",x"48",x"c1"),
   614 => (x"1e",x"72",x"4a",x"70"),
   615 => (x"00",x"0a",x"2c",x"27"),
   616 => (x"9a",x"27",x"1e",x"00"),
   617 => (x"0f",x"00",x"00",x"00"),
   618 => (x"48",x"c1",x"86",x"c8"),
   619 => (x"a6",x"c4",x"30",x"6e"),
   620 => (x"73",x"83",x"c1",x"58"),
   621 => (x"6e",x"95",x"72",x"4d"),
   622 => (x"27",x"1e",x"75",x"1e"),
   623 => (x"00",x"00",x"0a",x"35"),
   624 => (x"00",x"9a",x"27",x"1e"),
   625 => (x"cc",x"0f",x"00",x"00"),
   626 => (x"c8",x"49",x"6e",x"86"),
   627 => (x"06",x"a9",x"b7",x"c0"),
   628 => (x"6e",x"87",x"cf",x"c0"),
   629 => (x"c1",x"35",x"c1",x"4a"),
   630 => (x"c0",x"c8",x"2a",x"b7"),
   631 => (x"ff",x"01",x"aa",x"b7"),
   632 => (x"1e",x"75",x"87",x"f3"),
   633 => (x"00",x"0a",x"4b",x"27"),
   634 => (x"9a",x"27",x"1e",x"00"),
   635 => (x"0f",x"00",x"00",x"00"),
   636 => (x"48",x"75",x"86",x"c8"),
   637 => (x"26",x"4d",x"26",x"26"),
   638 => (x"26",x"4b",x"26",x"4c"),
   639 => (x"63",x"4f",x"26",x"4a"),
   640 => (x"7a",x"69",x"73",x"5f"),
   641 => (x"75",x"6d",x"5f",x"65"),
   642 => (x"20",x"3a",x"74",x"6c"),
   643 => (x"20",x"2c",x"64",x"25"),
   644 => (x"64",x"61",x"65",x"72"),
   645 => (x"5f",x"6c",x"62",x"5f"),
   646 => (x"3a",x"6e",x"65",x"6c"),
   647 => (x"2c",x"64",x"25",x"20"),
   648 => (x"69",x"73",x"63",x"20"),
   649 => (x"20",x"3a",x"65",x"7a"),
   650 => (x"00",x"0a",x"64",x"25"),
   651 => (x"74",x"6c",x"75",x"4d"),
   652 => (x"0a",x"64",x"25",x"20"),
   653 => (x"20",x"64",x"25",x"00"),
   654 => (x"63",x"6f",x"6c",x"62"),
   655 => (x"6f",x"20",x"73",x"6b"),
   656 => (x"69",x"73",x"20",x"66"),
   657 => (x"25",x"20",x"65",x"7a"),
   658 => (x"25",x"00",x"0a",x"64"),
   659 => (x"6c",x"62",x"20",x"64"),
   660 => (x"73",x"6b",x"63",x"6f"),
   661 => (x"20",x"66",x"6f",x"20"),
   662 => (x"20",x"32",x"31",x"35"),
   663 => (x"65",x"74",x"79",x"62"),
   664 => (x"0e",x"00",x"0a",x"73"),
   665 => (x"5c",x"5b",x"5a",x"5e"),
   666 => (x"66",x"d4",x"0e",x"5d"),
   667 => (x"dc",x"4c",x"c0",x"4d"),
   668 => (x"b7",x"c0",x"49",x"66"),
   669 => (x"fb",x"c0",x"06",x"a9"),
   670 => (x"c1",x"4b",x"15",x"87"),
   671 => (x"c0",x"c0",x"c0",x"c0"),
   672 => (x"b7",x"c0",x"c4",x"93"),
   673 => (x"66",x"d8",x"4b",x"93"),
   674 => (x"c1",x"4a",x"bf",x"97"),
   675 => (x"c0",x"c0",x"c0",x"c0"),
   676 => (x"b7",x"c0",x"c4",x"92"),
   677 => (x"66",x"d8",x"4a",x"92"),
   678 => (x"dc",x"80",x"c1",x"48"),
   679 => (x"b7",x"72",x"58",x"a6"),
   680 => (x"c5",x"c0",x"02",x"ab"),
   681 => (x"c0",x"48",x"c1",x"87"),
   682 => (x"84",x"c1",x"87",x"cc"),
   683 => (x"ac",x"b7",x"66",x"dc"),
   684 => (x"87",x"c5",x"ff",x"04"),
   685 => (x"4d",x"26",x"48",x"c0"),
   686 => (x"4b",x"26",x"4c",x"26"),
   687 => (x"4f",x"26",x"4a",x"26"),
   688 => (x"5b",x"5a",x"5e",x"0e"),
   689 => (x"27",x"0e",x"5d",x"5c"),
   690 => (x"00",x"00",x"1b",x"80"),
   691 => (x"27",x"79",x"c0",x"49"),
   692 => (x"00",x"00",x"18",x"94"),
   693 => (x"00",x"61",x"27",x"1e"),
   694 => (x"c4",x"0f",x"00",x"00"),
   695 => (x"19",x"78",x"27",x"86"),
   696 => (x"c0",x"1e",x"00",x"00"),
   697 => (x"07",x"f6",x"27",x"1e"),
   698 => (x"c8",x"0f",x"00",x"00"),
   699 => (x"72",x"4a",x"70",x"86"),
   700 => (x"d3",x"c0",x"05",x"9a"),
   701 => (x"17",x"c0",x"27",x"87"),
   702 => (x"27",x"1e",x"00",x"00"),
   703 => (x"00",x"00",x"00",x"61"),
   704 => (x"c0",x"86",x"c4",x"0f"),
   705 => (x"87",x"e6",x"d0",x"48"),
   706 => (x"00",x"18",x"a1",x"27"),
   707 => (x"61",x"27",x"1e",x"00"),
   708 => (x"0f",x"00",x"00",x"00"),
   709 => (x"4c",x"c0",x"86",x"c4"),
   710 => (x"00",x"1b",x"ac",x"27"),
   711 => (x"79",x"c1",x"49",x"00"),
   712 => (x"b8",x"27",x"1e",x"c8"),
   713 => (x"1e",x"00",x"00",x"18"),
   714 => (x"00",x"19",x"ae",x"27"),
   715 => (x"63",x"27",x"1e",x"00"),
   716 => (x"0f",x"00",x"00",x"0a"),
   717 => (x"4a",x"70",x"86",x"cc"),
   718 => (x"c0",x"05",x"9a",x"72"),
   719 => (x"ac",x"27",x"87",x"c8"),
   720 => (x"49",x"00",x"00",x"1b"),
   721 => (x"1e",x"c8",x"79",x"c0"),
   722 => (x"00",x"18",x"c1",x"27"),
   723 => (x"ca",x"27",x"1e",x"00"),
   724 => (x"1e",x"00",x"00",x"19"),
   725 => (x"00",x"0a",x"63",x"27"),
   726 => (x"86",x"cc",x"0f",x"00"),
   727 => (x"9a",x"72",x"4a",x"70"),
   728 => (x"87",x"c8",x"c0",x"05"),
   729 => (x"00",x"1b",x"ac",x"27"),
   730 => (x"79",x"c0",x"49",x"00"),
   731 => (x"00",x"1b",x"ac",x"27"),
   732 => (x"27",x"1e",x"bf",x"00"),
   733 => (x"00",x"00",x"18",x"ca"),
   734 => (x"00",x"9a",x"27",x"1e"),
   735 => (x"c8",x"0f",x"00",x"00"),
   736 => (x"1b",x"ac",x"27",x"86"),
   737 => (x"02",x"bf",x"00",x"00"),
   738 => (x"27",x"87",x"cc",x"c3"),
   739 => (x"00",x"00",x"19",x"78"),
   740 => (x"1b",x"36",x"27",x"4d"),
   741 => (x"27",x"4b",x"00",x"00"),
   742 => (x"00",x"00",x"1b",x"76"),
   743 => (x"cf",x"4a",x"bf",x"9f"),
   744 => (x"72",x"9a",x"ff",x"ff"),
   745 => (x"1b",x"76",x"27",x"1e"),
   746 => (x"27",x"4a",x"00",x"00"),
   747 => (x"00",x"00",x"19",x"78"),
   748 => (x"d0",x"1e",x"72",x"8a"),
   749 => (x"1e",x"c0",x"c8",x"1e"),
   750 => (x"00",x"17",x"f2",x"27"),
   751 => (x"9a",x"27",x"1e",x"00"),
   752 => (x"0f",x"00",x"00",x"00"),
   753 => (x"4a",x"73",x"86",x"d4"),
   754 => (x"4c",x"6a",x"82",x"c8"),
   755 => (x"00",x"1b",x"76",x"27"),
   756 => (x"4a",x"bf",x"9f",x"00"),
   757 => (x"9a",x"ff",x"ff",x"cf"),
   758 => (x"b7",x"ea",x"d6",x"c5"),
   759 => (x"d3",x"c0",x"05",x"aa"),
   760 => (x"c8",x"4a",x"73",x"87"),
   761 => (x"27",x"1e",x"6a",x"82"),
   762 => (x"00",x"00",x"12",x"ae"),
   763 => (x"70",x"86",x"c4",x"0f"),
   764 => (x"87",x"e8",x"c0",x"4c"),
   765 => (x"fe",x"c7",x"4a",x"75"),
   766 => (x"4a",x"6a",x"9f",x"82"),
   767 => (x"9a",x"ff",x"ff",x"cf"),
   768 => (x"b7",x"d5",x"e9",x"ca"),
   769 => (x"d3",x"c0",x"02",x"aa"),
   770 => (x"17",x"d4",x"27",x"87"),
   771 => (x"27",x"1e",x"00",x"00"),
   772 => (x"00",x"00",x"00",x"61"),
   773 => (x"c0",x"86",x"c4",x"0f"),
   774 => (x"87",x"d2",x"cc",x"48"),
   775 => (x"2f",x"27",x"1e",x"74"),
   776 => (x"1e",x"00",x"00",x"18"),
   777 => (x"00",x"00",x"9a",x"27"),
   778 => (x"86",x"c8",x"0f",x"00"),
   779 => (x"00",x"19",x"78",x"27"),
   780 => (x"1e",x"74",x"1e",x"00"),
   781 => (x"00",x"07",x"f6",x"27"),
   782 => (x"86",x"c8",x"0f",x"00"),
   783 => (x"9a",x"72",x"4a",x"70"),
   784 => (x"87",x"c5",x"c0",x"05"),
   785 => (x"e5",x"cb",x"48",x"c0"),
   786 => (x"18",x"47",x"27",x"87"),
   787 => (x"27",x"1e",x"00",x"00"),
   788 => (x"00",x"00",x"00",x"61"),
   789 => (x"27",x"86",x"c4",x"0f"),
   790 => (x"00",x"00",x"18",x"dd"),
   791 => (x"00",x"9a",x"27",x"1e"),
   792 => (x"c4",x"0f",x"00",x"00"),
   793 => (x"27",x"1e",x"c8",x"86"),
   794 => (x"00",x"00",x"18",x"f5"),
   795 => (x"19",x"ca",x"27",x"1e"),
   796 => (x"27",x"1e",x"00",x"00"),
   797 => (x"00",x"00",x"0a",x"63"),
   798 => (x"70",x"86",x"cc",x"0f"),
   799 => (x"05",x"9a",x"72",x"4a"),
   800 => (x"27",x"87",x"cb",x"c0"),
   801 => (x"00",x"00",x"1b",x"80"),
   802 => (x"c0",x"79",x"c1",x"49"),
   803 => (x"1e",x"c8",x"87",x"f1"),
   804 => (x"00",x"18",x"fe",x"27"),
   805 => (x"ae",x"27",x"1e",x"00"),
   806 => (x"1e",x"00",x"00",x"19"),
   807 => (x"00",x"0a",x"63",x"27"),
   808 => (x"86",x"cc",x"0f",x"00"),
   809 => (x"9a",x"72",x"4a",x"70"),
   810 => (x"87",x"d3",x"c0",x"02"),
   811 => (x"00",x"18",x"6e",x"27"),
   812 => (x"9a",x"27",x"1e",x"00"),
   813 => (x"0f",x"00",x"00",x"00"),
   814 => (x"48",x"c0",x"86",x"c4"),
   815 => (x"27",x"87",x"ef",x"c9"),
   816 => (x"00",x"00",x"1b",x"76"),
   817 => (x"c3",x"4a",x"bf",x"97"),
   818 => (x"d5",x"c1",x"9a",x"ff"),
   819 => (x"c0",x"05",x"aa",x"b7"),
   820 => (x"77",x"27",x"87",x"d3"),
   821 => (x"97",x"00",x"00",x"1b"),
   822 => (x"ff",x"c3",x"4a",x"bf"),
   823 => (x"b7",x"ea",x"c2",x"9a"),
   824 => (x"c5",x"c0",x"02",x"aa"),
   825 => (x"c9",x"48",x"c0",x"87"),
   826 => (x"78",x"27",x"87",x"c4"),
   827 => (x"97",x"00",x"00",x"19"),
   828 => (x"ff",x"c3",x"4a",x"bf"),
   829 => (x"b7",x"e9",x"c3",x"9a"),
   830 => (x"d8",x"c0",x"02",x"aa"),
   831 => (x"19",x"78",x"27",x"87"),
   832 => (x"bf",x"97",x"00",x"00"),
   833 => (x"9a",x"ff",x"c3",x"4a"),
   834 => (x"aa",x"b7",x"eb",x"c3"),
   835 => (x"87",x"c5",x"c0",x"02"),
   836 => (x"d9",x"c8",x"48",x"c0"),
   837 => (x"19",x"83",x"27",x"87"),
   838 => (x"bf",x"97",x"00",x"00"),
   839 => (x"9a",x"ff",x"c3",x"4a"),
   840 => (x"c0",x"05",x"9a",x"72"),
   841 => (x"84",x"27",x"87",x"d2"),
   842 => (x"97",x"00",x"00",x"19"),
   843 => (x"ff",x"c3",x"4a",x"bf"),
   844 => (x"aa",x"b7",x"c2",x"9a"),
   845 => (x"87",x"c5",x"c0",x"02"),
   846 => (x"f1",x"c7",x"48",x"c0"),
   847 => (x"19",x"85",x"27",x"87"),
   848 => (x"bf",x"97",x"00",x"00"),
   849 => (x"98",x"ff",x"c3",x"48"),
   850 => (x"00",x"1b",x"7c",x"27"),
   851 => (x"78",x"27",x"58",x"00"),
   852 => (x"bf",x"00",x"00",x"1b"),
   853 => (x"c1",x"4b",x"72",x"4a"),
   854 => (x"1b",x"7c",x"27",x"8b"),
   855 => (x"73",x"49",x"00",x"00"),
   856 => (x"72",x"1e",x"73",x"79"),
   857 => (x"19",x"07",x"27",x"1e"),
   858 => (x"27",x"1e",x"00",x"00"),
   859 => (x"00",x"00",x"00",x"9a"),
   860 => (x"27",x"86",x"cc",x"0f"),
   861 => (x"00",x"00",x"19",x"86"),
   862 => (x"c3",x"4a",x"bf",x"97"),
   863 => (x"82",x"74",x"9a",x"ff"),
   864 => (x"00",x"19",x"87",x"27"),
   865 => (x"4b",x"bf",x"97",x"00"),
   866 => (x"c8",x"9b",x"ff",x"c3"),
   867 => (x"72",x"48",x"73",x"33"),
   868 => (x"1b",x"90",x"27",x"80"),
   869 => (x"27",x"58",x"00",x"00"),
   870 => (x"00",x"00",x"19",x"88"),
   871 => (x"c3",x"48",x"bf",x"97"),
   872 => (x"a4",x"27",x"98",x"ff"),
   873 => (x"58",x"00",x"00",x"1b"),
   874 => (x"00",x"1b",x"80",x"27"),
   875 => (x"c3",x"02",x"bf",x"00"),
   876 => (x"1e",x"c8",x"87",x"f7"),
   877 => (x"00",x"18",x"8b",x"27"),
   878 => (x"ca",x"27",x"1e",x"00"),
   879 => (x"1e",x"00",x"00",x"19"),
   880 => (x"00",x"0a",x"63",x"27"),
   881 => (x"86",x"cc",x"0f",x"00"),
   882 => (x"9a",x"72",x"4a",x"70"),
   883 => (x"87",x"c5",x"c0",x"02"),
   884 => (x"d9",x"c5",x"48",x"c0"),
   885 => (x"1b",x"78",x"27",x"87"),
   886 => (x"4b",x"bf",x"00",x"00"),
   887 => (x"30",x"c4",x"48",x"73"),
   888 => (x"00",x"1b",x"a8",x"27"),
   889 => (x"9c",x"27",x"58",x"00"),
   890 => (x"49",x"00",x"00",x"1b"),
   891 => (x"9d",x"27",x"79",x"73"),
   892 => (x"97",x"00",x"00",x"19"),
   893 => (x"ff",x"c3",x"4a",x"bf"),
   894 => (x"27",x"32",x"c8",x"9a"),
   895 => (x"00",x"00",x"19",x"9c"),
   896 => (x"c3",x"4c",x"bf",x"97"),
   897 => (x"4a",x"72",x"9c",x"ff"),
   898 => (x"9e",x"27",x"82",x"74"),
   899 => (x"97",x"00",x"00",x"19"),
   900 => (x"ff",x"c3",x"4c",x"bf"),
   901 => (x"72",x"34",x"d0",x"9c"),
   902 => (x"27",x"82",x"74",x"4a"),
   903 => (x"00",x"00",x"19",x"9f"),
   904 => (x"c3",x"4c",x"bf",x"97"),
   905 => (x"34",x"d8",x"9c",x"ff"),
   906 => (x"82",x"74",x"4a",x"72"),
   907 => (x"00",x"1b",x"a8",x"27"),
   908 => (x"79",x"72",x"49",x"00"),
   909 => (x"a0",x"27",x"4a",x"72"),
   910 => (x"bf",x"00",x"00",x"1b"),
   911 => (x"27",x"4a",x"72",x"92"),
   912 => (x"00",x"00",x"1b",x"8c"),
   913 => (x"90",x"27",x"82",x"bf"),
   914 => (x"49",x"00",x"00",x"1b"),
   915 => (x"a5",x"27",x"79",x"72"),
   916 => (x"97",x"00",x"00",x"19"),
   917 => (x"ff",x"c3",x"4c",x"bf"),
   918 => (x"27",x"34",x"c8",x"9c"),
   919 => (x"00",x"00",x"19",x"a4"),
   920 => (x"c3",x"4d",x"bf",x"97"),
   921 => (x"4c",x"74",x"9d",x"ff"),
   922 => (x"a6",x"27",x"84",x"75"),
   923 => (x"97",x"00",x"00",x"19"),
   924 => (x"ff",x"c3",x"4d",x"bf"),
   925 => (x"74",x"35",x"d0",x"9d"),
   926 => (x"27",x"84",x"75",x"4c"),
   927 => (x"00",x"00",x"19",x"a7"),
   928 => (x"c3",x"4d",x"bf",x"97"),
   929 => (x"9d",x"cf",x"9d",x"ff"),
   930 => (x"4c",x"74",x"35",x"d8"),
   931 => (x"94",x"27",x"84",x"75"),
   932 => (x"49",x"00",x"00",x"1b"),
   933 => (x"8c",x"c2",x"79",x"74"),
   934 => (x"93",x"74",x"4b",x"73"),
   935 => (x"80",x"72",x"48",x"73"),
   936 => (x"00",x"1b",x"9c",x"27"),
   937 => (x"c3",x"c2",x"58",x"00"),
   938 => (x"19",x"8a",x"27",x"87"),
   939 => (x"bf",x"97",x"00",x"00"),
   940 => (x"9a",x"ff",x"c3",x"4a"),
   941 => (x"89",x"27",x"32",x"c8"),
   942 => (x"97",x"00",x"00",x"19"),
   943 => (x"ff",x"c3",x"4b",x"bf"),
   944 => (x"73",x"4a",x"72",x"9b"),
   945 => (x"1b",x"a4",x"27",x"82"),
   946 => (x"72",x"49",x"00",x"00"),
   947 => (x"c7",x"32",x"c5",x"79"),
   948 => (x"2a",x"c9",x"82",x"ff"),
   949 => (x"00",x"1b",x"9c",x"27"),
   950 => (x"79",x"72",x"49",x"00"),
   951 => (x"00",x"19",x"8f",x"27"),
   952 => (x"4b",x"bf",x"97",x"00"),
   953 => (x"c8",x"9b",x"ff",x"c3"),
   954 => (x"19",x"8e",x"27",x"33"),
   955 => (x"bf",x"97",x"00",x"00"),
   956 => (x"9c",x"ff",x"c3",x"4c"),
   957 => (x"83",x"74",x"4b",x"73"),
   958 => (x"00",x"1b",x"a8",x"27"),
   959 => (x"79",x"73",x"49",x"00"),
   960 => (x"a0",x"27",x"4b",x"73"),
   961 => (x"bf",x"00",x"00",x"1b"),
   962 => (x"27",x"4b",x"73",x"93"),
   963 => (x"00",x"00",x"1b",x"8c"),
   964 => (x"98",x"27",x"83",x"bf"),
   965 => (x"49",x"00",x"00",x"1b"),
   966 => (x"94",x"27",x"79",x"73"),
   967 => (x"49",x"00",x"00",x"1b"),
   968 => (x"48",x"73",x"79",x"c0"),
   969 => (x"94",x"27",x"80",x"72"),
   970 => (x"58",x"00",x"00",x"1b"),
   971 => (x"4d",x"26",x"48",x"c1"),
   972 => (x"4b",x"26",x"4c",x"26"),
   973 => (x"4f",x"26",x"4a",x"26"),
   974 => (x"5b",x"5a",x"5e",x"0e"),
   975 => (x"27",x"0e",x"5d",x"5c"),
   976 => (x"00",x"00",x"1b",x"80"),
   977 => (x"cf",x"c0",x"02",x"bf"),
   978 => (x"4d",x"66",x"d4",x"87"),
   979 => (x"d4",x"2d",x"b7",x"c7"),
   980 => (x"ff",x"c1",x"4b",x"66"),
   981 => (x"87",x"cc",x"c0",x"9b"),
   982 => (x"c8",x"4d",x"66",x"d4"),
   983 => (x"66",x"d4",x"2d",x"b7"),
   984 => (x"9b",x"ff",x"c3",x"4b"),
   985 => (x"00",x"19",x"78",x"27"),
   986 => (x"8c",x"27",x"1e",x"00"),
   987 => (x"bf",x"00",x"00",x"1b"),
   988 => (x"72",x"82",x"75",x"4a"),
   989 => (x"07",x"f6",x"27",x"1e"),
   990 => (x"c8",x"0f",x"00",x"00"),
   991 => (x"72",x"4a",x"70",x"86"),
   992 => (x"c5",x"c0",x"05",x"9a"),
   993 => (x"c0",x"48",x"c0",x"87"),
   994 => (x"80",x"27",x"87",x"f6"),
   995 => (x"bf",x"00",x"00",x"1b"),
   996 => (x"87",x"d7",x"c0",x"02"),
   997 => (x"92",x"c4",x"4a",x"73"),
   998 => (x"78",x"27",x"4a",x"72"),
   999 => (x"82",x"00",x"00",x"19"),
  1000 => (x"ff",x"cf",x"4c",x"6a"),
  1001 => (x"9c",x"ff",x"ff",x"ff"),
  1002 => (x"73",x"87",x"d3",x"c0"),
  1003 => (x"72",x"92",x"c2",x"4a"),
  1004 => (x"19",x"78",x"27",x"4a"),
  1005 => (x"9f",x"82",x"00",x"00"),
  1006 => (x"ff",x"cf",x"4c",x"6a"),
  1007 => (x"48",x"74",x"9c",x"ff"),
  1008 => (x"4c",x"26",x"4d",x"26"),
  1009 => (x"4a",x"26",x"4b",x"26"),
  1010 => (x"5e",x"0e",x"4f",x"26"),
  1011 => (x"5d",x"5c",x"5b",x"5a"),
  1012 => (x"cf",x"8e",x"cc",x"0e"),
  1013 => (x"f8",x"ff",x"ff",x"ff"),
  1014 => (x"76",x"4c",x"c0",x"4d"),
  1015 => (x"1b",x"94",x"27",x"49"),
  1016 => (x"79",x"bf",x"00",x"00"),
  1017 => (x"27",x"49",x"a6",x"c4"),
  1018 => (x"00",x"00",x"1b",x"98"),
  1019 => (x"80",x"27",x"79",x"bf"),
  1020 => (x"bf",x"00",x"00",x"1b"),
  1021 => (x"87",x"cc",x"c0",x"02"),
  1022 => (x"00",x"1b",x"78",x"27"),
  1023 => (x"c4",x"4a",x"bf",x"00"),
  1024 => (x"87",x"c9",x"c0",x"32"),
  1025 => (x"00",x"1b",x"9c",x"27"),
  1026 => (x"c4",x"4a",x"bf",x"00"),
  1027 => (x"49",x"a6",x"c8",x"32"),
  1028 => (x"4b",x"c0",x"79",x"72"),
  1029 => (x"c0",x"49",x"66",x"c8"),
  1030 => (x"e1",x"c3",x"06",x"a9"),
  1031 => (x"cf",x"4a",x"73",x"87"),
  1032 => (x"05",x"9a",x"72",x"9a"),
  1033 => (x"27",x"87",x"e4",x"c0"),
  1034 => (x"00",x"00",x"19",x"78"),
  1035 => (x"4a",x"66",x"c8",x"1e"),
  1036 => (x"c1",x"48",x"66",x"c8"),
  1037 => (x"58",x"a6",x"cc",x"80"),
  1038 => (x"f6",x"27",x"1e",x"72"),
  1039 => (x"0f",x"00",x"00",x"07"),
  1040 => (x"78",x"27",x"86",x"c8"),
  1041 => (x"4c",x"00",x"00",x"19"),
  1042 => (x"c0",x"87",x"c3",x"c0"),
  1043 => (x"6c",x"97",x"84",x"e0"),
  1044 => (x"9a",x"ff",x"c3",x"4a"),
  1045 => (x"c2",x"02",x"9a",x"72"),
  1046 => (x"6c",x"97",x"87",x"db"),
  1047 => (x"9a",x"ff",x"c3",x"4a"),
  1048 => (x"aa",x"b7",x"e5",x"c3"),
  1049 => (x"87",x"cd",x"c2",x"02"),
  1050 => (x"82",x"cb",x"4a",x"74"),
  1051 => (x"c3",x"4a",x"6a",x"97"),
  1052 => (x"9a",x"d8",x"9a",x"ff"),
  1053 => (x"c1",x"05",x"9a",x"72"),
  1054 => (x"1e",x"74",x"87",x"fb"),
  1055 => (x"00",x"00",x"61",x"27"),
  1056 => (x"86",x"c4",x"0f",x"00"),
  1057 => (x"e8",x"c0",x"1e",x"cb"),
  1058 => (x"1e",x"74",x"1e",x"66"),
  1059 => (x"00",x"0a",x"63",x"27"),
  1060 => (x"86",x"cc",x"0f",x"00"),
  1061 => (x"9a",x"72",x"4a",x"70"),
  1062 => (x"87",x"d9",x"c1",x"05"),
  1063 => (x"83",x"dc",x"4b",x"74"),
  1064 => (x"4a",x"66",x"e0",x"c0"),
  1065 => (x"7a",x"6b",x"82",x"c4"),
  1066 => (x"83",x"da",x"4b",x"74"),
  1067 => (x"4a",x"66",x"e0",x"c0"),
  1068 => (x"6b",x"9f",x"82",x"c8"),
  1069 => (x"ff",x"ff",x"cf",x"48"),
  1070 => (x"72",x"7a",x"70",x"98"),
  1071 => (x"1b",x"80",x"27",x"4d"),
  1072 => (x"02",x"bf",x"00",x"00"),
  1073 => (x"74",x"87",x"d9",x"c0"),
  1074 => (x"9f",x"82",x"d4",x"4a"),
  1075 => (x"ff",x"cf",x"4a",x"6a"),
  1076 => (x"ff",x"c0",x"9a",x"ff"),
  1077 => (x"48",x"72",x"9a",x"ff"),
  1078 => (x"a6",x"c4",x"30",x"d0"),
  1079 => (x"87",x"c4",x"c0",x"58"),
  1080 => (x"79",x"c0",x"49",x"76"),
  1081 => (x"80",x"6d",x"48",x"6e"),
  1082 => (x"e0",x"c0",x"7d",x"70"),
  1083 => (x"79",x"c0",x"49",x"66"),
  1084 => (x"ce",x"c1",x"48",x"c1"),
  1085 => (x"c8",x"83",x"c1",x"87"),
  1086 => (x"fc",x"04",x"ab",x"66"),
  1087 => (x"ff",x"cf",x"87",x"df"),
  1088 => (x"4d",x"f8",x"ff",x"ff"),
  1089 => (x"00",x"1b",x"80",x"27"),
  1090 => (x"c0",x"02",x"bf",x"00"),
  1091 => (x"1e",x"6e",x"87",x"f3"),
  1092 => (x"00",x"0f",x"38",x"27"),
  1093 => (x"86",x"c4",x"0f",x"00"),
  1094 => (x"6e",x"58",x"a6",x"c4"),
  1095 => (x"75",x"9a",x"75",x"4a"),
  1096 => (x"dc",x"c0",x"02",x"aa"),
  1097 => (x"c2",x"4a",x"6e",x"87"),
  1098 => (x"27",x"4a",x"72",x"8a"),
  1099 => (x"00",x"00",x"1b",x"78"),
  1100 => (x"90",x"27",x"92",x"bf"),
  1101 => (x"bf",x"00",x"00",x"1b"),
  1102 => (x"c8",x"80",x"72",x"48"),
  1103 => (x"d1",x"fb",x"58",x"a6"),
  1104 => (x"cf",x"48",x"c0",x"87"),
  1105 => (x"f8",x"ff",x"ff",x"ff"),
  1106 => (x"26",x"86",x"cc",x"4d"),
  1107 => (x"26",x"4c",x"26",x"4d"),
  1108 => (x"26",x"4a",x"26",x"4b"),
  1109 => (x"5a",x"5e",x"0e",x"4f"),
  1110 => (x"66",x"cc",x"0e",x"5b"),
  1111 => (x"82",x"c1",x"4a",x"bf"),
  1112 => (x"72",x"49",x"66",x"cc"),
  1113 => (x"27",x"4a",x"72",x"79"),
  1114 => (x"00",x"00",x"1b",x"7c"),
  1115 => (x"9a",x"72",x"9a",x"bf"),
  1116 => (x"87",x"d3",x"c0",x"05"),
  1117 => (x"c8",x"4a",x"66",x"cc"),
  1118 => (x"27",x"1e",x"6a",x"82"),
  1119 => (x"00",x"00",x"0f",x"38"),
  1120 => (x"70",x"86",x"c4",x"0f"),
  1121 => (x"c1",x"7a",x"73",x"4b"),
  1122 => (x"26",x"4b",x"26",x"48"),
  1123 => (x"0e",x"4f",x"26",x"4a"),
  1124 => (x"0e",x"5b",x"5a",x"5e"),
  1125 => (x"00",x"1b",x"90",x"27"),
  1126 => (x"cc",x"4a",x"bf",x"00"),
  1127 => (x"83",x"c8",x"4b",x"66"),
  1128 => (x"8b",x"c2",x"4b",x"6b"),
  1129 => (x"78",x"27",x"4b",x"73"),
  1130 => (x"bf",x"00",x"00",x"1b"),
  1131 => (x"73",x"4a",x"72",x"93"),
  1132 => (x"1b",x"7c",x"27",x"82"),
  1133 => (x"4b",x"bf",x"00",x"00"),
  1134 => (x"9b",x"bf",x"66",x"cc"),
  1135 => (x"82",x"73",x"4a",x"72"),
  1136 => (x"72",x"1e",x"66",x"d0"),
  1137 => (x"07",x"f6",x"27",x"1e"),
  1138 => (x"c8",x"0f",x"00",x"00"),
  1139 => (x"72",x"4a",x"70",x"86"),
  1140 => (x"c5",x"c0",x"05",x"9a"),
  1141 => (x"c0",x"48",x"c0",x"87"),
  1142 => (x"48",x"c1",x"87",x"c2"),
  1143 => (x"4a",x"26",x"4b",x"26"),
  1144 => (x"5e",x"0e",x"4f",x"26"),
  1145 => (x"5d",x"5c",x"5b",x"5a"),
  1146 => (x"4c",x"66",x"d8",x"0e"),
  1147 => (x"27",x"1e",x"66",x"d4"),
  1148 => (x"00",x"00",x"1b",x"b0"),
  1149 => (x"0f",x"ca",x"27",x"1e"),
  1150 => (x"c8",x"0f",x"00",x"00"),
  1151 => (x"72",x"4a",x"70",x"86"),
  1152 => (x"df",x"c1",x"02",x"9a"),
  1153 => (x"1b",x"b4",x"27",x"87"),
  1154 => (x"4a",x"bf",x"00",x"00"),
  1155 => (x"c9",x"82",x"ff",x"c7"),
  1156 => (x"c0",x"4d",x"72",x"2a"),
  1157 => (x"12",x"86",x"27",x"4b"),
  1158 => (x"27",x"1e",x"00",x"00"),
  1159 => (x"00",x"00",x"00",x"61"),
  1160 => (x"c0",x"86",x"c4",x"0f"),
  1161 => (x"c1",x"06",x"ad",x"b7"),
  1162 => (x"1e",x"74",x"87",x"d0"),
  1163 => (x"00",x"1b",x"b0",x"27"),
  1164 => (x"8f",x"27",x"1e",x"00"),
  1165 => (x"0f",x"00",x"00",x"11"),
  1166 => (x"4a",x"70",x"86",x"c8"),
  1167 => (x"c0",x"05",x"9a",x"72"),
  1168 => (x"48",x"c0",x"87",x"c5"),
  1169 => (x"27",x"87",x"f5",x"c0"),
  1170 => (x"00",x"00",x"1b",x"b0"),
  1171 => (x"11",x"55",x"27",x"1e"),
  1172 => (x"c4",x"0f",x"00",x"00"),
  1173 => (x"84",x"c0",x"c8",x"86"),
  1174 => (x"b7",x"75",x"83",x"c1"),
  1175 => (x"c9",x"ff",x"04",x"ab"),
  1176 => (x"87",x"d6",x"c0",x"87"),
  1177 => (x"27",x"1e",x"66",x"d4"),
  1178 => (x"00",x"00",x"12",x"9f"),
  1179 => (x"00",x"9a",x"27",x"1e"),
  1180 => (x"c8",x"0f",x"00",x"00"),
  1181 => (x"c0",x"48",x"c0",x"86"),
  1182 => (x"48",x"c1",x"87",x"c2"),
  1183 => (x"4c",x"26",x"4d",x"26"),
  1184 => (x"4a",x"26",x"4b",x"26"),
  1185 => (x"70",x"4f",x"4f",x"26"),
  1186 => (x"64",x"65",x"6e",x"65"),
  1187 => (x"6c",x"69",x"66",x"20"),
  1188 => (x"6c",x"20",x"2c",x"65"),
  1189 => (x"69",x"64",x"61",x"6f"),
  1190 => (x"2e",x"2e",x"67",x"6e"),
  1191 => (x"43",x"00",x"0a",x"2e"),
  1192 => (x"74",x"27",x"6e",x"61"),
  1193 => (x"65",x"70",x"6f",x"20"),
  1194 => (x"73",x"25",x"20",x"6e"),
  1195 => (x"5e",x"0e",x"00",x"0a"),
  1196 => (x"cc",x"0e",x"5b",x"5a"),
  1197 => (x"2a",x"d8",x"4a",x"66"),
  1198 => (x"cc",x"9a",x"ff",x"c3"),
  1199 => (x"2b",x"c8",x"4b",x"66"),
  1200 => (x"9b",x"c0",x"fc",x"cf"),
  1201 => (x"b2",x"73",x"4a",x"72"),
  1202 => (x"c8",x"4b",x"66",x"cc"),
  1203 => (x"f0",x"ff",x"c0",x"33"),
  1204 => (x"72",x"9b",x"c0",x"c0"),
  1205 => (x"cc",x"b2",x"73",x"4a"),
  1206 => (x"33",x"d8",x"4b",x"66"),
  1207 => (x"c0",x"c0",x"c0",x"ff"),
  1208 => (x"4a",x"72",x"9b",x"c0"),
  1209 => (x"48",x"72",x"b2",x"73"),
  1210 => (x"4a",x"26",x"4b",x"26"),
  1211 => (x"5e",x"0e",x"4f",x"26"),
  1212 => (x"cc",x"0e",x"5b",x"5a"),
  1213 => (x"2b",x"c8",x"4b",x"66"),
  1214 => (x"cc",x"9b",x"ff",x"c3"),
  1215 => (x"32",x"c8",x"4a",x"66"),
  1216 => (x"9a",x"c0",x"fc",x"cf"),
  1217 => (x"9b",x"ff",x"ff",x"cf"),
  1218 => (x"b2",x"73",x"4a",x"72"),
  1219 => (x"9a",x"ff",x"ff",x"cf"),
  1220 => (x"4b",x"26",x"48",x"72"),
  1221 => (x"4f",x"26",x"4a",x"26"),
  1222 => (x"5b",x"5a",x"5e",x"0e"),
  1223 => (x"4a",x"66",x"cc",x"0e"),
  1224 => (x"ff",x"cf",x"2a",x"d0"),
  1225 => (x"66",x"cc",x"9a",x"ff"),
  1226 => (x"f0",x"33",x"d0",x"4b"),
  1227 => (x"72",x"9b",x"c0",x"c0"),
  1228 => (x"72",x"b2",x"73",x"4a"),
  1229 => (x"26",x"4b",x"26",x"48"),
  1230 => (x"1e",x"4f",x"26",x"4a"),
  1231 => (x"c0",x"d0",x"1e",x"72"),
  1232 => (x"4a",x"c0",x"c0",x"c0"),
  1233 => (x"fd",x"ff",x"0f",x"72"),
  1234 => (x"26",x"4a",x"26",x"87"),
  1235 => (x"1e",x"72",x"1e",x"4f"),
  1236 => (x"c3",x"4a",x"66",x"cc"),
  1237 => (x"f7",x"c0",x"9a",x"df"),
  1238 => (x"aa",x"b7",x"c0",x"8a"),
  1239 => (x"87",x"c3",x"c0",x"03"),
  1240 => (x"c8",x"82",x"e7",x"c0"),
  1241 => (x"30",x"c4",x"48",x"66"),
  1242 => (x"c8",x"58",x"a6",x"cc"),
  1243 => (x"b0",x"72",x"48",x"66"),
  1244 => (x"c8",x"58",x"a6",x"cc"),
  1245 => (x"4a",x"26",x"48",x"66"),
  1246 => (x"5e",x"0e",x"4f",x"26"),
  1247 => (x"5d",x"5c",x"5b",x"5a"),
  1248 => (x"c0",x"c0",x"d0",x"0e"),
  1249 => (x"27",x"4d",x"c0",x"c0"),
  1250 => (x"00",x"00",x"1b",x"bc"),
  1251 => (x"80",x"c1",x"48",x"bf"),
  1252 => (x"00",x"1b",x"c0",x"27"),
  1253 => (x"d4",x"97",x"58",x"00"),
  1254 => (x"c0",x"c1",x"4a",x"66"),
  1255 => (x"92",x"c0",x"c0",x"c0"),
  1256 => (x"92",x"b7",x"c0",x"c4"),
  1257 => (x"b7",x"d3",x"c1",x"4a"),
  1258 => (x"e9",x"c0",x"05",x"aa"),
  1259 => (x"1b",x"bc",x"27",x"87"),
  1260 => (x"c0",x"49",x"00",x"00"),
  1261 => (x"1b",x"c0",x"27",x"79"),
  1262 => (x"c0",x"49",x"00",x"00"),
  1263 => (x"1b",x"c8",x"27",x"79"),
  1264 => (x"c0",x"49",x"00",x"00"),
  1265 => (x"1b",x"cc",x"27",x"79"),
  1266 => (x"c0",x"49",x"00",x"00"),
  1267 => (x"49",x"c0",x"ff",x"79"),
  1268 => (x"ca",x"79",x"d3",x"c1"),
  1269 => (x"bc",x"27",x"87",x"cb"),
  1270 => (x"bf",x"00",x"00",x"1b"),
  1271 => (x"a9",x"b7",x"c1",x"49"),
  1272 => (x"87",x"db",x"c1",x"05"),
  1273 => (x"c1",x"49",x"c0",x"ff"),
  1274 => (x"d4",x"97",x"79",x"f4"),
  1275 => (x"c0",x"c1",x"4a",x"66"),
  1276 => (x"92",x"c0",x"c0",x"c0"),
  1277 => (x"92",x"b7",x"c0",x"c4"),
  1278 => (x"27",x"1e",x"72",x"4a"),
  1279 => (x"00",x"00",x"1b",x"cc"),
  1280 => (x"4d",x"27",x"1e",x"bf"),
  1281 => (x"0f",x"00",x"00",x"13"),
  1282 => (x"d0",x"27",x"86",x"c8"),
  1283 => (x"58",x"00",x"00",x"1b"),
  1284 => (x"00",x"1b",x"cc",x"27"),
  1285 => (x"c3",x"4c",x"bf",x"00"),
  1286 => (x"c0",x"06",x"ac",x"b7"),
  1287 => (x"48",x"ca",x"87",x"c6"),
  1288 => (x"4c",x"70",x"88",x"74"),
  1289 => (x"82",x"c1",x"4a",x"74"),
  1290 => (x"30",x"c1",x"48",x"72"),
  1291 => (x"00",x"1b",x"c8",x"27"),
  1292 => (x"48",x"74",x"58",x"00"),
  1293 => (x"ff",x"80",x"f0",x"c0"),
  1294 => (x"79",x"70",x"49",x"c0"),
  1295 => (x"27",x"87",x"e2",x"c8"),
  1296 => (x"00",x"00",x"1b",x"cc"),
  1297 => (x"b7",x"c9",x"49",x"bf"),
  1298 => (x"d4",x"c8",x"01",x"a9"),
  1299 => (x"1b",x"cc",x"27",x"87"),
  1300 => (x"49",x"bf",x"00",x"00"),
  1301 => (x"06",x"a9",x"b7",x"c0"),
  1302 => (x"27",x"87",x"c6",x"c8"),
  1303 => (x"00",x"00",x"1b",x"cc"),
  1304 => (x"f0",x"c0",x"48",x"bf"),
  1305 => (x"49",x"c0",x"ff",x"80"),
  1306 => (x"bc",x"27",x"79",x"70"),
  1307 => (x"bf",x"00",x"00",x"1b"),
  1308 => (x"a9",x"b7",x"c3",x"49"),
  1309 => (x"87",x"e9",x"c0",x"01"),
  1310 => (x"4a",x"66",x"d4",x"97"),
  1311 => (x"c0",x"c0",x"c0",x"c1"),
  1312 => (x"c0",x"c4",x"92",x"c0"),
  1313 => (x"72",x"4a",x"92",x"b7"),
  1314 => (x"1b",x"c8",x"27",x"1e"),
  1315 => (x"1e",x"bf",x"00",x"00"),
  1316 => (x"00",x"13",x"4d",x"27"),
  1317 => (x"86",x"c8",x"0f",x"00"),
  1318 => (x"00",x"1b",x"cc",x"27"),
  1319 => (x"c0",x"c7",x"58",x"00"),
  1320 => (x"1b",x"c4",x"27",x"87"),
  1321 => (x"4a",x"bf",x"00",x"00"),
  1322 => (x"bc",x"27",x"82",x"c3"),
  1323 => (x"bf",x"00",x"00",x"1b"),
  1324 => (x"a9",x"b7",x"72",x"49"),
  1325 => (x"87",x"f1",x"c0",x"01"),
  1326 => (x"4a",x"66",x"d4",x"97"),
  1327 => (x"c0",x"c0",x"c0",x"c1"),
  1328 => (x"c0",x"c4",x"92",x"c0"),
  1329 => (x"72",x"4a",x"92",x"b7"),
  1330 => (x"1b",x"c0",x"27",x"1e"),
  1331 => (x"1e",x"bf",x"00",x"00"),
  1332 => (x"00",x"13",x"4d",x"27"),
  1333 => (x"86",x"c8",x"0f",x"00"),
  1334 => (x"00",x"1b",x"c4",x"27"),
  1335 => (x"d0",x"27",x"58",x"00"),
  1336 => (x"49",x"00",x"00",x"1b"),
  1337 => (x"f8",x"c5",x"79",x"c1"),
  1338 => (x"1b",x"cc",x"27",x"87"),
  1339 => (x"49",x"bf",x"00",x"00"),
  1340 => (x"06",x"a9",x"b7",x"c0"),
  1341 => (x"27",x"87",x"d0",x"c3"),
  1342 => (x"00",x"00",x"1b",x"cc"),
  1343 => (x"b7",x"c3",x"49",x"bf"),
  1344 => (x"c2",x"c3",x"01",x"a9"),
  1345 => (x"1b",x"c8",x"27",x"87"),
  1346 => (x"4a",x"bf",x"00",x"00"),
  1347 => (x"82",x"c1",x"32",x"c1"),
  1348 => (x"00",x"1b",x"bc",x"27"),
  1349 => (x"72",x"49",x"bf",x"00"),
  1350 => (x"c2",x"01",x"a9",x"b7"),
  1351 => (x"d4",x"97",x"87",x"c2"),
  1352 => (x"c0",x"c1",x"4a",x"66"),
  1353 => (x"92",x"c0",x"c0",x"c0"),
  1354 => (x"92",x"b7",x"c0",x"c4"),
  1355 => (x"27",x"1e",x"72",x"4a"),
  1356 => (x"00",x"00",x"1b",x"d4"),
  1357 => (x"4d",x"27",x"1e",x"bf"),
  1358 => (x"0f",x"00",x"00",x"13"),
  1359 => (x"d8",x"27",x"86",x"c8"),
  1360 => (x"58",x"00",x"00",x"1b"),
  1361 => (x"00",x"1b",x"d0",x"27"),
  1362 => (x"c1",x"4a",x"bf",x"00"),
  1363 => (x"1b",x"d0",x"27",x"8a"),
  1364 => (x"72",x"49",x"00",x"00"),
  1365 => (x"aa",x"b7",x"c0",x"79"),
  1366 => (x"87",x"c5",x"c4",x"03"),
  1367 => (x"00",x"1b",x"c0",x"27"),
  1368 => (x"27",x"4a",x"bf",x"00"),
  1369 => (x"00",x"00",x"1b",x"d4"),
  1370 => (x"27",x"52",x"bf",x"97"),
  1371 => (x"00",x"00",x"1b",x"c0"),
  1372 => (x"82",x"c1",x"4a",x"bf"),
  1373 => (x"00",x"1b",x"c0",x"27"),
  1374 => (x"79",x"72",x"49",x"00"),
  1375 => (x"00",x"1b",x"d8",x"27"),
  1376 => (x"aa",x"b7",x"bf",x"00"),
  1377 => (x"87",x"cd",x"c0",x"06"),
  1378 => (x"00",x"1b",x"d8",x"27"),
  1379 => (x"c0",x"27",x"49",x"00"),
  1380 => (x"bf",x"00",x"00",x"1b"),
  1381 => (x"1b",x"d0",x"27",x"79"),
  1382 => (x"c1",x"49",x"00",x"00"),
  1383 => (x"87",x"c1",x"c3",x"79"),
  1384 => (x"00",x"1b",x"d0",x"27"),
  1385 => (x"c2",x"05",x"bf",x"00"),
  1386 => (x"d4",x"27",x"87",x"f7"),
  1387 => (x"bf",x"00",x"00",x"1b"),
  1388 => (x"27",x"32",x"c4",x"4a"),
  1389 => (x"00",x"00",x"1b",x"d4"),
  1390 => (x"27",x"79",x"72",x"49"),
  1391 => (x"00",x"00",x"1b",x"c0"),
  1392 => (x"51",x"72",x"49",x"bf"),
  1393 => (x"27",x"87",x"da",x"c2"),
  1394 => (x"00",x"00",x"1b",x"cc"),
  1395 => (x"b7",x"c7",x"49",x"bf"),
  1396 => (x"fd",x"c1",x"04",x"a9"),
  1397 => (x"fe",x"4b",x"c0",x"87"),
  1398 => (x"79",x"c1",x"49",x"f4"),
  1399 => (x"00",x"1b",x"d8",x"27"),
  1400 => (x"75",x"1e",x"bf",x"00"),
  1401 => (x"19",x"2b",x"27",x"1e"),
  1402 => (x"27",x"1e",x"00",x"00"),
  1403 => (x"00",x"00",x"00",x"9a"),
  1404 => (x"27",x"86",x"cc",x"0f"),
  1405 => (x"00",x"00",x"1b",x"c0"),
  1406 => (x"27",x"79",x"75",x"49"),
  1407 => (x"00",x"00",x"1b",x"c0"),
  1408 => (x"d8",x"27",x"49",x"bf"),
  1409 => (x"bf",x"00",x"00",x"1b"),
  1410 => (x"c0",x"03",x"a9",x"b7"),
  1411 => (x"c0",x"27",x"87",x"e5"),
  1412 => (x"bf",x"00",x"00",x"1b"),
  1413 => (x"c0",x"27",x"83",x"bf"),
  1414 => (x"bf",x"00",x"00",x"1b"),
  1415 => (x"27",x"82",x"c4",x"4a"),
  1416 => (x"00",x"00",x"1b",x"c0"),
  1417 => (x"27",x"79",x"72",x"49"),
  1418 => (x"00",x"00",x"1b",x"d8"),
  1419 => (x"04",x"aa",x"b7",x"bf"),
  1420 => (x"73",x"87",x"db",x"ff"),
  1421 => (x"19",x"4a",x"27",x"1e"),
  1422 => (x"27",x"1e",x"00",x"00"),
  1423 => (x"00",x"00",x"00",x"9a"),
  1424 => (x"ff",x"86",x"c8",x"0f"),
  1425 => (x"c2",x"c1",x"49",x"c0"),
  1426 => (x"13",x"3b",x"27",x"79"),
  1427 => (x"c0",x"0f",x"00",x"00"),
  1428 => (x"cc",x"27",x"87",x"cf"),
  1429 => (x"bf",x"00",x"00",x"1b"),
  1430 => (x"80",x"f0",x"c0",x"48"),
  1431 => (x"70",x"49",x"c0",x"ff"),
  1432 => (x"26",x"4d",x"26",x"79"),
  1433 => (x"26",x"4b",x"26",x"4c"),
  1434 => (x"0e",x"4f",x"26",x"4a"),
  1435 => (x"5c",x"5b",x"5a",x"5e"),
  1436 => (x"27",x"1e",x"0e",x"5d"),
  1437 => (x"00",x"00",x"17",x"7e"),
  1438 => (x"00",x"61",x"27",x"1e"),
  1439 => (x"c4",x"0f",x"00",x"00"),
  1440 => (x"04",x"ff",x"27",x"86"),
  1441 => (x"70",x"0f",x"00",x"00"),
  1442 => (x"02",x"9a",x"72",x"4a"),
  1443 => (x"27",x"87",x"d3",x"c0"),
  1444 => (x"00",x"00",x"0a",x"c0"),
  1445 => (x"72",x"4a",x"70",x"0f"),
  1446 => (x"c5",x"c0",x"02",x"9a"),
  1447 => (x"c0",x"4a",x"c1",x"87"),
  1448 => (x"4a",x"c0",x"87",x"c2"),
  1449 => (x"79",x"72",x"49",x"76"),
  1450 => (x"00",x"17",x"94",x"27"),
  1451 => (x"61",x"27",x"1e",x"00"),
  1452 => (x"0f",x"00",x"00",x"00"),
  1453 => (x"d8",x"27",x"86",x"c4"),
  1454 => (x"49",x"00",x"00",x"1b"),
  1455 => (x"ee",x"c0",x"79",x"c0"),
  1456 => (x"00",x"42",x"27",x"1e"),
  1457 => (x"c4",x"0f",x"00",x"00"),
  1458 => (x"c8",x"f4",x"c3",x"86"),
  1459 => (x"c0",x"ff",x"4b",x"ff"),
  1460 => (x"4a",x"74",x"4c",x"bf"),
  1461 => (x"72",x"9a",x"c0",x"c8"),
  1462 => (x"e1",x"c1",x"02",x"9a"),
  1463 => (x"c3",x"4d",x"74",x"87"),
  1464 => (x"b7",x"db",x"9d",x"ff"),
  1465 => (x"c6",x"c1",x"05",x"ad"),
  1466 => (x"c0",x"02",x"6e",x"87"),
  1467 => (x"c0",x"d0",x"87",x"f3"),
  1468 => (x"1e",x"c0",x"c0",x"c0"),
  1469 => (x"00",x"17",x"62",x"27"),
  1470 => (x"e2",x"27",x"1e",x"00"),
  1471 => (x"0f",x"00",x"00",x"11"),
  1472 => (x"4a",x"70",x"86",x"c8"),
  1473 => (x"c0",x"02",x"9a",x"72"),
  1474 => (x"56",x"27",x"87",x"d7"),
  1475 => (x"1e",x"00",x"00",x"17"),
  1476 => (x"00",x"00",x"61",x"27"),
  1477 => (x"86",x"c4",x"0f",x"00"),
  1478 => (x"00",x"13",x"3b",x"27"),
  1479 => (x"ce",x"c0",x"0f",x"00"),
  1480 => (x"17",x"6e",x"27",x"87"),
  1481 => (x"27",x"1e",x"00",x"00"),
  1482 => (x"00",x"00",x"00",x"61"),
  1483 => (x"75",x"86",x"c4",x"0f"),
  1484 => (x"13",x"7a",x"27",x"1e"),
  1485 => (x"c4",x"0f",x"00",x"00"),
  1486 => (x"c9",x"f4",x"c3",x"86"),
  1487 => (x"4a",x"73",x"4b",x"c0"),
  1488 => (x"9a",x"72",x"8b",x"c1"),
  1489 => (x"87",x"c6",x"fe",x"05"),
  1490 => (x"26",x"87",x"f3",x"fd"),
  1491 => (x"4c",x"26",x"4d",x"26"),
  1492 => (x"4a",x"26",x"4b",x"26"),
  1493 => (x"6f",x"42",x"4f",x"26"),
  1494 => (x"6e",x"69",x"74",x"6f"),
  1495 => (x"2e",x"2e",x"2e",x"67"),
  1496 => (x"4f",x"42",x"00",x"0a"),
  1497 => (x"33",x"38",x"54",x"4f"),
  1498 => (x"49",x"42",x"20",x"32"),
  1499 => (x"44",x"53",x"00",x"4e"),
  1500 => (x"6f",x"6f",x"62",x"20"),
  1501 => (x"61",x"66",x"20",x"74"),
  1502 => (x"64",x"65",x"6c",x"69"),
  1503 => (x"6e",x"49",x"00",x"0a"),
  1504 => (x"61",x"69",x"74",x"69"),
  1505 => (x"69",x"7a",x"69",x"6c"),
  1506 => (x"53",x"20",x"67",x"6e"),
  1507 => (x"61",x"63",x"20",x"44"),
  1508 => (x"00",x"0a",x"64",x"72"),
  1509 => (x"33",x"32",x"53",x"52"),
  1510 => (x"6f",x"62",x"20",x"32"),
  1511 => (x"2d",x"20",x"74",x"6f"),
  1512 => (x"65",x"72",x"70",x"20"),
  1513 => (x"45",x"20",x"73",x"73"),
  1514 => (x"74",x"20",x"43",x"53"),
  1515 => (x"6f",x"62",x"20",x"6f"),
  1516 => (x"66",x"20",x"74",x"6f"),
  1517 => (x"20",x"6d",x"6f",x"72"),
  1518 => (x"00",x"2e",x"44",x"53"),
  1519 => (x"00",x"44",x"4d",x"43"),
  1520 => (x"64",x"61",x"65",x"52"),
  1521 => (x"20",x"66",x"6f",x"20"),
  1522 => (x"20",x"52",x"42",x"4d"),
  1523 => (x"6c",x"69",x"61",x"66"),
  1524 => (x"00",x"0a",x"64",x"65"),
  1525 => (x"70",x"20",x"6f",x"4e"),
  1526 => (x"69",x"74",x"72",x"61"),
  1527 => (x"6e",x"6f",x"69",x"74"),
  1528 => (x"67",x"69",x"73",x"20"),
  1529 => (x"75",x"74",x"61",x"6e"),
  1530 => (x"66",x"20",x"65",x"72"),
  1531 => (x"64",x"6e",x"75",x"6f"),
  1532 => (x"42",x"4d",x"00",x"0a"),
  1533 => (x"7a",x"69",x"73",x"52"),
  1534 => (x"25",x"20",x"3a",x"65"),
  1535 => (x"70",x"20",x"2c",x"64"),
  1536 => (x"69",x"74",x"72",x"61"),
  1537 => (x"6e",x"6f",x"69",x"74"),
  1538 => (x"65",x"7a",x"69",x"73"),
  1539 => (x"64",x"25",x"20",x"3a"),
  1540 => (x"66",x"6f",x"20",x"2c"),
  1541 => (x"74",x"65",x"73",x"66"),
  1542 => (x"20",x"66",x"6f",x"20"),
  1543 => (x"3a",x"67",x"69",x"73"),
  1544 => (x"2c",x"64",x"25",x"20"),
  1545 => (x"67",x"69",x"73",x"20"),
  1546 => (x"25",x"78",x"30",x"20"),
  1547 => (x"52",x"00",x"0a",x"78"),
  1548 => (x"69",x"64",x"61",x"65"),
  1549 => (x"62",x"20",x"67",x"6e"),
  1550 => (x"20",x"74",x"6f",x"6f"),
  1551 => (x"74",x"63",x"65",x"73"),
  1552 => (x"25",x"20",x"72",x"6f"),
  1553 => (x"52",x"00",x"0a",x"64"),
  1554 => (x"20",x"64",x"61",x"65"),
  1555 => (x"74",x"6f",x"6f",x"62"),
  1556 => (x"63",x"65",x"73",x"20"),
  1557 => (x"20",x"72",x"6f",x"74"),
  1558 => (x"6d",x"6f",x"72",x"66"),
  1559 => (x"72",x"69",x"66",x"20"),
  1560 => (x"70",x"20",x"74",x"73"),
  1561 => (x"69",x"74",x"72",x"61"),
  1562 => (x"6e",x"6f",x"69",x"74"),
  1563 => (x"6e",x"55",x"00",x"0a"),
  1564 => (x"70",x"70",x"75",x"73"),
  1565 => (x"65",x"74",x"72",x"6f"),
  1566 => (x"61",x"70",x"20",x"64"),
  1567 => (x"74",x"69",x"74",x"72"),
  1568 => (x"20",x"6e",x"6f",x"69"),
  1569 => (x"65",x"70",x"79",x"74"),
  1570 => (x"46",x"00",x"0d",x"21"),
  1571 => (x"32",x"33",x"54",x"41"),
  1572 => (x"00",x"20",x"20",x"20"),
  1573 => (x"64",x"61",x"65",x"52"),
  1574 => (x"20",x"67",x"6e",x"69"),
  1575 => (x"0a",x"52",x"42",x"4d"),
  1576 => (x"52",x"42",x"4d",x"00"),
  1577 => (x"63",x"75",x"73",x"20"),
  1578 => (x"73",x"73",x"65",x"63"),
  1579 => (x"6c",x"6c",x"75",x"66"),
  1580 => (x"65",x"72",x"20",x"79"),
  1581 => (x"00",x"0a",x"64",x"61"),
  1582 => (x"31",x"54",x"41",x"46"),
  1583 => (x"20",x"20",x"20",x"36"),
  1584 => (x"54",x"41",x"46",x"00"),
  1585 => (x"20",x"20",x"32",x"33"),
  1586 => (x"61",x"50",x"00",x"20"),
  1587 => (x"74",x"69",x"74",x"72"),
  1588 => (x"63",x"6e",x"6f",x"69"),
  1589 => (x"74",x"6e",x"75",x"6f"),
  1590 => (x"0a",x"64",x"25",x"20"),
  1591 => (x"6e",x"75",x"48",x"00"),
  1592 => (x"67",x"6e",x"69",x"74"),
  1593 => (x"72",x"6f",x"66",x"20"),
  1594 => (x"6c",x"69",x"66",x"20"),
  1595 => (x"73",x"79",x"73",x"65"),
  1596 => (x"0a",x"6d",x"65",x"74"),
  1597 => (x"54",x"41",x"46",x"00"),
  1598 => (x"20",x"20",x"32",x"33"),
  1599 => (x"41",x"46",x"00",x"20"),
  1600 => (x"20",x"36",x"31",x"54"),
  1601 => (x"43",x"00",x"20",x"20"),
  1602 => (x"74",x"73",x"75",x"6c"),
  1603 => (x"73",x"20",x"72",x"65"),
  1604 => (x"3a",x"65",x"7a",x"69"),
  1605 => (x"2c",x"64",x"25",x"20"),
  1606 => (x"75",x"6c",x"43",x"20"),
  1607 => (x"72",x"65",x"74",x"73"),
  1608 => (x"73",x"61",x"6d",x"20"),
  1609 => (x"25",x"20",x"2c",x"6b"),
  1610 => (x"43",x"00",x"0a",x"64"),
  1611 => (x"6b",x"63",x"65",x"68"),
  1612 => (x"6d",x"6d",x"75",x"73"),
  1613 => (x"20",x"67",x"6e",x"69"),
  1614 => (x"6d",x"6f",x"72",x"66"),
  1615 => (x"20",x"64",x"25",x"20"),
  1616 => (x"25",x"20",x"6f",x"74"),
  1617 => (x"2e",x"2e",x"2e",x"64"),
  1618 => (x"64",x"25",x"00",x"20"),
  1619 => (x"64",x"25",x"00",x"0a"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
