
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"c9",x"01"),
     1 => (x"cf",x"03",x"87",x"cc"),
     2 => (x"87",x"fd",x"00",x"87"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"36",x"27",x"4f",x"00"),
     5 => (x"4f",x"00",x"00",x"00"),
     6 => (x"0e",x"1e",x"18",x"0e"),
     7 => (x"00",x"00",x"44",x"27"),
     8 => (x"48",x"26",x"0f",x"00"),
     9 => (x"08",x"26",x"80",x"ff"),
    10 => (x"c0",x"c0",x"c2",x"4f"),
    11 => (x"16",x"58",x"27",x"4e"),
    12 => (x"00",x"0f",x"00",x"00"),
    13 => (x"f0",x"c1",x"87",x"fd"),
    14 => (x"43",x"27",x"4e",x"c0"),
    15 => (x"0f",x"00",x"00",x"00"),
    16 => (x"4f",x"87",x"fd",x"00"),
    17 => (x"0e",x"1e",x"18",x"0e"),
    18 => (x"80",x"ff",x"48",x"26"),
    19 => (x"1e",x"4f",x"08",x"26"),
    20 => (x"ff",x"1e",x"1e",x"72"),
    21 => (x"48",x"6a",x"4a",x"c0"),
    22 => (x"c4",x"98",x"c0",x"c4"),
    23 => (x"02",x"6e",x"58",x"a6"),
    24 => (x"cc",x"87",x"f3",x"ff"),
    25 => (x"66",x"cc",x"7a",x"66"),
    26 => (x"4a",x"26",x"26",x"48"),
    27 => (x"5e",x"0e",x"4f",x"26"),
    28 => (x"5d",x"5c",x"5b",x"5a"),
    29 => (x"4b",x"66",x"d4",x"0e"),
    30 => (x"4c",x"13",x"4d",x"c0"),
    31 => (x"c0",x"02",x"9c",x"74"),
    32 => (x"4a",x"74",x"87",x"d6"),
    33 => (x"4f",x"27",x"1e",x"72"),
    34 => (x"0f",x"00",x"00",x"00"),
    35 => (x"85",x"c1",x"86",x"c4"),
    36 => (x"9c",x"74",x"4c",x"13"),
    37 => (x"87",x"ea",x"ff",x"05"),
    38 => (x"4d",x"26",x"48",x"75"),
    39 => (x"4b",x"26",x"4c",x"26"),
    40 => (x"4f",x"26",x"4a",x"26"),
    41 => (x"5b",x"5a",x"5e",x"0e"),
    42 => (x"1e",x"0e",x"5d",x"5c"),
    43 => (x"27",x"4d",x"66",x"d8"),
    44 => (x"00",x"00",x"1a",x"48"),
    45 => (x"27",x"49",x"76",x"4b"),
    46 => (x"00",x"00",x"18",x"b4"),
    47 => (x"c0",x"4c",x"c0",x"79"),
    48 => (x"c0",x"03",x"ad",x"b7"),
    49 => (x"ed",x"c0",x"87",x"cd"),
    50 => (x"00",x"4f",x"27",x"1e"),
    51 => (x"c4",x"0f",x"00",x"00"),
    52 => (x"75",x"8d",x"0d",x"86"),
    53 => (x"c6",x"c0",x"05",x"9d"),
    54 => (x"53",x"f0",x"c0",x"87"),
    55 => (x"75",x"87",x"f6",x"c0"),
    56 => (x"f0",x"c0",x"02",x"9d"),
    57 => (x"72",x"49",x"75",x"87"),
    58 => (x"66",x"e4",x"c0",x"1e"),
    59 => (x"18",x"6a",x"27",x"4a"),
    60 => (x"26",x"0f",x"00",x"00"),
    61 => (x"72",x"4a",x"71",x"4a"),
    62 => (x"12",x"82",x"6e",x"4a"),
    63 => (x"72",x"49",x"75",x"53"),
    64 => (x"66",x"e4",x"c0",x"1e"),
    65 => (x"18",x"6a",x"27",x"4a"),
    66 => (x"26",x"0f",x"00",x"00"),
    67 => (x"75",x"4d",x"70",x"4a"),
    68 => (x"d0",x"ff",x"05",x"9d"),
    69 => (x"1a",x"48",x"27",x"87"),
    70 => (x"ab",x"b7",x"00",x"00"),
    71 => (x"87",x"de",x"c0",x"02"),
    72 => (x"66",x"dc",x"8b",x"c1"),
    73 => (x"51",x"6b",x"97",x"49"),
    74 => (x"c1",x"48",x"66",x"dc"),
    75 => (x"a6",x"e0",x"c0",x"80"),
    76 => (x"27",x"84",x"c1",x"58"),
    77 => (x"00",x"00",x"1a",x"48"),
    78 => (x"ff",x"05",x"ab",x"b7"),
    79 => (x"66",x"dc",x"87",x"e2"),
    80 => (x"74",x"51",x"c0",x"49"),
    81 => (x"4d",x"26",x"26",x"48"),
    82 => (x"4b",x"26",x"4c",x"26"),
    83 => (x"4f",x"26",x"4a",x"26"),
    84 => (x"5b",x"5a",x"5e",x"0e"),
    85 => (x"1e",x"0e",x"5d",x"5c"),
    86 => (x"49",x"76",x"4c",x"c0"),
    87 => (x"a6",x"dc",x"79",x"c0"),
    88 => (x"4a",x"66",x"d8",x"4b"),
    89 => (x"c1",x"48",x"66",x"d8"),
    90 => (x"58",x"a6",x"dc",x"80"),
    91 => (x"35",x"d8",x"4d",x"12"),
    92 => (x"9d",x"75",x"2d",x"b7"),
    93 => (x"87",x"cb",x"c4",x"02"),
    94 => (x"d7",x"c3",x"02",x"6e"),
    95 => (x"c0",x"49",x"76",x"87"),
    96 => (x"c1",x"4a",x"75",x"79"),
    97 => (x"c2",x"02",x"ad",x"e3"),
    98 => (x"e4",x"c1",x"87",x"dd"),
    99 => (x"d8",x"c0",x"02",x"aa"),
   100 => (x"aa",x"ec",x"c1",x"87"),
   101 => (x"87",x"c8",x"c2",x"02"),
   102 => (x"02",x"aa",x"f3",x"c1"),
   103 => (x"c1",x"87",x"e8",x"c1"),
   104 => (x"c0",x"02",x"aa",x"f8"),
   105 => (x"d3",x"c2",x"87",x"f2"),
   106 => (x"27",x"1e",x"ca",x"87"),
   107 => (x"00",x"00",x"1a",x"98"),
   108 => (x"73",x"83",x"c4",x"1e"),
   109 => (x"6a",x"8a",x"c4",x"4a"),
   110 => (x"00",x"a4",x"27",x"1e"),
   111 => (x"cc",x"0f",x"00",x"00"),
   112 => (x"74",x"4a",x"70",x"86"),
   113 => (x"27",x"84",x"72",x"4c"),
   114 => (x"00",x"00",x"1a",x"98"),
   115 => (x"00",x"6e",x"27",x"1e"),
   116 => (x"c4",x"0f",x"00",x"00"),
   117 => (x"87",x"d4",x"c2",x"86"),
   118 => (x"98",x"27",x"1e",x"d0"),
   119 => (x"1e",x"00",x"00",x"1a"),
   120 => (x"4a",x"73",x"83",x"c4"),
   121 => (x"1e",x"6a",x"8a",x"c4"),
   122 => (x"00",x"00",x"a4",x"27"),
   123 => (x"86",x"cc",x"0f",x"00"),
   124 => (x"4c",x"74",x"4a",x"70"),
   125 => (x"98",x"27",x"84",x"72"),
   126 => (x"1e",x"00",x"00",x"1a"),
   127 => (x"00",x"00",x"6e",x"27"),
   128 => (x"86",x"c4",x"0f",x"00"),
   129 => (x"c4",x"87",x"e5",x"c1"),
   130 => (x"c4",x"4a",x"73",x"83"),
   131 => (x"27",x"1e",x"6a",x"8a"),
   132 => (x"00",x"00",x"00",x"6e"),
   133 => (x"70",x"86",x"c4",x"0f"),
   134 => (x"72",x"4c",x"74",x"4a"),
   135 => (x"87",x"cc",x"c1",x"84"),
   136 => (x"79",x"c1",x"49",x"76"),
   137 => (x"c4",x"87",x"c5",x"c1"),
   138 => (x"c4",x"4a",x"73",x"83"),
   139 => (x"27",x"1e",x"6a",x"8a"),
   140 => (x"00",x"00",x"00",x"4f"),
   141 => (x"c1",x"86",x"c4",x"0f"),
   142 => (x"87",x"f0",x"c0",x"84"),
   143 => (x"27",x"1e",x"e5",x"c0"),
   144 => (x"00",x"00",x"00",x"4f"),
   145 => (x"75",x"86",x"c4",x"0f"),
   146 => (x"00",x"4f",x"27",x"1e"),
   147 => (x"c4",x"0f",x"00",x"00"),
   148 => (x"87",x"d8",x"c0",x"86"),
   149 => (x"05",x"ad",x"e5",x"c0"),
   150 => (x"76",x"87",x"c7",x"c0"),
   151 => (x"c0",x"79",x"c1",x"49"),
   152 => (x"1e",x"75",x"87",x"ca"),
   153 => (x"00",x"00",x"4f",x"27"),
   154 => (x"86",x"c4",x"0f",x"00"),
   155 => (x"d8",x"4a",x"66",x"d8"),
   156 => (x"80",x"c1",x"48",x"66"),
   157 => (x"12",x"58",x"a6",x"dc"),
   158 => (x"b7",x"35",x"d8",x"4d"),
   159 => (x"05",x"9d",x"75",x"2d"),
   160 => (x"74",x"87",x"f5",x"fb"),
   161 => (x"4d",x"26",x"26",x"48"),
   162 => (x"4b",x"26",x"4c",x"26"),
   163 => (x"4f",x"26",x"4a",x"26"),
   164 => (x"00",x"00",x"00",x"00"),
   165 => (x"ff",x"1e",x"75",x"1e"),
   166 => (x"ff",x"c3",x"4d",x"d4"),
   167 => (x"48",x"6d",x"7d",x"49"),
   168 => (x"7d",x"71",x"38",x"c8"),
   169 => (x"38",x"c8",x"b0",x"6d"),
   170 => (x"b0",x"6d",x"7d",x"71"),
   171 => (x"7d",x"71",x"38",x"c8"),
   172 => (x"38",x"c8",x"b0",x"6d"),
   173 => (x"4f",x"26",x"4d",x"26"),
   174 => (x"ff",x"1e",x"75",x"1e"),
   175 => (x"ff",x"c3",x"4d",x"d4"),
   176 => (x"48",x"6d",x"7d",x"49"),
   177 => (x"7d",x"71",x"30",x"c8"),
   178 => (x"30",x"c8",x"b0",x"6d"),
   179 => (x"b0",x"6d",x"7d",x"71"),
   180 => (x"7d",x"71",x"30",x"c8"),
   181 => (x"4d",x"26",x"b0",x"6d"),
   182 => (x"75",x"1e",x"4f",x"26"),
   183 => (x"4d",x"d4",x"ff",x"1e"),
   184 => (x"c8",x"49",x"66",x"cc"),
   185 => (x"fe",x"7d",x"48",x"66"),
   186 => (x"c9",x"02",x"67",x"e6"),
   187 => (x"39",x"d8",x"07",x"31"),
   188 => (x"39",x"09",x"7d",x"09"),
   189 => (x"39",x"09",x"7d",x"09"),
   190 => (x"39",x"09",x"7d",x"09"),
   191 => (x"38",x"d0",x"7d",x"09"),
   192 => (x"f1",x"c9",x"7d",x"70"),
   193 => (x"ff",x"c3",x"49",x"c0"),
   194 => (x"a8",x"08",x"6d",x"48"),
   195 => (x"08",x"87",x"c7",x"05"),
   196 => (x"05",x"89",x"c1",x"7d"),
   197 => (x"4d",x"26",x"87",x"f3"),
   198 => (x"72",x"1e",x"4f",x"26"),
   199 => (x"ff",x"4a",x"c0",x"1e"),
   200 => (x"ff",x"c3",x"49",x"d4"),
   201 => (x"c3",x"82",x"c1",x"79"),
   202 => (x"04",x"aa",x"b7",x"c8"),
   203 => (x"26",x"87",x"f0",x"ff"),
   204 => (x"0e",x"4f",x"26",x"4a"),
   205 => (x"5c",x"5b",x"5a",x"5e"),
   206 => (x"ff",x"c0",x"0e",x"5d"),
   207 => (x"4d",x"f7",x"c1",x"f0"),
   208 => (x"c0",x"c0",x"c0",x"c1"),
   209 => (x"27",x"4b",x"c0",x"c0"),
   210 => (x"00",x"00",x"03",x"1a"),
   211 => (x"df",x"f8",x"c4",x"0f"),
   212 => (x"75",x"1e",x"c0",x"4c"),
   213 => (x"02",x"da",x"27",x"1e"),
   214 => (x"c8",x"0f",x"00",x"00"),
   215 => (x"c1",x"4a",x"70",x"86"),
   216 => (x"c0",x"05",x"aa",x"b7"),
   217 => (x"d4",x"ff",x"87",x"ef"),
   218 => (x"79",x"ff",x"c3",x"49"),
   219 => (x"e1",x"c0",x"1e",x"73"),
   220 => (x"1e",x"e9",x"c1",x"f0"),
   221 => (x"00",x"02",x"da",x"27"),
   222 => (x"86",x"c8",x"0f",x"00"),
   223 => (x"9a",x"72",x"4a",x"70"),
   224 => (x"87",x"cb",x"c0",x"05"),
   225 => (x"c3",x"49",x"d4",x"ff"),
   226 => (x"48",x"c1",x"79",x"ff"),
   227 => (x"27",x"87",x"d0",x"c0"),
   228 => (x"00",x"00",x"03",x"1a"),
   229 => (x"74",x"8c",x"c1",x"0f"),
   230 => (x"f4",x"fe",x"05",x"9c"),
   231 => (x"26",x"48",x"c0",x"87"),
   232 => (x"26",x"4c",x"26",x"4d"),
   233 => (x"26",x"4a",x"26",x"4b"),
   234 => (x"5a",x"5e",x"0e",x"4f"),
   235 => (x"c0",x"0e",x"5c",x"5b"),
   236 => (x"c1",x"c1",x"f0",x"ff"),
   237 => (x"49",x"d4",x"ff",x"4c"),
   238 => (x"27",x"79",x"ff",x"c3"),
   239 => (x"00",x"00",x"18",x"c5"),
   240 => (x"00",x"6e",x"27",x"1e"),
   241 => (x"c4",x"0f",x"00",x"00"),
   242 => (x"c0",x"4b",x"d3",x"86"),
   243 => (x"27",x"1e",x"74",x"1e"),
   244 => (x"00",x"00",x"02",x"da"),
   245 => (x"70",x"86",x"c8",x"0f"),
   246 => (x"05",x"9a",x"72",x"4a"),
   247 => (x"ff",x"87",x"cb",x"c0"),
   248 => (x"ff",x"c3",x"49",x"d4"),
   249 => (x"c0",x"48",x"c1",x"79"),
   250 => (x"1a",x"27",x"87",x"d0"),
   251 => (x"0f",x"00",x"00",x"03"),
   252 => (x"9b",x"73",x"8b",x"c1"),
   253 => (x"87",x"d3",x"ff",x"05"),
   254 => (x"4c",x"26",x"48",x"c0"),
   255 => (x"4a",x"26",x"4b",x"26"),
   256 => (x"5e",x"0e",x"4f",x"26"),
   257 => (x"5d",x"5c",x"5b",x"5a"),
   258 => (x"ff",x"c3",x"1e",x"0e"),
   259 => (x"4c",x"d4",x"ff",x"4d"),
   260 => (x"00",x"03",x"1a",x"27"),
   261 => (x"ea",x"c6",x"0f",x"00"),
   262 => (x"f0",x"e1",x"c0",x"1e"),
   263 => (x"27",x"1e",x"c8",x"c1"),
   264 => (x"00",x"00",x"02",x"da"),
   265 => (x"70",x"86",x"c8",x"0f"),
   266 => (x"27",x"1e",x"72",x"4a"),
   267 => (x"00",x"00",x"05",x"61"),
   268 => (x"01",x"50",x"27",x"1e"),
   269 => (x"c8",x"0f",x"00",x"00"),
   270 => (x"aa",x"b7",x"c1",x"86"),
   271 => (x"87",x"cb",x"c0",x"02"),
   272 => (x"00",x"03",x"a9",x"27"),
   273 => (x"48",x"c0",x"0f",x"00"),
   274 => (x"27",x"87",x"c9",x"c3"),
   275 => (x"00",x"00",x"02",x"b8"),
   276 => (x"cf",x"4a",x"70",x"0f"),
   277 => (x"c6",x"9a",x"ff",x"ff"),
   278 => (x"02",x"aa",x"b7",x"ea"),
   279 => (x"27",x"87",x"cb",x"c0"),
   280 => (x"00",x"00",x"03",x"a9"),
   281 => (x"c2",x"48",x"c0",x"0f"),
   282 => (x"7c",x"75",x"87",x"ea"),
   283 => (x"f1",x"c0",x"49",x"76"),
   284 => (x"03",x"33",x"27",x"79"),
   285 => (x"70",x"0f",x"00",x"00"),
   286 => (x"02",x"9a",x"72",x"4a"),
   287 => (x"c0",x"87",x"eb",x"c1"),
   288 => (x"f0",x"ff",x"c0",x"1e"),
   289 => (x"27",x"1e",x"fa",x"c1"),
   290 => (x"00",x"00",x"02",x"da"),
   291 => (x"70",x"86",x"c8",x"0f"),
   292 => (x"05",x"9b",x"73",x"4b"),
   293 => (x"73",x"87",x"c3",x"c1"),
   294 => (x"05",x"1f",x"27",x"1e"),
   295 => (x"27",x"1e",x"00",x"00"),
   296 => (x"00",x"00",x"01",x"50"),
   297 => (x"75",x"86",x"c8",x"0f"),
   298 => (x"75",x"4b",x"6c",x"7c"),
   299 => (x"27",x"1e",x"73",x"9b"),
   300 => (x"00",x"00",x"05",x"2b"),
   301 => (x"01",x"50",x"27",x"1e"),
   302 => (x"c8",x"0f",x"00",x"00"),
   303 => (x"75",x"7c",x"75",x"86"),
   304 => (x"75",x"7c",x"75",x"7c"),
   305 => (x"c1",x"4a",x"73",x"7c"),
   306 => (x"9a",x"72",x"9a",x"c0"),
   307 => (x"87",x"c5",x"c0",x"02"),
   308 => (x"ff",x"c0",x"48",x"c1"),
   309 => (x"c0",x"48",x"c0",x"87"),
   310 => (x"1e",x"73",x"87",x"fa"),
   311 => (x"00",x"05",x"39",x"27"),
   312 => (x"50",x"27",x"1e",x"00"),
   313 => (x"0f",x"00",x"00",x"01"),
   314 => (x"49",x"6e",x"86",x"c8"),
   315 => (x"05",x"a9",x"b7",x"c2"),
   316 => (x"27",x"87",x"d3",x"c0"),
   317 => (x"00",x"00",x"05",x"45"),
   318 => (x"01",x"50",x"27",x"1e"),
   319 => (x"c4",x"0f",x"00",x"00"),
   320 => (x"c0",x"48",x"c0",x"86"),
   321 => (x"48",x"6e",x"87",x"ce"),
   322 => (x"a6",x"c4",x"88",x"c1"),
   323 => (x"fd",x"05",x"6e",x"58"),
   324 => (x"48",x"c0",x"87",x"df"),
   325 => (x"26",x"4d",x"26",x"26"),
   326 => (x"26",x"4b",x"26",x"4c"),
   327 => (x"43",x"4f",x"26",x"4a"),
   328 => (x"38",x"35",x"44",x"4d"),
   329 => (x"0a",x"64",x"25",x"20"),
   330 => (x"43",x"00",x"20",x"20"),
   331 => (x"38",x"35",x"44",x"4d"),
   332 => (x"25",x"20",x"32",x"5f"),
   333 => (x"20",x"20",x"0a",x"64"),
   334 => (x"44",x"4d",x"43",x"00"),
   335 => (x"25",x"20",x"38",x"35"),
   336 => (x"20",x"20",x"0a",x"64"),
   337 => (x"48",x"44",x"53",x"00"),
   338 => (x"6e",x"49",x"20",x"43"),
   339 => (x"61",x"69",x"74",x"69"),
   340 => (x"61",x"7a",x"69",x"6c"),
   341 => (x"6e",x"6f",x"69",x"74"),
   342 => (x"72",x"72",x"65",x"20"),
   343 => (x"0a",x"21",x"72",x"6f"),
   344 => (x"64",x"6d",x"63",x"00"),
   345 => (x"44",x"4d",x"43",x"5f"),
   346 => (x"65",x"72",x"20",x"38"),
   347 => (x"6e",x"6f",x"70",x"73"),
   348 => (x"20",x"3a",x"65",x"73"),
   349 => (x"00",x"0a",x"64",x"25"),
   350 => (x"5b",x"5a",x"5e",x"0e"),
   351 => (x"1e",x"0e",x"5d",x"5c"),
   352 => (x"c8",x"4c",x"d0",x"ff"),
   353 => (x"27",x"4b",x"c0",x"c0"),
   354 => (x"00",x"00",x"02",x"90"),
   355 => (x"27",x"79",x"c1",x"49"),
   356 => (x"00",x"00",x"06",x"95"),
   357 => (x"00",x"6e",x"27",x"1e"),
   358 => (x"c4",x"0f",x"00",x"00"),
   359 => (x"6c",x"4d",x"c7",x"86"),
   360 => (x"c4",x"98",x"73",x"48"),
   361 => (x"02",x"6e",x"58",x"a6"),
   362 => (x"6c",x"87",x"cc",x"c0"),
   363 => (x"c4",x"98",x"73",x"48"),
   364 => (x"05",x"6e",x"58",x"a6"),
   365 => (x"c0",x"87",x"f4",x"ff"),
   366 => (x"03",x"1a",x"27",x"7c"),
   367 => (x"6c",x"0f",x"00",x"00"),
   368 => (x"c4",x"98",x"73",x"48"),
   369 => (x"02",x"6e",x"58",x"a6"),
   370 => (x"6c",x"87",x"cc",x"c0"),
   371 => (x"c4",x"98",x"73",x"48"),
   372 => (x"05",x"6e",x"58",x"a6"),
   373 => (x"c1",x"87",x"f4",x"ff"),
   374 => (x"c0",x"1e",x"c0",x"7c"),
   375 => (x"c0",x"c1",x"d0",x"e5"),
   376 => (x"02",x"da",x"27",x"1e"),
   377 => (x"c8",x"0f",x"00",x"00"),
   378 => (x"c1",x"4a",x"70",x"86"),
   379 => (x"c0",x"05",x"aa",x"b7"),
   380 => (x"4d",x"c1",x"87",x"c2"),
   381 => (x"05",x"ad",x"b7",x"c2"),
   382 => (x"27",x"87",x"d3",x"c0"),
   383 => (x"00",x"00",x"06",x"90"),
   384 => (x"00",x"6e",x"27",x"1e"),
   385 => (x"c4",x"0f",x"00",x"00"),
   386 => (x"c1",x"48",x"c0",x"86"),
   387 => (x"8d",x"c1",x"87",x"f7"),
   388 => (x"fe",x"05",x"9d",x"75"),
   389 => (x"02",x"27",x"87",x"c9"),
   390 => (x"0f",x"00",x"00",x"04"),
   391 => (x"00",x"02",x"94",x"27"),
   392 => (x"90",x"27",x"58",x"00"),
   393 => (x"bf",x"00",x"00",x"02"),
   394 => (x"87",x"d0",x"c0",x"05"),
   395 => (x"ff",x"c0",x"1e",x"c1"),
   396 => (x"1e",x"d0",x"c1",x"f0"),
   397 => (x"00",x"02",x"da",x"27"),
   398 => (x"86",x"c8",x"0f",x"00"),
   399 => (x"c3",x"49",x"d4",x"ff"),
   400 => (x"2b",x"27",x"79",x"ff"),
   401 => (x"0f",x"00",x"00",x"09"),
   402 => (x"00",x"1a",x"c0",x"27"),
   403 => (x"bc",x"27",x"58",x"00"),
   404 => (x"bf",x"00",x"00",x"1a"),
   405 => (x"06",x"99",x"27",x"1e"),
   406 => (x"27",x"1e",x"00",x"00"),
   407 => (x"00",x"00",x"01",x"50"),
   408 => (x"6c",x"86",x"c8",x"0f"),
   409 => (x"c4",x"98",x"73",x"48"),
   410 => (x"02",x"6e",x"58",x"a6"),
   411 => (x"6c",x"87",x"cc",x"c0"),
   412 => (x"c4",x"98",x"73",x"48"),
   413 => (x"05",x"6e",x"58",x"a6"),
   414 => (x"c0",x"87",x"f4",x"ff"),
   415 => (x"49",x"d4",x"ff",x"7c"),
   416 => (x"c1",x"79",x"ff",x"c3"),
   417 => (x"4d",x"26",x"26",x"48"),
   418 => (x"4b",x"26",x"4c",x"26"),
   419 => (x"4f",x"26",x"4a",x"26"),
   420 => (x"52",x"52",x"45",x"49"),
   421 => (x"49",x"50",x"53",x"00"),
   422 => (x"20",x"44",x"53",x"00"),
   423 => (x"64",x"72",x"61",x"63"),
   424 => (x"7a",x"69",x"73",x"20"),
   425 => (x"73",x"69",x"20",x"65"),
   426 => (x"0a",x"64",x"25",x"20"),
   427 => (x"5a",x"5e",x"0e",x"00"),
   428 => (x"0e",x"5d",x"5c",x"5b"),
   429 => (x"4d",x"ff",x"c3",x"1e"),
   430 => (x"75",x"4c",x"d4",x"ff"),
   431 => (x"bf",x"d0",x"ff",x"7c"),
   432 => (x"c0",x"c0",x"c8",x"48"),
   433 => (x"58",x"a6",x"c4",x"98"),
   434 => (x"d2",x"c0",x"02",x"6e"),
   435 => (x"c0",x"c0",x"c8",x"87"),
   436 => (x"bf",x"d0",x"ff",x"4a"),
   437 => (x"c4",x"98",x"72",x"48"),
   438 => (x"05",x"6e",x"58",x"a6"),
   439 => (x"ff",x"87",x"f2",x"ff"),
   440 => (x"c1",x"c4",x"49",x"d0"),
   441 => (x"d8",x"7c",x"75",x"79"),
   442 => (x"ff",x"c0",x"1e",x"66"),
   443 => (x"1e",x"d8",x"c1",x"f0"),
   444 => (x"00",x"02",x"da",x"27"),
   445 => (x"86",x"c8",x"0f",x"00"),
   446 => (x"9a",x"72",x"4a",x"70"),
   447 => (x"87",x"d3",x"c0",x"02"),
   448 => (x"00",x"07",x"b5",x"27"),
   449 => (x"6e",x"27",x"1e",x"00"),
   450 => (x"0f",x"00",x"00",x"00"),
   451 => (x"48",x"c1",x"86",x"c4"),
   452 => (x"75",x"87",x"d7",x"c2"),
   453 => (x"7c",x"fe",x"c3",x"7c"),
   454 => (x"79",x"c0",x"49",x"76"),
   455 => (x"4a",x"bf",x"66",x"dc"),
   456 => (x"b7",x"d8",x"4b",x"72"),
   457 => (x"75",x"48",x"73",x"2b"),
   458 => (x"72",x"7c",x"70",x"98"),
   459 => (x"2b",x"b7",x"d0",x"4b"),
   460 => (x"98",x"75",x"48",x"73"),
   461 => (x"4b",x"72",x"7c",x"70"),
   462 => (x"73",x"2b",x"b7",x"c8"),
   463 => (x"70",x"98",x"75",x"48"),
   464 => (x"75",x"48",x"72",x"7c"),
   465 => (x"dc",x"7c",x"70",x"98"),
   466 => (x"80",x"c4",x"48",x"66"),
   467 => (x"58",x"a6",x"e0",x"c0"),
   468 => (x"80",x"c1",x"48",x"6e"),
   469 => (x"6e",x"58",x"a6",x"c4"),
   470 => (x"b7",x"c0",x"c2",x"49"),
   471 => (x"fb",x"fe",x"04",x"a9"),
   472 => (x"75",x"7c",x"75",x"87"),
   473 => (x"d8",x"7c",x"75",x"7c"),
   474 => (x"75",x"4b",x"e0",x"da"),
   475 => (x"75",x"4a",x"6c",x"7c"),
   476 => (x"05",x"9a",x"72",x"9a"),
   477 => (x"c1",x"87",x"c8",x"c0"),
   478 => (x"05",x"9b",x"73",x"8b"),
   479 => (x"75",x"87",x"ec",x"ff"),
   480 => (x"bf",x"d0",x"ff",x"7c"),
   481 => (x"c0",x"c0",x"c8",x"48"),
   482 => (x"58",x"a6",x"c4",x"98"),
   483 => (x"d2",x"c0",x"02",x"6e"),
   484 => (x"c0",x"c0",x"c8",x"87"),
   485 => (x"bf",x"d0",x"ff",x"4a"),
   486 => (x"c4",x"98",x"72",x"48"),
   487 => (x"05",x"6e",x"58",x"a6"),
   488 => (x"ff",x"87",x"f2",x"ff"),
   489 => (x"79",x"c0",x"49",x"d0"),
   490 => (x"26",x"26",x"48",x"c0"),
   491 => (x"26",x"4c",x"26",x"4d"),
   492 => (x"26",x"4a",x"26",x"4b"),
   493 => (x"69",x"72",x"57",x"4f"),
   494 => (x"66",x"20",x"65",x"74"),
   495 => (x"65",x"6c",x"69",x"61"),
   496 => (x"0e",x"00",x"0a",x"64"),
   497 => (x"5c",x"5b",x"5a",x"5e"),
   498 => (x"d8",x"1e",x"0e",x"5d"),
   499 => (x"66",x"dc",x"4c",x"66"),
   500 => (x"c0",x"49",x"76",x"4b"),
   501 => (x"cd",x"ee",x"c5",x"79"),
   502 => (x"d4",x"ff",x"4d",x"df"),
   503 => (x"79",x"ff",x"c3",x"49"),
   504 => (x"4a",x"bf",x"d4",x"ff"),
   505 => (x"c3",x"9a",x"ff",x"c3"),
   506 => (x"05",x"aa",x"b7",x"fe"),
   507 => (x"27",x"87",x"e5",x"c1"),
   508 => (x"00",x"00",x"1a",x"b8"),
   509 => (x"c4",x"79",x"c0",x"49"),
   510 => (x"c0",x"04",x"ab",x"b7"),
   511 => (x"94",x"27",x"87",x"e4"),
   512 => (x"0f",x"00",x"00",x"02"),
   513 => (x"7c",x"72",x"4a",x"70"),
   514 => (x"b8",x"27",x"84",x"c4"),
   515 => (x"bf",x"00",x"00",x"1a"),
   516 => (x"27",x"80",x"72",x"48"),
   517 => (x"00",x"00",x"1a",x"bc"),
   518 => (x"c4",x"8b",x"c4",x"58"),
   519 => (x"ff",x"03",x"ab",x"b7"),
   520 => (x"b7",x"c0",x"87",x"dc"),
   521 => (x"e5",x"c0",x"06",x"ab"),
   522 => (x"4d",x"d4",x"ff",x"87"),
   523 => (x"6d",x"7d",x"ff",x"c3"),
   524 => (x"7c",x"97",x"72",x"4a"),
   525 => (x"b8",x"27",x"84",x"c1"),
   526 => (x"bf",x"00",x"00",x"1a"),
   527 => (x"27",x"80",x"72",x"48"),
   528 => (x"00",x"00",x"1a",x"bc"),
   529 => (x"c0",x"8b",x"c1",x"58"),
   530 => (x"ff",x"01",x"ab",x"b7"),
   531 => (x"4d",x"c1",x"87",x"de"),
   532 => (x"79",x"c1",x"49",x"76"),
   533 => (x"9d",x"75",x"8d",x"c1"),
   534 => (x"87",x"fe",x"fd",x"05"),
   535 => (x"c3",x"49",x"d4",x"ff"),
   536 => (x"48",x"6e",x"79",x"ff"),
   537 => (x"26",x"4d",x"26",x"26"),
   538 => (x"26",x"4b",x"26",x"4c"),
   539 => (x"0e",x"4f",x"26",x"4a"),
   540 => (x"5c",x"5b",x"5a",x"5e"),
   541 => (x"ff",x"1e",x"0e",x"5d"),
   542 => (x"c0",x"c8",x"4b",x"d0"),
   543 => (x"4c",x"c0",x"4a",x"c0"),
   544 => (x"c3",x"49",x"d4",x"ff"),
   545 => (x"48",x"6b",x"79",x"ff"),
   546 => (x"a6",x"c4",x"98",x"72"),
   547 => (x"c0",x"02",x"6e",x"58"),
   548 => (x"48",x"6b",x"87",x"cc"),
   549 => (x"a6",x"c4",x"98",x"72"),
   550 => (x"ff",x"05",x"6e",x"58"),
   551 => (x"c1",x"c4",x"87",x"f4"),
   552 => (x"49",x"d4",x"ff",x"7b"),
   553 => (x"d8",x"79",x"ff",x"c3"),
   554 => (x"ff",x"c0",x"1e",x"66"),
   555 => (x"1e",x"d1",x"c1",x"f0"),
   556 => (x"00",x"02",x"da",x"27"),
   557 => (x"86",x"c8",x"0f",x"00"),
   558 => (x"9d",x"75",x"4d",x"70"),
   559 => (x"87",x"d6",x"c0",x"02"),
   560 => (x"66",x"dc",x"1e",x"75"),
   561 => (x"09",x"0b",x"27",x"1e"),
   562 => (x"27",x"1e",x"00",x"00"),
   563 => (x"00",x"00",x"01",x"50"),
   564 => (x"c0",x"86",x"cc",x"0f"),
   565 => (x"c0",x"c8",x"87",x"e8"),
   566 => (x"66",x"e0",x"c0",x"1e"),
   567 => (x"87",x"e3",x"fb",x"1e"),
   568 => (x"4c",x"70",x"86",x"c8"),
   569 => (x"98",x"72",x"48",x"6b"),
   570 => (x"6e",x"58",x"a6",x"c4"),
   571 => (x"87",x"cc",x"c0",x"02"),
   572 => (x"98",x"72",x"48",x"6b"),
   573 => (x"6e",x"58",x"a6",x"c4"),
   574 => (x"87",x"f4",x"ff",x"05"),
   575 => (x"48",x"74",x"7b",x"c0"),
   576 => (x"26",x"4d",x"26",x"26"),
   577 => (x"26",x"4b",x"26",x"4c"),
   578 => (x"52",x"4f",x"26",x"4a"),
   579 => (x"20",x"64",x"61",x"65"),
   580 => (x"6d",x"6d",x"6f",x"63"),
   581 => (x"20",x"64",x"6e",x"61"),
   582 => (x"6c",x"69",x"61",x"66"),
   583 => (x"61",x"20",x"64",x"65"),
   584 => (x"64",x"25",x"20",x"74"),
   585 => (x"64",x"25",x"28",x"20"),
   586 => (x"0e",x"00",x"0a",x"29"),
   587 => (x"5c",x"5b",x"5a",x"5e"),
   588 => (x"c0",x"1e",x"0e",x"5d"),
   589 => (x"f0",x"ff",x"c0",x"1e"),
   590 => (x"27",x"1e",x"c9",x"c1"),
   591 => (x"00",x"00",x"02",x"da"),
   592 => (x"d2",x"86",x"c8",x"0f"),
   593 => (x"1a",x"c8",x"27",x"1e"),
   594 => (x"f9",x"1e",x"00",x"00"),
   595 => (x"86",x"c8",x"87",x"f5"),
   596 => (x"85",x"c1",x"4d",x"c0"),
   597 => (x"04",x"ad",x"b7",x"d2"),
   598 => (x"27",x"87",x"f7",x"ff"),
   599 => (x"00",x"00",x"1a",x"c8"),
   600 => (x"c3",x"4a",x"bf",x"97"),
   601 => (x"c0",x"c1",x"9a",x"c0"),
   602 => (x"c0",x"05",x"aa",x"b7"),
   603 => (x"cf",x"27",x"87",x"f2"),
   604 => (x"97",x"00",x"00",x"1a"),
   605 => (x"32",x"d0",x"4a",x"bf"),
   606 => (x"00",x"1a",x"d0",x"27"),
   607 => (x"4b",x"bf",x"97",x"00"),
   608 => (x"4a",x"72",x"33",x"c8"),
   609 => (x"d1",x"27",x"b2",x"73"),
   610 => (x"97",x"00",x"00",x"1a"),
   611 => (x"4a",x"72",x"4b",x"bf"),
   612 => (x"ff",x"cf",x"b2",x"73"),
   613 => (x"72",x"9a",x"ff",x"ff"),
   614 => (x"ca",x"85",x"c1",x"4d"),
   615 => (x"87",x"cb",x"c3",x"35"),
   616 => (x"00",x"1a",x"d1",x"27"),
   617 => (x"4a",x"bf",x"97",x"00"),
   618 => (x"9a",x"c6",x"32",x"c1"),
   619 => (x"00",x"1a",x"d2",x"27"),
   620 => (x"4b",x"bf",x"97",x"00"),
   621 => (x"72",x"2b",x"b7",x"c7"),
   622 => (x"27",x"b2",x"73",x"4a"),
   623 => (x"00",x"00",x"1a",x"cd"),
   624 => (x"73",x"4b",x"bf",x"97"),
   625 => (x"c4",x"98",x"cf",x"48"),
   626 => (x"ce",x"27",x"58",x"a6"),
   627 => (x"97",x"00",x"00",x"1a"),
   628 => (x"9b",x"c3",x"4b",x"bf"),
   629 => (x"cf",x"27",x"33",x"ca"),
   630 => (x"97",x"00",x"00",x"1a"),
   631 => (x"34",x"c2",x"4c",x"bf"),
   632 => (x"b3",x"74",x"4b",x"73"),
   633 => (x"00",x"1a",x"d0",x"27"),
   634 => (x"4c",x"bf",x"97",x"00"),
   635 => (x"c6",x"9c",x"c0",x"c3"),
   636 => (x"4b",x"73",x"2c",x"b7"),
   637 => (x"1e",x"73",x"b3",x"74"),
   638 => (x"72",x"1e",x"66",x"c4"),
   639 => (x"0a",x"78",x"27",x"1e"),
   640 => (x"27",x"1e",x"00",x"00"),
   641 => (x"00",x"00",x"01",x"50"),
   642 => (x"c2",x"86",x"d0",x"0f"),
   643 => (x"72",x"48",x"c1",x"82"),
   644 => (x"72",x"4a",x"70",x"30"),
   645 => (x"0a",x"a5",x"27",x"1e"),
   646 => (x"27",x"1e",x"00",x"00"),
   647 => (x"00",x"00",x"01",x"50"),
   648 => (x"c1",x"86",x"c8",x"0f"),
   649 => (x"c4",x"30",x"6e",x"48"),
   650 => (x"83",x"c1",x"58",x"a6"),
   651 => (x"95",x"72",x"4d",x"73"),
   652 => (x"1e",x"75",x"1e",x"6e"),
   653 => (x"00",x"0a",x"ae",x"27"),
   654 => (x"50",x"27",x"1e",x"00"),
   655 => (x"0f",x"00",x"00",x"01"),
   656 => (x"49",x"6e",x"86",x"cc"),
   657 => (x"a9",x"b7",x"c0",x"c8"),
   658 => (x"87",x"cf",x"c0",x"06"),
   659 => (x"35",x"c1",x"4a",x"6e"),
   660 => (x"c8",x"2a",x"b7",x"c1"),
   661 => (x"01",x"aa",x"b7",x"c0"),
   662 => (x"75",x"87",x"f3",x"ff"),
   663 => (x"0a",x"c4",x"27",x"1e"),
   664 => (x"27",x"1e",x"00",x"00"),
   665 => (x"00",x"00",x"01",x"50"),
   666 => (x"75",x"86",x"c8",x"0f"),
   667 => (x"4d",x"26",x"26",x"48"),
   668 => (x"4b",x"26",x"4c",x"26"),
   669 => (x"4f",x"26",x"4a",x"26"),
   670 => (x"69",x"73",x"5f",x"63"),
   671 => (x"6d",x"5f",x"65",x"7a"),
   672 => (x"3a",x"74",x"6c",x"75"),
   673 => (x"2c",x"64",x"25",x"20"),
   674 => (x"61",x"65",x"72",x"20"),
   675 => (x"6c",x"62",x"5f",x"64"),
   676 => (x"6e",x"65",x"6c",x"5f"),
   677 => (x"64",x"25",x"20",x"3a"),
   678 => (x"73",x"63",x"20",x"2c"),
   679 => (x"3a",x"65",x"7a",x"69"),
   680 => (x"0a",x"64",x"25",x"20"),
   681 => (x"6c",x"75",x"4d",x"00"),
   682 => (x"64",x"25",x"20",x"74"),
   683 => (x"64",x"25",x"00",x"0a"),
   684 => (x"6f",x"6c",x"62",x"20"),
   685 => (x"20",x"73",x"6b",x"63"),
   686 => (x"73",x"20",x"66",x"6f"),
   687 => (x"20",x"65",x"7a",x"69"),
   688 => (x"00",x"0a",x"64",x"25"),
   689 => (x"62",x"20",x"64",x"25"),
   690 => (x"6b",x"63",x"6f",x"6c"),
   691 => (x"66",x"6f",x"20",x"73"),
   692 => (x"32",x"31",x"35",x"20"),
   693 => (x"74",x"79",x"62",x"20"),
   694 => (x"00",x"0a",x"73",x"65"),
   695 => (x"5b",x"5a",x"5e",x"0e"),
   696 => (x"d4",x"0e",x"5d",x"5c"),
   697 => (x"4c",x"c0",x"4d",x"66"),
   698 => (x"c0",x"49",x"66",x"dc"),
   699 => (x"c0",x"06",x"a9",x"b7"),
   700 => (x"4b",x"15",x"87",x"fb"),
   701 => (x"c0",x"c0",x"c0",x"c1"),
   702 => (x"c0",x"c4",x"93",x"c0"),
   703 => (x"d8",x"4b",x"93",x"b7"),
   704 => (x"4a",x"bf",x"97",x"66"),
   705 => (x"c0",x"c0",x"c0",x"c1"),
   706 => (x"c0",x"c4",x"92",x"c0"),
   707 => (x"d8",x"4a",x"92",x"b7"),
   708 => (x"80",x"c1",x"48",x"66"),
   709 => (x"72",x"58",x"a6",x"dc"),
   710 => (x"c0",x"02",x"ab",x"b7"),
   711 => (x"48",x"c1",x"87",x"c5"),
   712 => (x"c1",x"87",x"cc",x"c0"),
   713 => (x"b7",x"66",x"dc",x"84"),
   714 => (x"c5",x"ff",x"04",x"ac"),
   715 => (x"26",x"48",x"c0",x"87"),
   716 => (x"26",x"4c",x"26",x"4d"),
   717 => (x"26",x"4a",x"26",x"4b"),
   718 => (x"5a",x"5e",x"0e",x"4f"),
   719 => (x"0e",x"5d",x"5c",x"5b"),
   720 => (x"00",x"1c",x"f0",x"27"),
   721 => (x"79",x"c0",x"49",x"00"),
   722 => (x"00",x"19",x"9d",x"27"),
   723 => (x"6e",x"27",x"1e",x"00"),
   724 => (x"0f",x"00",x"00",x"00"),
   725 => (x"e8",x"27",x"86",x"c4"),
   726 => (x"1e",x"00",x"00",x"1a"),
   727 => (x"6f",x"27",x"1e",x"c0"),
   728 => (x"0f",x"00",x"00",x"08"),
   729 => (x"4a",x"70",x"86",x"c8"),
   730 => (x"c0",x"05",x"9a",x"72"),
   731 => (x"c9",x"27",x"87",x"d3"),
   732 => (x"1e",x"00",x"00",x"18"),
   733 => (x"00",x"00",x"6e",x"27"),
   734 => (x"86",x"c4",x"0f",x"00"),
   735 => (x"d8",x"cf",x"48",x"c0"),
   736 => (x"19",x"aa",x"27",x"87"),
   737 => (x"27",x"1e",x"00",x"00"),
   738 => (x"00",x"00",x"00",x"6e"),
   739 => (x"c0",x"86",x"c4",x"0f"),
   740 => (x"1d",x"1c",x"27",x"4c"),
   741 => (x"c1",x"49",x"00",x"00"),
   742 => (x"27",x"1e",x"c8",x"79"),
   743 => (x"00",x"00",x"19",x"c1"),
   744 => (x"1b",x"1e",x"27",x"1e"),
   745 => (x"27",x"1e",x"00",x"00"),
   746 => (x"00",x"00",x"0a",x"dc"),
   747 => (x"70",x"86",x"cc",x"0f"),
   748 => (x"05",x"9a",x"72",x"4a"),
   749 => (x"27",x"87",x"c8",x"c0"),
   750 => (x"00",x"00",x"1d",x"1c"),
   751 => (x"c8",x"79",x"c0",x"49"),
   752 => (x"19",x"ca",x"27",x"1e"),
   753 => (x"27",x"1e",x"00",x"00"),
   754 => (x"00",x"00",x"1b",x"3a"),
   755 => (x"0a",x"dc",x"27",x"1e"),
   756 => (x"cc",x"0f",x"00",x"00"),
   757 => (x"72",x"4a",x"70",x"86"),
   758 => (x"c8",x"c0",x"05",x"9a"),
   759 => (x"1d",x"1c",x"27",x"87"),
   760 => (x"c0",x"49",x"00",x"00"),
   761 => (x"1d",x"1c",x"27",x"79"),
   762 => (x"1e",x"bf",x"00",x"00"),
   763 => (x"00",x"19",x"d3",x"27"),
   764 => (x"50",x"27",x"1e",x"00"),
   765 => (x"0f",x"00",x"00",x"01"),
   766 => (x"1c",x"27",x"86",x"c8"),
   767 => (x"bf",x"00",x"00",x"1d"),
   768 => (x"87",x"c0",x"c3",x"02"),
   769 => (x"00",x"1a",x"e8",x"27"),
   770 => (x"a6",x"27",x"4d",x"00"),
   771 => (x"4b",x"00",x"00",x"1c"),
   772 => (x"00",x"1c",x"e6",x"27"),
   773 => (x"4a",x"bf",x"9f",x"00"),
   774 => (x"e6",x"27",x"1e",x"72"),
   775 => (x"4a",x"00",x"00",x"1c"),
   776 => (x"00",x"1a",x"e8",x"27"),
   777 => (x"1e",x"72",x"8a",x"00"),
   778 => (x"c0",x"c8",x"1e",x"d0"),
   779 => (x"18",x"fb",x"27",x"1e"),
   780 => (x"27",x"1e",x"00",x"00"),
   781 => (x"00",x"00",x"01",x"50"),
   782 => (x"73",x"86",x"d4",x"0f"),
   783 => (x"6a",x"82",x"c8",x"4a"),
   784 => (x"1c",x"e6",x"27",x"4c"),
   785 => (x"bf",x"9f",x"00",x"00"),
   786 => (x"ea",x"d6",x"c5",x"4a"),
   787 => (x"c0",x"05",x"aa",x"b7"),
   788 => (x"4a",x"73",x"87",x"d3"),
   789 => (x"1e",x"6a",x"82",x"c8"),
   790 => (x"00",x"12",x"c4",x"27"),
   791 => (x"86",x"c4",x"0f",x"00"),
   792 => (x"e4",x"c0",x"4c",x"70"),
   793 => (x"c7",x"4a",x"75",x"87"),
   794 => (x"6a",x"9f",x"82",x"fe"),
   795 => (x"d5",x"e9",x"ca",x"4a"),
   796 => (x"c0",x"02",x"aa",x"b7"),
   797 => (x"dd",x"27",x"87",x"d3"),
   798 => (x"1e",x"00",x"00",x"18"),
   799 => (x"00",x"00",x"6e",x"27"),
   800 => (x"86",x"c4",x"0f",x"00"),
   801 => (x"d0",x"cb",x"48",x"c0"),
   802 => (x"27",x"1e",x"74",x"87"),
   803 => (x"00",x"00",x"19",x"38"),
   804 => (x"01",x"50",x"27",x"1e"),
   805 => (x"c8",x"0f",x"00",x"00"),
   806 => (x"1a",x"e8",x"27",x"86"),
   807 => (x"74",x"1e",x"00",x"00"),
   808 => (x"08",x"6f",x"27",x"1e"),
   809 => (x"c8",x"0f",x"00",x"00"),
   810 => (x"72",x"4a",x"70",x"86"),
   811 => (x"c5",x"c0",x"05",x"9a"),
   812 => (x"ca",x"48",x"c0",x"87"),
   813 => (x"50",x"27",x"87",x"e3"),
   814 => (x"1e",x"00",x"00",x"19"),
   815 => (x"00",x"00",x"6e",x"27"),
   816 => (x"86",x"c4",x"0f",x"00"),
   817 => (x"00",x"19",x"e6",x"27"),
   818 => (x"50",x"27",x"1e",x"00"),
   819 => (x"0f",x"00",x"00",x"01"),
   820 => (x"1e",x"c8",x"86",x"c4"),
   821 => (x"00",x"19",x"fe",x"27"),
   822 => (x"3a",x"27",x"1e",x"00"),
   823 => (x"1e",x"00",x"00",x"1b"),
   824 => (x"00",x"0a",x"dc",x"27"),
   825 => (x"86",x"cc",x"0f",x"00"),
   826 => (x"9a",x"72",x"4a",x"70"),
   827 => (x"87",x"cb",x"c0",x"05"),
   828 => (x"00",x"1c",x"f0",x"27"),
   829 => (x"79",x"c1",x"49",x"00"),
   830 => (x"c8",x"87",x"f1",x"c0"),
   831 => (x"1a",x"07",x"27",x"1e"),
   832 => (x"27",x"1e",x"00",x"00"),
   833 => (x"00",x"00",x"1b",x"1e"),
   834 => (x"0a",x"dc",x"27",x"1e"),
   835 => (x"cc",x"0f",x"00",x"00"),
   836 => (x"72",x"4a",x"70",x"86"),
   837 => (x"d3",x"c0",x"02",x"9a"),
   838 => (x"19",x"77",x"27",x"87"),
   839 => (x"27",x"1e",x"00",x"00"),
   840 => (x"00",x"00",x"01",x"50"),
   841 => (x"c0",x"86",x"c4",x"0f"),
   842 => (x"87",x"ed",x"c8",x"48"),
   843 => (x"00",x"1c",x"e6",x"27"),
   844 => (x"4a",x"bf",x"97",x"00"),
   845 => (x"aa",x"b7",x"d5",x"c1"),
   846 => (x"87",x"d0",x"c0",x"05"),
   847 => (x"00",x"1c",x"e7",x"27"),
   848 => (x"4a",x"bf",x"97",x"00"),
   849 => (x"aa",x"b7",x"ea",x"c2"),
   850 => (x"87",x"c5",x"c0",x"02"),
   851 => (x"c8",x"c8",x"48",x"c0"),
   852 => (x"1a",x"e8",x"27",x"87"),
   853 => (x"bf",x"97",x"00",x"00"),
   854 => (x"b7",x"e9",x"c3",x"4a"),
   855 => (x"d5",x"c0",x"02",x"aa"),
   856 => (x"1a",x"e8",x"27",x"87"),
   857 => (x"bf",x"97",x"00",x"00"),
   858 => (x"b7",x"eb",x"c3",x"4a"),
   859 => (x"c5",x"c0",x"02",x"aa"),
   860 => (x"c7",x"48",x"c0",x"87"),
   861 => (x"f3",x"27",x"87",x"e3"),
   862 => (x"97",x"00",x"00",x"1a"),
   863 => (x"9a",x"72",x"4a",x"bf"),
   864 => (x"87",x"cf",x"c0",x"05"),
   865 => (x"00",x"1a",x"f4",x"27"),
   866 => (x"4a",x"bf",x"97",x"00"),
   867 => (x"02",x"aa",x"b7",x"c2"),
   868 => (x"c0",x"87",x"c5",x"c0"),
   869 => (x"87",x"c1",x"c7",x"48"),
   870 => (x"00",x"1a",x"f5",x"27"),
   871 => (x"48",x"bf",x"97",x"00"),
   872 => (x"00",x"1c",x"ec",x"27"),
   873 => (x"e8",x"27",x"58",x"00"),
   874 => (x"bf",x"00",x"00",x"1c"),
   875 => (x"c1",x"4b",x"72",x"4a"),
   876 => (x"1c",x"ec",x"27",x"8b"),
   877 => (x"73",x"49",x"00",x"00"),
   878 => (x"72",x"1e",x"73",x"79"),
   879 => (x"1a",x"10",x"27",x"1e"),
   880 => (x"27",x"1e",x"00",x"00"),
   881 => (x"00",x"00",x"01",x"50"),
   882 => (x"27",x"86",x"cc",x"0f"),
   883 => (x"00",x"00",x"1a",x"f6"),
   884 => (x"74",x"4a",x"bf",x"97"),
   885 => (x"1a",x"f7",x"27",x"82"),
   886 => (x"bf",x"97",x"00",x"00"),
   887 => (x"73",x"33",x"c8",x"4b"),
   888 => (x"27",x"80",x"72",x"48"),
   889 => (x"00",x"00",x"1d",x"00"),
   890 => (x"1a",x"f8",x"27",x"58"),
   891 => (x"bf",x"97",x"00",x"00"),
   892 => (x"1d",x"14",x"27",x"48"),
   893 => (x"27",x"58",x"00",x"00"),
   894 => (x"00",x"00",x"1c",x"f0"),
   895 => (x"df",x"c3",x"02",x"bf"),
   896 => (x"27",x"1e",x"c8",x"87"),
   897 => (x"00",x"00",x"19",x"94"),
   898 => (x"1b",x"3a",x"27",x"1e"),
   899 => (x"27",x"1e",x"00",x"00"),
   900 => (x"00",x"00",x"0a",x"dc"),
   901 => (x"70",x"86",x"cc",x"0f"),
   902 => (x"02",x"9a",x"72",x"4a"),
   903 => (x"c0",x"87",x"c5",x"c0"),
   904 => (x"87",x"f5",x"c4",x"48"),
   905 => (x"00",x"1c",x"e8",x"27"),
   906 => (x"73",x"4b",x"bf",x"00"),
   907 => (x"27",x"30",x"c4",x"48"),
   908 => (x"00",x"00",x"1d",x"18"),
   909 => (x"1d",x"0c",x"27",x"58"),
   910 => (x"73",x"49",x"00",x"00"),
   911 => (x"1b",x"0d",x"27",x"79"),
   912 => (x"bf",x"97",x"00",x"00"),
   913 => (x"27",x"32",x"c8",x"4a"),
   914 => (x"00",x"00",x"1b",x"0c"),
   915 => (x"72",x"4c",x"bf",x"97"),
   916 => (x"27",x"82",x"74",x"4a"),
   917 => (x"00",x"00",x"1b",x"0e"),
   918 => (x"d0",x"4c",x"bf",x"97"),
   919 => (x"74",x"4a",x"72",x"34"),
   920 => (x"1b",x"0f",x"27",x"82"),
   921 => (x"bf",x"97",x"00",x"00"),
   922 => (x"72",x"34",x"d8",x"4c"),
   923 => (x"27",x"82",x"74",x"4a"),
   924 => (x"00",x"00",x"1d",x"18"),
   925 => (x"72",x"79",x"72",x"49"),
   926 => (x"1d",x"10",x"27",x"4a"),
   927 => (x"92",x"bf",x"00",x"00"),
   928 => (x"fc",x"27",x"4a",x"72"),
   929 => (x"bf",x"00",x"00",x"1c"),
   930 => (x"1d",x"00",x"27",x"82"),
   931 => (x"72",x"49",x"00",x"00"),
   932 => (x"1b",x"15",x"27",x"79"),
   933 => (x"bf",x"97",x"00",x"00"),
   934 => (x"27",x"34",x"c8",x"4c"),
   935 => (x"00",x"00",x"1b",x"14"),
   936 => (x"74",x"4d",x"bf",x"97"),
   937 => (x"27",x"84",x"75",x"4c"),
   938 => (x"00",x"00",x"1b",x"16"),
   939 => (x"d0",x"4d",x"bf",x"97"),
   940 => (x"75",x"4c",x"74",x"35"),
   941 => (x"1b",x"17",x"27",x"84"),
   942 => (x"bf",x"97",x"00",x"00"),
   943 => (x"d8",x"9d",x"cf",x"4d"),
   944 => (x"75",x"4c",x"74",x"35"),
   945 => (x"1d",x"04",x"27",x"84"),
   946 => (x"74",x"49",x"00",x"00"),
   947 => (x"73",x"8c",x"c2",x"79"),
   948 => (x"73",x"93",x"74",x"4b"),
   949 => (x"27",x"80",x"72",x"48"),
   950 => (x"00",x"00",x"1d",x"0c"),
   951 => (x"87",x"f7",x"c1",x"58"),
   952 => (x"00",x"1a",x"fa",x"27"),
   953 => (x"4a",x"bf",x"97",x"00"),
   954 => (x"f9",x"27",x"32",x"c8"),
   955 => (x"97",x"00",x"00",x"1a"),
   956 => (x"4a",x"72",x"4b",x"bf"),
   957 => (x"14",x"27",x"82",x"73"),
   958 => (x"49",x"00",x"00",x"1d"),
   959 => (x"32",x"c5",x"79",x"72"),
   960 => (x"c9",x"82",x"ff",x"c7"),
   961 => (x"1d",x"0c",x"27",x"2a"),
   962 => (x"72",x"49",x"00",x"00"),
   963 => (x"1a",x"ff",x"27",x"79"),
   964 => (x"bf",x"97",x"00",x"00"),
   965 => (x"27",x"33",x"c8",x"4b"),
   966 => (x"00",x"00",x"1a",x"fe"),
   967 => (x"73",x"4c",x"bf",x"97"),
   968 => (x"27",x"83",x"74",x"4b"),
   969 => (x"00",x"00",x"1d",x"18"),
   970 => (x"73",x"79",x"73",x"49"),
   971 => (x"1d",x"10",x"27",x"4b"),
   972 => (x"93",x"bf",x"00",x"00"),
   973 => (x"fc",x"27",x"4b",x"73"),
   974 => (x"bf",x"00",x"00",x"1c"),
   975 => (x"1d",x"08",x"27",x"83"),
   976 => (x"73",x"49",x"00",x"00"),
   977 => (x"1d",x"04",x"27",x"79"),
   978 => (x"c0",x"49",x"00",x"00"),
   979 => (x"72",x"48",x"73",x"79"),
   980 => (x"1d",x"04",x"27",x"80"),
   981 => (x"c1",x"58",x"00",x"00"),
   982 => (x"26",x"4d",x"26",x"48"),
   983 => (x"26",x"4b",x"26",x"4c"),
   984 => (x"0e",x"4f",x"26",x"4a"),
   985 => (x"5c",x"5b",x"5a",x"5e"),
   986 => (x"f0",x"27",x"0e",x"5d"),
   987 => (x"bf",x"00",x"00",x"1c"),
   988 => (x"87",x"cf",x"c0",x"02"),
   989 => (x"c7",x"4c",x"66",x"d4"),
   990 => (x"66",x"d4",x"2c",x"b7"),
   991 => (x"9b",x"ff",x"c1",x"4b"),
   992 => (x"d4",x"87",x"cc",x"c0"),
   993 => (x"b7",x"c8",x"4c",x"66"),
   994 => (x"4b",x"66",x"d4",x"2c"),
   995 => (x"27",x"9b",x"ff",x"c3"),
   996 => (x"00",x"00",x"1a",x"e8"),
   997 => (x"1c",x"fc",x"27",x"1e"),
   998 => (x"4a",x"bf",x"00",x"00"),
   999 => (x"1e",x"72",x"82",x"74"),
  1000 => (x"00",x"08",x"6f",x"27"),
  1001 => (x"86",x"c8",x"0f",x"00"),
  1002 => (x"9a",x"72",x"4a",x"70"),
  1003 => (x"87",x"c5",x"c0",x"05"),
  1004 => (x"f2",x"c0",x"48",x"c0"),
  1005 => (x"1c",x"f0",x"27",x"87"),
  1006 => (x"02",x"bf",x"00",x"00"),
  1007 => (x"73",x"87",x"d7",x"c0"),
  1008 => (x"72",x"92",x"c4",x"4a"),
  1009 => (x"1a",x"e8",x"27",x"4a"),
  1010 => (x"6a",x"82",x"00",x"00"),
  1011 => (x"ff",x"ff",x"cf",x"4d"),
  1012 => (x"c0",x"9d",x"ff",x"ff"),
  1013 => (x"4a",x"73",x"87",x"cf"),
  1014 => (x"4a",x"72",x"92",x"c2"),
  1015 => (x"00",x"1a",x"e8",x"27"),
  1016 => (x"6a",x"9f",x"82",x"00"),
  1017 => (x"26",x"48",x"75",x"4d"),
  1018 => (x"26",x"4c",x"26",x"4d"),
  1019 => (x"26",x"4a",x"26",x"4b"),
  1020 => (x"5a",x"5e",x"0e",x"4f"),
  1021 => (x"0e",x"5d",x"5c",x"5b"),
  1022 => (x"ff",x"cf",x"8e",x"cc"),
  1023 => (x"4d",x"f8",x"ff",x"ff"),
  1024 => (x"49",x"76",x"4c",x"c0"),
  1025 => (x"00",x"1d",x"04",x"27"),
  1026 => (x"c4",x"79",x"bf",x"00"),
  1027 => (x"08",x"27",x"49",x"a6"),
  1028 => (x"bf",x"00",x"00",x"1d"),
  1029 => (x"1c",x"f0",x"27",x"79"),
  1030 => (x"02",x"bf",x"00",x"00"),
  1031 => (x"27",x"87",x"cc",x"c0"),
  1032 => (x"00",x"00",x"1c",x"e8"),
  1033 => (x"32",x"c4",x"4a",x"bf"),
  1034 => (x"27",x"87",x"c9",x"c0"),
  1035 => (x"00",x"00",x"1d",x"0c"),
  1036 => (x"32",x"c4",x"4a",x"bf"),
  1037 => (x"72",x"49",x"a6",x"c8"),
  1038 => (x"c8",x"4b",x"c0",x"79"),
  1039 => (x"a9",x"c0",x"49",x"66"),
  1040 => (x"87",x"d0",x"c3",x"06"),
  1041 => (x"9a",x"cf",x"4a",x"73"),
  1042 => (x"c0",x"05",x"9a",x"72"),
  1043 => (x"e8",x"27",x"87",x"e4"),
  1044 => (x"1e",x"00",x"00",x"1a"),
  1045 => (x"c8",x"4a",x"66",x"c8"),
  1046 => (x"80",x"c1",x"48",x"66"),
  1047 => (x"72",x"58",x"a6",x"cc"),
  1048 => (x"08",x"6f",x"27",x"1e"),
  1049 => (x"c8",x"0f",x"00",x"00"),
  1050 => (x"1a",x"e8",x"27",x"86"),
  1051 => (x"c0",x"4c",x"00",x"00"),
  1052 => (x"e0",x"c0",x"87",x"c3"),
  1053 => (x"4a",x"6c",x"97",x"84"),
  1054 => (x"c2",x"02",x"9a",x"72"),
  1055 => (x"6c",x"97",x"87",x"cd"),
  1056 => (x"b7",x"e5",x"c3",x"4a"),
  1057 => (x"c2",x"c2",x"02",x"aa"),
  1058 => (x"cb",x"4a",x"74",x"87"),
  1059 => (x"4a",x"6a",x"97",x"82"),
  1060 => (x"9a",x"72",x"9a",x"d8"),
  1061 => (x"87",x"f3",x"c1",x"05"),
  1062 => (x"6e",x"27",x"1e",x"74"),
  1063 => (x"0f",x"00",x"00",x"00"),
  1064 => (x"1e",x"cb",x"86",x"c4"),
  1065 => (x"1e",x"66",x"e8",x"c0"),
  1066 => (x"dc",x"27",x"1e",x"74"),
  1067 => (x"0f",x"00",x"00",x"0a"),
  1068 => (x"4a",x"70",x"86",x"cc"),
  1069 => (x"c1",x"05",x"9a",x"72"),
  1070 => (x"4b",x"74",x"87",x"d1"),
  1071 => (x"e0",x"c0",x"83",x"dc"),
  1072 => (x"82",x"c4",x"4a",x"66"),
  1073 => (x"4b",x"74",x"7a",x"6b"),
  1074 => (x"e0",x"c0",x"83",x"da"),
  1075 => (x"82",x"c8",x"4a",x"66"),
  1076 => (x"70",x"48",x"6b",x"9f"),
  1077 => (x"27",x"4d",x"72",x"7a"),
  1078 => (x"00",x"00",x"1c",x"f0"),
  1079 => (x"d5",x"c0",x"02",x"bf"),
  1080 => (x"d4",x"4a",x"74",x"87"),
  1081 => (x"4a",x"6a",x"9f",x"82"),
  1082 => (x"9a",x"ff",x"ff",x"c0"),
  1083 => (x"30",x"d0",x"48",x"72"),
  1084 => (x"c0",x"58",x"a6",x"c4"),
  1085 => (x"49",x"76",x"87",x"c4"),
  1086 => (x"48",x"6e",x"79",x"c0"),
  1087 => (x"7d",x"70",x"80",x"6d"),
  1088 => (x"49",x"66",x"e0",x"c0"),
  1089 => (x"48",x"c1",x"79",x"c0"),
  1090 => (x"c1",x"87",x"ce",x"c1"),
  1091 => (x"ab",x"66",x"c8",x"83"),
  1092 => (x"87",x"f0",x"fc",x"04"),
  1093 => (x"ff",x"ff",x"ff",x"cf"),
  1094 => (x"f0",x"27",x"4d",x"f8"),
  1095 => (x"bf",x"00",x"00",x"1c"),
  1096 => (x"87",x"f3",x"c0",x"02"),
  1097 => (x"63",x"27",x"1e",x"6e"),
  1098 => (x"0f",x"00",x"00",x"0f"),
  1099 => (x"a6",x"c4",x"86",x"c4"),
  1100 => (x"75",x"4a",x"6e",x"58"),
  1101 => (x"02",x"aa",x"75",x"9a"),
  1102 => (x"6e",x"87",x"dc",x"c0"),
  1103 => (x"72",x"8a",x"c2",x"4a"),
  1104 => (x"1c",x"e8",x"27",x"4a"),
  1105 => (x"92",x"bf",x"00",x"00"),
  1106 => (x"00",x"1d",x"00",x"27"),
  1107 => (x"72",x"48",x"bf",x"00"),
  1108 => (x"58",x"a6",x"c8",x"80"),
  1109 => (x"c0",x"87",x"e2",x"fb"),
  1110 => (x"ff",x"ff",x"cf",x"48"),
  1111 => (x"cc",x"4d",x"f8",x"ff"),
  1112 => (x"26",x"4d",x"26",x"86"),
  1113 => (x"26",x"4b",x"26",x"4c"),
  1114 => (x"0e",x"4f",x"26",x"4a"),
  1115 => (x"0e",x"5b",x"5a",x"5e"),
  1116 => (x"4a",x"bf",x"66",x"cc"),
  1117 => (x"66",x"cc",x"82",x"c1"),
  1118 => (x"72",x"79",x"72",x"49"),
  1119 => (x"1c",x"ec",x"27",x"4a"),
  1120 => (x"9a",x"bf",x"00",x"00"),
  1121 => (x"c0",x"05",x"9a",x"72"),
  1122 => (x"66",x"cc",x"87",x"d3"),
  1123 => (x"6a",x"82",x"c8",x"4a"),
  1124 => (x"0f",x"63",x"27",x"1e"),
  1125 => (x"c4",x"0f",x"00",x"00"),
  1126 => (x"73",x"4b",x"70",x"86"),
  1127 => (x"26",x"48",x"c1",x"7a"),
  1128 => (x"26",x"4a",x"26",x"4b"),
  1129 => (x"5a",x"5e",x"0e",x"4f"),
  1130 => (x"00",x"27",x"0e",x"5b"),
  1131 => (x"bf",x"00",x"00",x"1d"),
  1132 => (x"4b",x"66",x"cc",x"4a"),
  1133 => (x"4b",x"6b",x"83",x"c8"),
  1134 => (x"4b",x"73",x"8b",x"c2"),
  1135 => (x"00",x"1c",x"e8",x"27"),
  1136 => (x"72",x"93",x"bf",x"00"),
  1137 => (x"27",x"82",x"73",x"4a"),
  1138 => (x"00",x"00",x"1c",x"ec"),
  1139 => (x"66",x"cc",x"4b",x"bf"),
  1140 => (x"4a",x"72",x"9b",x"bf"),
  1141 => (x"66",x"d0",x"82",x"73"),
  1142 => (x"27",x"1e",x"72",x"1e"),
  1143 => (x"00",x"00",x"08",x"6f"),
  1144 => (x"70",x"86",x"c8",x"0f"),
  1145 => (x"05",x"9a",x"72",x"4a"),
  1146 => (x"c0",x"87",x"c5",x"c0"),
  1147 => (x"87",x"c2",x"c0",x"48"),
  1148 => (x"4b",x"26",x"48",x"c1"),
  1149 => (x"4f",x"26",x"4a",x"26"),
  1150 => (x"5b",x"5a",x"5e",x"0e"),
  1151 => (x"d8",x"0e",x"5d",x"5c"),
  1152 => (x"66",x"d4",x"4c",x"66"),
  1153 => (x"1d",x"20",x"27",x"1e"),
  1154 => (x"27",x"1e",x"00",x"00"),
  1155 => (x"00",x"00",x"0f",x"f1"),
  1156 => (x"70",x"86",x"c8",x"0f"),
  1157 => (x"02",x"9a",x"72",x"4a"),
  1158 => (x"27",x"87",x"df",x"c1"),
  1159 => (x"00",x"00",x"1d",x"24"),
  1160 => (x"ff",x"c7",x"4a",x"bf"),
  1161 => (x"72",x"2a",x"c9",x"82"),
  1162 => (x"27",x"4b",x"c0",x"4d"),
  1163 => (x"00",x"00",x"12",x"9c"),
  1164 => (x"00",x"6e",x"27",x"1e"),
  1165 => (x"c4",x"0f",x"00",x"00"),
  1166 => (x"ad",x"b7",x"c0",x"86"),
  1167 => (x"87",x"d0",x"c1",x"06"),
  1168 => (x"20",x"27",x"1e",x"74"),
  1169 => (x"1e",x"00",x"00",x"1d"),
  1170 => (x"00",x"11",x"a5",x"27"),
  1171 => (x"86",x"c8",x"0f",x"00"),
  1172 => (x"9a",x"72",x"4a",x"70"),
  1173 => (x"87",x"c5",x"c0",x"05"),
  1174 => (x"f5",x"c0",x"48",x"c0"),
  1175 => (x"1d",x"20",x"27",x"87"),
  1176 => (x"27",x"1e",x"00",x"00"),
  1177 => (x"00",x"00",x"11",x"6b"),
  1178 => (x"c8",x"86",x"c4",x"0f"),
  1179 => (x"83",x"c1",x"84",x"c0"),
  1180 => (x"04",x"ab",x"b7",x"75"),
  1181 => (x"c0",x"87",x"c9",x"ff"),
  1182 => (x"66",x"d4",x"87",x"d6"),
  1183 => (x"12",x"b5",x"27",x"1e"),
  1184 => (x"27",x"1e",x"00",x"00"),
  1185 => (x"00",x"00",x"01",x"50"),
  1186 => (x"c0",x"86",x"c8",x"0f"),
  1187 => (x"87",x"c2",x"c0",x"48"),
  1188 => (x"4d",x"26",x"48",x"c1"),
  1189 => (x"4b",x"26",x"4c",x"26"),
  1190 => (x"4f",x"26",x"4a",x"26"),
  1191 => (x"6e",x"65",x"70",x"4f"),
  1192 => (x"66",x"20",x"64",x"65"),
  1193 => (x"2c",x"65",x"6c",x"69"),
  1194 => (x"61",x"6f",x"6c",x"20"),
  1195 => (x"67",x"6e",x"69",x"64"),
  1196 => (x"0a",x"2e",x"2e",x"2e"),
  1197 => (x"6e",x"61",x"43",x"00"),
  1198 => (x"6f",x"20",x"74",x"27"),
  1199 => (x"20",x"6e",x"65",x"70"),
  1200 => (x"00",x"0a",x"73",x"25"),
  1201 => (x"5b",x"5a",x"5e",x"0e"),
  1202 => (x"4a",x"66",x"cc",x"0e"),
  1203 => (x"ff",x"c3",x"2a",x"d8"),
  1204 => (x"4b",x"66",x"cc",x"9a"),
  1205 => (x"fc",x"cf",x"2b",x"c8"),
  1206 => (x"4a",x"72",x"9b",x"c0"),
  1207 => (x"66",x"cc",x"b2",x"73"),
  1208 => (x"c0",x"33",x"c8",x"4b"),
  1209 => (x"c0",x"c0",x"f0",x"ff"),
  1210 => (x"73",x"4a",x"72",x"9b"),
  1211 => (x"4b",x"66",x"cc",x"b2"),
  1212 => (x"c0",x"ff",x"33",x"d8"),
  1213 => (x"9b",x"c0",x"c0",x"c0"),
  1214 => (x"b2",x"73",x"4a",x"72"),
  1215 => (x"4b",x"26",x"48",x"72"),
  1216 => (x"4f",x"26",x"4a",x"26"),
  1217 => (x"5b",x"5a",x"5e",x"0e"),
  1218 => (x"4b",x"66",x"cc",x"0e"),
  1219 => (x"ff",x"c3",x"2b",x"c8"),
  1220 => (x"66",x"cc",x"4b",x"9b"),
  1221 => (x"cf",x"32",x"c8",x"4a"),
  1222 => (x"72",x"9a",x"c0",x"fc"),
  1223 => (x"4a",x"b2",x"73",x"4a"),
  1224 => (x"4b",x"26",x"48",x"72"),
  1225 => (x"4f",x"26",x"4a",x"26"),
  1226 => (x"5b",x"5a",x"5e",x"0e"),
  1227 => (x"4a",x"66",x"cc",x"0e"),
  1228 => (x"ff",x"cf",x"2a",x"d0"),
  1229 => (x"cc",x"4a",x"9a",x"ff"),
  1230 => (x"33",x"d0",x"4b",x"66"),
  1231 => (x"9b",x"c0",x"c0",x"f0"),
  1232 => (x"b2",x"73",x"4a",x"72"),
  1233 => (x"4b",x"26",x"48",x"72"),
  1234 => (x"4f",x"26",x"4a",x"26"),
  1235 => (x"87",x"fd",x"ff",x"1e"),
  1236 => (x"72",x"1e",x"4f",x"26"),
  1237 => (x"4a",x"66",x"cc",x"1e"),
  1238 => (x"c0",x"9a",x"df",x"c3"),
  1239 => (x"b7",x"c0",x"8a",x"f7"),
  1240 => (x"c3",x"c0",x"03",x"aa"),
  1241 => (x"82",x"e7",x"c0",x"87"),
  1242 => (x"c4",x"48",x"66",x"c8"),
  1243 => (x"58",x"a6",x"cc",x"30"),
  1244 => (x"72",x"48",x"66",x"c8"),
  1245 => (x"58",x"a6",x"cc",x"b0"),
  1246 => (x"26",x"48",x"66",x"c8"),
  1247 => (x"0e",x"4f",x"26",x"4a"),
  1248 => (x"5c",x"5b",x"5a",x"5e"),
  1249 => (x"1d",x"30",x"27",x"0e"),
  1250 => (x"48",x"bf",x"00",x"00"),
  1251 => (x"34",x"27",x"80",x"c1"),
  1252 => (x"58",x"00",x"00",x"1d"),
  1253 => (x"4a",x"66",x"d0",x"97"),
  1254 => (x"c0",x"c0",x"c0",x"c1"),
  1255 => (x"c0",x"c4",x"92",x"c0"),
  1256 => (x"c1",x"4a",x"92",x"b7"),
  1257 => (x"05",x"aa",x"b7",x"d3"),
  1258 => (x"27",x"87",x"e9",x"c0"),
  1259 => (x"00",x"00",x"1d",x"30"),
  1260 => (x"27",x"79",x"c0",x"49"),
  1261 => (x"00",x"00",x"1d",x"34"),
  1262 => (x"27",x"79",x"c0",x"49"),
  1263 => (x"00",x"00",x"1d",x"3c"),
  1264 => (x"27",x"79",x"c0",x"49"),
  1265 => (x"00",x"00",x"1d",x"40"),
  1266 => (x"ff",x"79",x"c0",x"49"),
  1267 => (x"d3",x"c1",x"49",x"c0"),
  1268 => (x"87",x"f6",x"c9",x"79"),
  1269 => (x"00",x"1d",x"30",x"27"),
  1270 => (x"c1",x"49",x"bf",x"00"),
  1271 => (x"c1",x"05",x"a9",x"b7"),
  1272 => (x"c0",x"ff",x"87",x"db"),
  1273 => (x"79",x"f4",x"c1",x"49"),
  1274 => (x"4a",x"66",x"d0",x"97"),
  1275 => (x"c0",x"c0",x"c0",x"c1"),
  1276 => (x"c0",x"c4",x"92",x"c0"),
  1277 => (x"72",x"4a",x"92",x"b7"),
  1278 => (x"1d",x"40",x"27",x"1e"),
  1279 => (x"1e",x"bf",x"00",x"00"),
  1280 => (x"00",x"13",x"52",x"27"),
  1281 => (x"86",x"c8",x"0f",x"00"),
  1282 => (x"00",x"1d",x"44",x"27"),
  1283 => (x"40",x"27",x"58",x"00"),
  1284 => (x"bf",x"00",x"00",x"1d"),
  1285 => (x"ac",x"b7",x"c3",x"4c"),
  1286 => (x"87",x"c6",x"c0",x"06"),
  1287 => (x"88",x"74",x"48",x"ca"),
  1288 => (x"4a",x"74",x"4c",x"70"),
  1289 => (x"48",x"72",x"82",x"c1"),
  1290 => (x"3c",x"27",x"30",x"c1"),
  1291 => (x"58",x"00",x"00",x"1d"),
  1292 => (x"f0",x"c0",x"48",x"74"),
  1293 => (x"49",x"c0",x"ff",x"80"),
  1294 => (x"cd",x"c8",x"79",x"70"),
  1295 => (x"1d",x"40",x"27",x"87"),
  1296 => (x"49",x"bf",x"00",x"00"),
  1297 => (x"01",x"a9",x"b7",x"c9"),
  1298 => (x"27",x"87",x"ff",x"c7"),
  1299 => (x"00",x"00",x"1d",x"40"),
  1300 => (x"b7",x"c0",x"49",x"bf"),
  1301 => (x"f1",x"c7",x"06",x"a9"),
  1302 => (x"1d",x"40",x"27",x"87"),
  1303 => (x"48",x"bf",x"00",x"00"),
  1304 => (x"ff",x"80",x"f0",x"c0"),
  1305 => (x"79",x"70",x"49",x"c0"),
  1306 => (x"00",x"1d",x"30",x"27"),
  1307 => (x"c3",x"49",x"bf",x"00"),
  1308 => (x"c0",x"01",x"a9",x"b7"),
  1309 => (x"d0",x"97",x"87",x"e9"),
  1310 => (x"c0",x"c1",x"4a",x"66"),
  1311 => (x"92",x"c0",x"c0",x"c0"),
  1312 => (x"92",x"b7",x"c0",x"c4"),
  1313 => (x"27",x"1e",x"72",x"4a"),
  1314 => (x"00",x"00",x"1d",x"3c"),
  1315 => (x"52",x"27",x"1e",x"bf"),
  1316 => (x"0f",x"00",x"00",x"13"),
  1317 => (x"40",x"27",x"86",x"c8"),
  1318 => (x"58",x"00",x"00",x"1d"),
  1319 => (x"27",x"87",x"eb",x"c6"),
  1320 => (x"00",x"00",x"1d",x"38"),
  1321 => (x"82",x"c3",x"4a",x"bf"),
  1322 => (x"00",x"1d",x"30",x"27"),
  1323 => (x"72",x"49",x"bf",x"00"),
  1324 => (x"c0",x"01",x"a9",x"b7"),
  1325 => (x"d0",x"97",x"87",x"f1"),
  1326 => (x"c0",x"c1",x"4a",x"66"),
  1327 => (x"92",x"c0",x"c0",x"c0"),
  1328 => (x"92",x"b7",x"c0",x"c4"),
  1329 => (x"27",x"1e",x"72",x"4a"),
  1330 => (x"00",x"00",x"1d",x"34"),
  1331 => (x"52",x"27",x"1e",x"bf"),
  1332 => (x"0f",x"00",x"00",x"13"),
  1333 => (x"38",x"27",x"86",x"c8"),
  1334 => (x"58",x"00",x"00",x"1d"),
  1335 => (x"00",x"1d",x"44",x"27"),
  1336 => (x"79",x"c1",x"49",x"00"),
  1337 => (x"27",x"87",x"e3",x"c5"),
  1338 => (x"00",x"00",x"1d",x"40"),
  1339 => (x"b7",x"c0",x"49",x"bf"),
  1340 => (x"d0",x"c3",x"06",x"a9"),
  1341 => (x"1d",x"40",x"27",x"87"),
  1342 => (x"49",x"bf",x"00",x"00"),
  1343 => (x"01",x"a9",x"b7",x"c3"),
  1344 => (x"27",x"87",x"c2",x"c3"),
  1345 => (x"00",x"00",x"1d",x"3c"),
  1346 => (x"32",x"c1",x"4a",x"bf"),
  1347 => (x"30",x"27",x"82",x"c1"),
  1348 => (x"bf",x"00",x"00",x"1d"),
  1349 => (x"a9",x"b7",x"72",x"49"),
  1350 => (x"87",x"c2",x"c2",x"01"),
  1351 => (x"4a",x"66",x"d0",x"97"),
  1352 => (x"c0",x"c0",x"c0",x"c1"),
  1353 => (x"c0",x"c4",x"92",x"c0"),
  1354 => (x"72",x"4a",x"92",x"b7"),
  1355 => (x"1d",x"48",x"27",x"1e"),
  1356 => (x"1e",x"bf",x"00",x"00"),
  1357 => (x"00",x"13",x"52",x"27"),
  1358 => (x"86",x"c8",x"0f",x"00"),
  1359 => (x"00",x"1d",x"4c",x"27"),
  1360 => (x"44",x"27",x"58",x"00"),
  1361 => (x"bf",x"00",x"00",x"1d"),
  1362 => (x"27",x"8a",x"c1",x"4a"),
  1363 => (x"00",x"00",x"1d",x"44"),
  1364 => (x"c0",x"79",x"72",x"49"),
  1365 => (x"c3",x"03",x"aa",x"b7"),
  1366 => (x"34",x"27",x"87",x"f0"),
  1367 => (x"bf",x"00",x"00",x"1d"),
  1368 => (x"1d",x"48",x"27",x"4a"),
  1369 => (x"bf",x"97",x"00",x"00"),
  1370 => (x"1d",x"34",x"27",x"52"),
  1371 => (x"4a",x"bf",x"00",x"00"),
  1372 => (x"34",x"27",x"82",x"c1"),
  1373 => (x"49",x"00",x"00",x"1d"),
  1374 => (x"4c",x"27",x"79",x"72"),
  1375 => (x"bf",x"00",x"00",x"1d"),
  1376 => (x"c0",x"06",x"aa",x"b7"),
  1377 => (x"4c",x"27",x"87",x"cd"),
  1378 => (x"49",x"00",x"00",x"1d"),
  1379 => (x"00",x"1d",x"34",x"27"),
  1380 => (x"27",x"79",x"bf",x"00"),
  1381 => (x"00",x"00",x"1d",x"44"),
  1382 => (x"c2",x"79",x"c1",x"49"),
  1383 => (x"44",x"27",x"87",x"ec"),
  1384 => (x"bf",x"00",x"00",x"1d"),
  1385 => (x"87",x"e2",x"c2",x"05"),
  1386 => (x"00",x"1d",x"48",x"27"),
  1387 => (x"c4",x"4b",x"bf",x"00"),
  1388 => (x"1d",x"48",x"27",x"33"),
  1389 => (x"73",x"49",x"00",x"00"),
  1390 => (x"1d",x"34",x"27",x"79"),
  1391 => (x"4a",x"bf",x"00",x"00"),
  1392 => (x"c5",x"c2",x"52",x"73"),
  1393 => (x"1d",x"40",x"27",x"87"),
  1394 => (x"49",x"bf",x"00",x"00"),
  1395 => (x"04",x"a9",x"b7",x"c7"),
  1396 => (x"c0",x"87",x"e8",x"c1"),
  1397 => (x"49",x"f4",x"fe",x"4b"),
  1398 => (x"34",x"27",x"79",x"c1"),
  1399 => (x"49",x"00",x"00",x"1d"),
  1400 => (x"4c",x"27",x"79",x"c0"),
  1401 => (x"bf",x"00",x"00",x"1d"),
  1402 => (x"a9",x"b7",x"c0",x"49"),
  1403 => (x"87",x"e5",x"c0",x"06"),
  1404 => (x"00",x"1d",x"34",x"27"),
  1405 => (x"83",x"bf",x"bf",x"00"),
  1406 => (x"00",x"1d",x"34",x"27"),
  1407 => (x"c4",x"4a",x"bf",x"00"),
  1408 => (x"1d",x"34",x"27",x"82"),
  1409 => (x"72",x"49",x"00",x"00"),
  1410 => (x"1d",x"4c",x"27",x"79"),
  1411 => (x"b7",x"bf",x"00",x"00"),
  1412 => (x"db",x"ff",x"04",x"aa"),
  1413 => (x"27",x"1e",x"73",x"87"),
  1414 => (x"00",x"00",x"1d",x"4c"),
  1415 => (x"34",x"27",x"1e",x"bf"),
  1416 => (x"1e",x"00",x"00",x"1a"),
  1417 => (x"00",x"01",x"50",x"27"),
  1418 => (x"86",x"cc",x"0f",x"00"),
  1419 => (x"c1",x"49",x"c0",x"ff"),
  1420 => (x"4c",x"27",x"79",x"c2"),
  1421 => (x"0f",x"00",x"00",x"13"),
  1422 => (x"27",x"87",x"cf",x"c0"),
  1423 => (x"00",x"00",x"1d",x"40"),
  1424 => (x"f0",x"c0",x"48",x"bf"),
  1425 => (x"49",x"c0",x"ff",x"80"),
  1426 => (x"4c",x"26",x"79",x"70"),
  1427 => (x"4a",x"26",x"4b",x"26"),
  1428 => (x"ff",x"1e",x"4f",x"26"),
  1429 => (x"4f",x"26",x"87",x"fd"),
  1430 => (x"5b",x"5a",x"5e",x"0e"),
  1431 => (x"27",x"0e",x"5d",x"5c"),
  1432 => (x"00",x"00",x"18",x"40"),
  1433 => (x"00",x"6e",x"27",x"1e"),
  1434 => (x"c4",x"0f",x"00",x"00"),
  1435 => (x"05",x"78",x"27",x"86"),
  1436 => (x"70",x"0f",x"00",x"00"),
  1437 => (x"02",x"9a",x"72",x"4a"),
  1438 => (x"27",x"87",x"ce",x"c4"),
  1439 => (x"00",x"00",x"18",x"1d"),
  1440 => (x"00",x"6e",x"27",x"1e"),
  1441 => (x"c4",x"0f",x"00",x"00"),
  1442 => (x"0b",x"39",x"27",x"86"),
  1443 => (x"27",x"0f",x"00",x"00"),
  1444 => (x"00",x"00",x"1d",x"50"),
  1445 => (x"18",x"34",x"27",x"1e"),
  1446 => (x"27",x"1e",x"00",x"00"),
  1447 => (x"00",x"00",x"11",x"f8"),
  1448 => (x"70",x"86",x"c8",x"0f"),
  1449 => (x"02",x"9a",x"72",x"4a"),
  1450 => (x"27",x"87",x"d0",x"c3"),
  1451 => (x"00",x"00",x"1d",x"50"),
  1452 => (x"17",x"f2",x"27",x"4b"),
  1453 => (x"27",x"1e",x"00",x"00"),
  1454 => (x"00",x"00",x"00",x"6e"),
  1455 => (x"c0",x"86",x"c4",x"0f"),
  1456 => (x"74",x"4c",x"13",x"4d"),
  1457 => (x"b7",x"e0",x"c0",x"4a"),
  1458 => (x"ed",x"c1",x"02",x"aa"),
  1459 => (x"ff",x"48",x"74",x"87"),
  1460 => (x"79",x"70",x"49",x"c0"),
  1461 => (x"e3",x"c0",x"4a",x"74"),
  1462 => (x"c1",x"02",x"aa",x"b7"),
  1463 => (x"4a",x"74",x"87",x"dc"),
  1464 => (x"aa",x"b7",x"c7",x"c1"),
  1465 => (x"87",x"c6",x"c0",x"05"),
  1466 => (x"00",x"13",x"4c",x"27"),
  1467 => (x"4a",x"74",x"0f",x"00"),
  1468 => (x"05",x"aa",x"b7",x"ca"),
  1469 => (x"27",x"87",x"c6",x"c0"),
  1470 => (x"00",x"00",x"16",x"52"),
  1471 => (x"c1",x"4a",x"74",x"0f"),
  1472 => (x"05",x"aa",x"b7",x"cc"),
  1473 => (x"27",x"87",x"c6",x"c0"),
  1474 => (x"00",x"00",x"1d",x"50"),
  1475 => (x"ff",x"4a",x"74",x"4b"),
  1476 => (x"8a",x"d0",x"9a",x"df"),
  1477 => (x"4a",x"74",x"4c",x"72"),
  1478 => (x"aa",x"b7",x"f9",x"c0"),
  1479 => (x"87",x"c6",x"c0",x"04"),
  1480 => (x"8a",x"d1",x"4a",x"74"),
  1481 => (x"35",x"c4",x"4c",x"72"),
  1482 => (x"4d",x"75",x"4a",x"74"),
  1483 => (x"4c",x"13",x"b5",x"72"),
  1484 => (x"e0",x"c0",x"4a",x"74"),
  1485 => (x"fe",x"05",x"aa",x"b7"),
  1486 => (x"4a",x"74",x"87",x"d3"),
  1487 => (x"aa",x"b7",x"e3",x"c0"),
  1488 => (x"87",x"e2",x"c0",x"02"),
  1489 => (x"e0",x"c0",x"4a",x"13"),
  1490 => (x"c0",x"05",x"aa",x"b7"),
  1491 => (x"4a",x"13",x"87",x"ca"),
  1492 => (x"aa",x"b7",x"e0",x"c0"),
  1493 => (x"87",x"f6",x"ff",x"02"),
  1494 => (x"1e",x"75",x"8b",x"c1"),
  1495 => (x"f8",x"27",x"1e",x"73"),
  1496 => (x"0f",x"00",x"00",x"11"),
  1497 => (x"4a",x"13",x"86",x"c8"),
  1498 => (x"02",x"aa",x"b7",x"ca"),
  1499 => (x"13",x"87",x"d0",x"fd"),
  1500 => (x"aa",x"b7",x"ca",x"4a"),
  1501 => (x"87",x"f7",x"ff",x"05"),
  1502 => (x"27",x"87",x"c4",x"fd"),
  1503 => (x"00",x"00",x"18",x"04"),
  1504 => (x"00",x"6e",x"27",x"1e"),
  1505 => (x"c4",x"0f",x"00",x"00"),
  1506 => (x"18",x"56",x"27",x"86"),
  1507 => (x"27",x"1e",x"00",x"00"),
  1508 => (x"00",x"00",x"00",x"6e"),
  1509 => (x"27",x"86",x"c4",x"0f"),
  1510 => (x"00",x"00",x"1d",x"4c"),
  1511 => (x"c3",x"79",x"c0",x"49"),
  1512 => (x"4d",x"ff",x"c8",x"f4"),
  1513 => (x"27",x"1e",x"ee",x"c0"),
  1514 => (x"00",x"00",x"00",x"4f"),
  1515 => (x"75",x"86",x"c4",x"0f"),
  1516 => (x"c9",x"f4",x"c3",x"4b"),
  1517 => (x"c0",x"ff",x"4d",x"c0"),
  1518 => (x"4a",x"74",x"4c",x"bf"),
  1519 => (x"72",x"9a",x"c0",x"c8"),
  1520 => (x"d1",x"c0",x"02",x"9a"),
  1521 => (x"c3",x"4a",x"74",x"87"),
  1522 => (x"1e",x"72",x"9a",x"ff"),
  1523 => (x"00",x"13",x"7f",x"27"),
  1524 => (x"86",x"c4",x"0f",x"00"),
  1525 => (x"4a",x"73",x"4b",x"75"),
  1526 => (x"9a",x"72",x"8b",x"c1"),
  1527 => (x"87",x"d6",x"ff",x"05"),
  1528 => (x"ff",x"c8",x"f4",x"c3"),
  1529 => (x"87",x"fc",x"fe",x"4d"),
  1530 => (x"4c",x"26",x"4d",x"26"),
  1531 => (x"4a",x"26",x"4b",x"26"),
  1532 => (x"61",x"50",x"4f",x"26"),
  1533 => (x"6e",x"69",x"73",x"72"),
  1534 => (x"61",x"6d",x"20",x"67"),
  1535 => (x"65",x"66",x"69",x"6e"),
  1536 => (x"00",x"0a",x"74",x"73"),
  1537 => (x"64",x"61",x"6f",x"4c"),
  1538 => (x"20",x"67",x"6e",x"69"),
  1539 => (x"69",x"6e",x"61",x"6d"),
  1540 => (x"74",x"73",x"65",x"66"),
  1541 => (x"69",x"61",x"66",x"20"),
  1542 => (x"0a",x"64",x"65",x"6c"),
  1543 => (x"6e",x"75",x"48",x"00"),
  1544 => (x"67",x"6e",x"69",x"74"),
  1545 => (x"72",x"6f",x"66",x"20"),
  1546 => (x"72",x"61",x"70",x"20"),
  1547 => (x"69",x"74",x"69",x"74"),
  1548 => (x"00",x"0a",x"6e",x"6f"),
  1549 => (x"49",x"4e",x"41",x"4d"),
  1550 => (x"54",x"53",x"45",x"46"),
  1551 => (x"00",x"54",x"53",x"4d"),
  1552 => (x"74",x"69",x"6e",x"49"),
  1553 => (x"69",x"6c",x"61",x"69"),
  1554 => (x"67",x"6e",x"69",x"7a"),
  1555 => (x"20",x"44",x"53",x"20"),
  1556 => (x"64",x"72",x"61",x"63"),
  1557 => (x"6f",x"42",x"00",x"0a"),
  1558 => (x"6e",x"69",x"74",x"6f"),
  1559 => (x"72",x"66",x"20",x"67"),
  1560 => (x"52",x"20",x"6d",x"6f"),
  1561 => (x"32",x"33",x"32",x"53"),
  1562 => (x"73",x"1e",x"00",x"2e"),
  1563 => (x"02",x"9a",x"72",x"1e"),
  1564 => (x"48",x"c0",x"87",x"d9"),
  1565 => (x"a9",x"72",x"4b",x"c1"),
  1566 => (x"83",x"73",x"82",x"01"),
  1567 => (x"a9",x"72",x"87",x"f8"),
  1568 => (x"80",x"73",x"89",x"03"),
  1569 => (x"2b",x"2a",x"c1",x"07"),
  1570 => (x"26",x"87",x"f3",x"05"),
  1571 => (x"1e",x"4f",x"26",x"4b"),
  1572 => (x"4d",x"c0",x"1e",x"75"),
  1573 => (x"ff",x"04",x"a1",x"71"),
  1574 => (x"bd",x"81",x"c1",x"b9"),
  1575 => (x"04",x"a2",x"72",x"07"),
  1576 => (x"82",x"c1",x"ba",x"ff"),
  1577 => (x"87",x"c2",x"07",x"bd"),
  1578 => (x"ff",x"05",x"9d",x"75"),
  1579 => (x"07",x"80",x"c1",x"b8"),
  1580 => (x"4f",x"26",x"4d",x"25"),
  1581 => (x"33",x"32",x"31",x"30"),
  1582 => (x"37",x"36",x"35",x"34"),
  1583 => (x"42",x"41",x"39",x"38"),
  1584 => (x"46",x"45",x"44",x"43"),
  1585 => (x"44",x"4d",x"43",x"00"),
  1586 => (x"61",x"65",x"52",x"00"),
  1587 => (x"66",x"6f",x"20",x"64"),
  1588 => (x"52",x"42",x"4d",x"20"),
  1589 => (x"69",x"61",x"66",x"20"),
  1590 => (x"0a",x"64",x"65",x"6c"),
  1591 => (x"20",x"6f",x"4e",x"00"),
  1592 => (x"74",x"72",x"61",x"70"),
  1593 => (x"6f",x"69",x"74",x"69"),
  1594 => (x"69",x"73",x"20",x"6e"),
  1595 => (x"74",x"61",x"6e",x"67"),
  1596 => (x"20",x"65",x"72",x"75"),
  1597 => (x"6e",x"75",x"6f",x"66"),
  1598 => (x"4d",x"00",x"0a",x"64"),
  1599 => (x"69",x"73",x"52",x"42"),
  1600 => (x"20",x"3a",x"65",x"7a"),
  1601 => (x"20",x"2c",x"64",x"25"),
  1602 => (x"74",x"72",x"61",x"70"),
  1603 => (x"6f",x"69",x"74",x"69"),
  1604 => (x"7a",x"69",x"73",x"6e"),
  1605 => (x"25",x"20",x"3a",x"65"),
  1606 => (x"6f",x"20",x"2c",x"64"),
  1607 => (x"65",x"73",x"66",x"66"),
  1608 => (x"66",x"6f",x"20",x"74"),
  1609 => (x"67",x"69",x"73",x"20"),
  1610 => (x"64",x"25",x"20",x"3a"),
  1611 => (x"69",x"73",x"20",x"2c"),
  1612 => (x"78",x"30",x"20",x"67"),
  1613 => (x"00",x"0a",x"78",x"25"),
  1614 => (x"64",x"61",x"65",x"52"),
  1615 => (x"20",x"67",x"6e",x"69"),
  1616 => (x"74",x"6f",x"6f",x"62"),
  1617 => (x"63",x"65",x"73",x"20"),
  1618 => (x"20",x"72",x"6f",x"74"),
  1619 => (x"00",x"0a",x"64",x"25"),
  1620 => (x"64",x"61",x"65",x"52"),
  1621 => (x"6f",x"6f",x"62",x"20"),
  1622 => (x"65",x"73",x"20",x"74"),
  1623 => (x"72",x"6f",x"74",x"63"),
  1624 => (x"6f",x"72",x"66",x"20"),
  1625 => (x"69",x"66",x"20",x"6d"),
  1626 => (x"20",x"74",x"73",x"72"),
  1627 => (x"74",x"72",x"61",x"70"),
  1628 => (x"6f",x"69",x"74",x"69"),
  1629 => (x"55",x"00",x"0a",x"6e"),
  1630 => (x"70",x"75",x"73",x"6e"),
  1631 => (x"74",x"72",x"6f",x"70"),
  1632 => (x"70",x"20",x"64",x"65"),
  1633 => (x"69",x"74",x"72",x"61"),
  1634 => (x"6e",x"6f",x"69",x"74"),
  1635 => (x"70",x"79",x"74",x"20"),
  1636 => (x"00",x"0d",x"21",x"65"),
  1637 => (x"33",x"54",x"41",x"46"),
  1638 => (x"20",x"20",x"20",x"32"),
  1639 => (x"61",x"65",x"52",x"00"),
  1640 => (x"67",x"6e",x"69",x"64"),
  1641 => (x"52",x"42",x"4d",x"20"),
  1642 => (x"42",x"4d",x"00",x"0a"),
  1643 => (x"75",x"73",x"20",x"52"),
  1644 => (x"73",x"65",x"63",x"63"),
  1645 => (x"6c",x"75",x"66",x"73"),
  1646 => (x"72",x"20",x"79",x"6c"),
  1647 => (x"0a",x"64",x"61",x"65"),
  1648 => (x"54",x"41",x"46",x"00"),
  1649 => (x"20",x"20",x"36",x"31"),
  1650 => (x"41",x"46",x"00",x"20"),
  1651 => (x"20",x"32",x"33",x"54"),
  1652 => (x"50",x"00",x"20",x"20"),
  1653 => (x"69",x"74",x"72",x"61"),
  1654 => (x"6e",x"6f",x"69",x"74"),
  1655 => (x"6e",x"75",x"6f",x"63"),
  1656 => (x"64",x"25",x"20",x"74"),
  1657 => (x"75",x"48",x"00",x"0a"),
  1658 => (x"6e",x"69",x"74",x"6e"),
  1659 => (x"6f",x"66",x"20",x"67"),
  1660 => (x"69",x"66",x"20",x"72"),
  1661 => (x"79",x"73",x"65",x"6c"),
  1662 => (x"6d",x"65",x"74",x"73"),
  1663 => (x"41",x"46",x"00",x"0a"),
  1664 => (x"20",x"32",x"33",x"54"),
  1665 => (x"46",x"00",x"20",x"20"),
  1666 => (x"36",x"31",x"54",x"41"),
  1667 => (x"00",x"20",x"20",x"20"),
  1668 => (x"73",x"75",x"6c",x"43"),
  1669 => (x"20",x"72",x"65",x"74"),
  1670 => (x"65",x"7a",x"69",x"73"),
  1671 => (x"64",x"25",x"20",x"3a"),
  1672 => (x"6c",x"43",x"20",x"2c"),
  1673 => (x"65",x"74",x"73",x"75"),
  1674 => (x"61",x"6d",x"20",x"72"),
  1675 => (x"20",x"2c",x"6b",x"73"),
  1676 => (x"00",x"0a",x"64",x"25"),
  1677 => (x"63",x"65",x"68",x"43"),
  1678 => (x"6d",x"75",x"73",x"6b"),
  1679 => (x"20",x"6f",x"74",x"20"),
  1680 => (x"20",x"3a",x"64",x"25"),
  1681 => (x"00",x"0a",x"64",x"25"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
