
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"2c",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"29"),
    10 => (x"87",x"fd",x"00",x"4f"),
    11 => (x"d8",x"f2",x"c3",x"4f"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"d8",x"f2",x"c3"),
    14 => (x"48",x"e0",x"cf",x"c1"),
    15 => (x"03",x"89",x"d0",x"89"),
    16 => (x"40",x"40",x"40",x"c0"),
    17 => (x"d0",x"87",x"f6",x"40"),
    18 => (x"50",x"c0",x"05",x"81"),
    19 => (x"f9",x"05",x"89",x"c1"),
    20 => (x"df",x"cf",x"c1",x"87"),
    21 => (x"df",x"cf",x"c1",x"4d"),
    22 => (x"02",x"ad",x"74",x"4c"),
    23 => (x"0f",x"24",x"87",x"c4"),
    24 => (x"e0",x"cb",x"87",x"f7"),
    25 => (x"df",x"cf",x"c1",x"87"),
    26 => (x"df",x"cf",x"c1",x"4d"),
    27 => (x"02",x"ad",x"74",x"4c"),
    28 => (x"8c",x"c4",x"87",x"c6"),
    29 => (x"87",x"f5",x"0f",x"6c"),
    30 => (x"1e",x"87",x"fd",x"00"),
    31 => (x"1e",x"74",x"1e",x"73"),
    32 => (x"66",x"d0",x"1e",x"75"),
    33 => (x"e0",x"cf",x"c1",x"4a"),
    34 => (x"4d",x"ef",x"c3",x"4b"),
    35 => (x"9a",x"72",x"4c",x"c0"),
    36 => (x"c0",x"87",x"c6",x"05"),
    37 => (x"eb",x"c0",x"53",x"f0"),
    38 => (x"02",x"9a",x"72",x"87"),
    39 => (x"72",x"87",x"e5",x"c0"),
    40 => (x"d8",x"49",x"72",x"1e"),
    41 => (x"e6",x"c8",x"4a",x"66"),
    42 => (x"75",x"4a",x"26",x"87"),
    43 => (x"53",x"11",x"49",x"a1"),
    44 => (x"49",x"72",x"1e",x"71"),
    45 => (x"c8",x"4a",x"66",x"d8"),
    46 => (x"4a",x"70",x"87",x"d5"),
    47 => (x"9a",x"72",x"49",x"26"),
    48 => (x"87",x"db",x"ff",x"05"),
    49 => (x"ab",x"e0",x"cf",x"c1"),
    50 => (x"d8",x"87",x"da",x"02"),
    51 => (x"66",x"dc",x"4d",x"66"),
    52 => (x"97",x"8b",x"c1",x"1e"),
    53 => (x"1e",x"71",x"49",x"6b"),
    54 => (x"86",x"c8",x"0f",x"75"),
    55 => (x"cf",x"c1",x"84",x"c1"),
    56 => (x"e9",x"05",x"ab",x"e0"),
    57 => (x"26",x"48",x"74",x"87"),
    58 => (x"26",x"4c",x"26",x"4d"),
    59 => (x"30",x"4f",x"26",x"4b"),
    60 => (x"34",x"33",x"32",x"31"),
    61 => (x"38",x"37",x"36",x"35"),
    62 => (x"43",x"42",x"41",x"39"),
    63 => (x"00",x"46",x"45",x"44"),
    64 => (x"74",x"1e",x"73",x"1e"),
    65 => (x"d0",x"1e",x"75",x"1e"),
    66 => (x"4d",x"ff",x"4c",x"66"),
    67 => (x"9b",x"73",x"4b",x"14"),
    68 => (x"c1",x"87",x"d8",x"02"),
    69 => (x"1e",x"66",x"d8",x"85"),
    70 => (x"66",x"dc",x"1e",x"73"),
    71 => (x"73",x"86",x"c8",x"0f"),
    72 => (x"87",x"c7",x"05",x"a8"),
    73 => (x"9b",x"73",x"4b",x"14"),
    74 => (x"75",x"87",x"e8",x"05"),
    75 => (x"26",x"4d",x"26",x"48"),
    76 => (x"26",x"4b",x"26",x"4c"),
    77 => (x"1e",x"73",x"1e",x"4f"),
    78 => (x"1e",x"75",x"1e",x"74"),
    79 => (x"e4",x"c0",x"86",x"f4"),
    80 => (x"4d",x"c0",x"4c",x"66"),
    81 => (x"c0",x"48",x"a6",x"c4"),
    82 => (x"97",x"66",x"dc",x"78"),
    83 => (x"66",x"dc",x"4b",x"bf"),
    84 => (x"c0",x"80",x"c1",x"48"),
    85 => (x"73",x"58",x"a6",x"e0"),
    86 => (x"f9",x"c4",x"02",x"9b"),
    87 => (x"02",x"66",x"c4",x"87"),
    88 => (x"c8",x"87",x"c8",x"c4"),
    89 => (x"78",x"c0",x"48",x"a6"),
    90 => (x"78",x"c0",x"80",x"fc"),
    91 => (x"f0",x"c0",x"49",x"73"),
    92 => (x"e5",x"c1",x"02",x"ab"),
    93 => (x"a9",x"e3",x"c1",x"87"),
    94 => (x"87",x"e6",x"c1",x"02"),
    95 => (x"02",x"a9",x"e4",x"c1"),
    96 => (x"c1",x"87",x"e2",x"c0"),
    97 => (x"c1",x"02",x"a9",x"ec"),
    98 => (x"f0",x"c1",x"87",x"d0"),
    99 => (x"87",x"dd",x"02",x"a9"),
   100 => (x"02",x"a9",x"f3",x"c1"),
   101 => (x"f5",x"c1",x"87",x"df"),
   102 => (x"87",x"c9",x"02",x"a9"),
   103 => (x"02",x"a9",x"f8",x"c1"),
   104 => (x"db",x"c1",x"87",x"cb"),
   105 => (x"48",x"a6",x"c8",x"87"),
   106 => (x"f0",x"c1",x"78",x"ca"),
   107 => (x"48",x"a6",x"c8",x"87"),
   108 => (x"e8",x"c1",x"78",x"d0"),
   109 => (x"66",x"e8",x"c0",x"87"),
   110 => (x"c0",x"1e",x"74",x"1e"),
   111 => (x"c4",x"48",x"66",x"e8"),
   112 => (x"a6",x"ec",x"c0",x"80"),
   113 => (x"66",x"e8",x"c0",x"58"),
   114 => (x"69",x"89",x"c4",x"49"),
   115 => (x"87",x"f0",x"fc",x"1e"),
   116 => (x"49",x"70",x"86",x"cc"),
   117 => (x"c1",x"4d",x"a5",x"71"),
   118 => (x"a6",x"c4",x"87",x"c3"),
   119 => (x"c0",x"78",x"c1",x"48"),
   120 => (x"e8",x"c0",x"87",x"fb"),
   121 => (x"e4",x"c0",x"1e",x"66"),
   122 => (x"80",x"c4",x"48",x"66"),
   123 => (x"58",x"a6",x"e8",x"c0"),
   124 => (x"49",x"66",x"e4",x"c0"),
   125 => (x"1e",x"69",x"89",x"c4"),
   126 => (x"86",x"c8",x"0f",x"74"),
   127 => (x"87",x"dd",x"85",x"c1"),
   128 => (x"02",x"ab",x"e5",x"c0"),
   129 => (x"e8",x"c0",x"87",x"cb"),
   130 => (x"e5",x"c0",x"1e",x"66"),
   131 => (x"c8",x"0f",x"74",x"1e"),
   132 => (x"66",x"e8",x"c0",x"86"),
   133 => (x"74",x"1e",x"73",x"1e"),
   134 => (x"c1",x"86",x"c8",x"0f"),
   135 => (x"02",x"66",x"c8",x"85"),
   136 => (x"c0",x"87",x"df",x"c1"),
   137 => (x"c4",x"48",x"66",x"e0"),
   138 => (x"a6",x"e4",x"c0",x"80"),
   139 => (x"66",x"e0",x"c0",x"58"),
   140 => (x"69",x"89",x"c4",x"49"),
   141 => (x"ab",x"e4",x"c1",x"7e"),
   142 => (x"6e",x"87",x"d8",x"05"),
   143 => (x"a8",x"b7",x"c0",x"48"),
   144 => (x"c0",x"87",x"d0",x"03"),
   145 => (x"ec",x"c1",x"1e",x"ed"),
   146 => (x"6e",x"86",x"c4",x"87"),
   147 => (x"88",x"08",x"c0",x"48"),
   148 => (x"c0",x"58",x"a6",x"c4"),
   149 => (x"74",x"1e",x"66",x"e8"),
   150 => (x"1e",x"66",x"d0",x"1e"),
   151 => (x"f8",x"1e",x"66",x"cc"),
   152 => (x"86",x"d0",x"87",x"d9"),
   153 => (x"a5",x"71",x"49",x"70"),
   154 => (x"c0",x"87",x"d7",x"4d"),
   155 => (x"c7",x"05",x"ab",x"e5"),
   156 => (x"48",x"a6",x"c4",x"87"),
   157 => (x"87",x"ca",x"78",x"c1"),
   158 => (x"1e",x"66",x"e8",x"c0"),
   159 => (x"0f",x"74",x"1e",x"73"),
   160 => (x"66",x"dc",x"86",x"c8"),
   161 => (x"dc",x"4b",x"bf",x"97"),
   162 => (x"80",x"c1",x"48",x"66"),
   163 => (x"58",x"a6",x"e0",x"c0"),
   164 => (x"fb",x"05",x"9b",x"73"),
   165 => (x"48",x"75",x"87",x"c7"),
   166 => (x"4d",x"26",x"8e",x"f4"),
   167 => (x"4b",x"26",x"4c",x"26"),
   168 => (x"c0",x"1e",x"4f",x"26"),
   169 => (x"1e",x"f5",x"ca",x"1e"),
   170 => (x"d0",x"1e",x"a6",x"d0"),
   171 => (x"c4",x"fa",x"1e",x"66"),
   172 => (x"26",x"86",x"d0",x"87"),
   173 => (x"86",x"fc",x"1e",x"4f"),
   174 => (x"69",x"49",x"c0",x"ff"),
   175 => (x"98",x"c0",x"c4",x"48"),
   176 => (x"6e",x"58",x"a6",x"c4"),
   177 => (x"c8",x"87",x"f4",x"02"),
   178 => (x"fc",x"48",x"79",x"66"),
   179 => (x"1e",x"4f",x"26",x"8e"),
   180 => (x"9a",x"72",x"1e",x"73"),
   181 => (x"87",x"e7",x"c0",x"02"),
   182 => (x"4b",x"c1",x"48",x"c0"),
   183 => (x"d1",x"06",x"a9",x"72"),
   184 => (x"06",x"82",x"72",x"87"),
   185 => (x"83",x"73",x"87",x"c9"),
   186 => (x"f4",x"01",x"a9",x"72"),
   187 => (x"c1",x"87",x"c3",x"87"),
   188 => (x"a9",x"72",x"3a",x"b2"),
   189 => (x"80",x"73",x"89",x"03"),
   190 => (x"2b",x"2a",x"c1",x"07"),
   191 => (x"26",x"87",x"f3",x"05"),
   192 => (x"1e",x"4f",x"26",x"4b"),
   193 => (x"4d",x"c4",x"1e",x"75"),
   194 => (x"04",x"a1",x"b7",x"71"),
   195 => (x"81",x"c1",x"b9",x"ff"),
   196 => (x"72",x"07",x"bd",x"c3"),
   197 => (x"ff",x"04",x"a2",x"b7"),
   198 => (x"c1",x"82",x"c1",x"ba"),
   199 => (x"ee",x"fe",x"07",x"bd"),
   200 => (x"04",x"2d",x"c1",x"87"),
   201 => (x"80",x"c1",x"b8",x"ff"),
   202 => (x"ff",x"04",x"2d",x"07"),
   203 => (x"07",x"81",x"c1",x"b9"),
   204 => (x"4f",x"26",x"4d",x"26"),
   205 => (x"12",x"1e",x"72",x"1e"),
   206 => (x"c4",x"02",x"11",x"48"),
   207 => (x"f6",x"02",x"88",x"87"),
   208 => (x"26",x"4a",x"26",x"87"),
   209 => (x"1e",x"73",x"1e",x"4f"),
   210 => (x"1e",x"75",x"1e",x"74"),
   211 => (x"c1",x"86",x"dc",x"ff"),
   212 => (x"c3",x"48",x"f4",x"cf"),
   213 => (x"c1",x"78",x"f8",x"ef"),
   214 => (x"c3",x"48",x"f0",x"cf"),
   215 => (x"48",x"78",x"e8",x"f0"),
   216 => (x"78",x"f8",x"ef",x"c3"),
   217 => (x"48",x"ec",x"f0",x"c3"),
   218 => (x"80",x"c4",x"78",x"c0"),
   219 => (x"f0",x"c3",x"78",x"c2"),
   220 => (x"e8",x"c0",x"48",x"f4"),
   221 => (x"c3",x"1e",x"71",x"78"),
   222 => (x"c0",x"49",x"f8",x"f0"),
   223 => (x"20",x"48",x"c8",x"ee"),
   224 => (x"20",x"41",x"20",x"41"),
   225 => (x"20",x"41",x"20",x"41"),
   226 => (x"20",x"41",x"20",x"41"),
   227 => (x"10",x"51",x"10",x"41"),
   228 => (x"26",x"51",x"10",x"51"),
   229 => (x"c3",x"1e",x"71",x"49"),
   230 => (x"c0",x"49",x"d8",x"f1"),
   231 => (x"20",x"48",x"e8",x"ee"),
   232 => (x"20",x"41",x"20",x"41"),
   233 => (x"20",x"41",x"20",x"41"),
   234 => (x"20",x"41",x"20",x"41"),
   235 => (x"10",x"51",x"10",x"41"),
   236 => (x"26",x"51",x"10",x"51"),
   237 => (x"ec",x"ec",x"c1",x"49"),
   238 => (x"c0",x"78",x"ca",x"48"),
   239 => (x"fb",x"1e",x"c8",x"ef"),
   240 => (x"86",x"c4",x"87",x"e0"),
   241 => (x"1e",x"cc",x"ef",x"c0"),
   242 => (x"c4",x"87",x"d7",x"fb"),
   243 => (x"fc",x"ef",x"c0",x"86"),
   244 => (x"87",x"ce",x"fb",x"1e"),
   245 => (x"e7",x"c0",x"86",x"c4"),
   246 => (x"d4",x"02",x"bf",x"ec"),
   247 => (x"f4",x"e7",x"c0",x"87"),
   248 => (x"87",x"fe",x"fa",x"1e"),
   249 => (x"e8",x"c0",x"86",x"c4"),
   250 => (x"f5",x"fa",x"1e",x"e0"),
   251 => (x"d2",x"86",x"c4",x"87"),
   252 => (x"e4",x"e8",x"c0",x"87"),
   253 => (x"87",x"ea",x"fa",x"1e"),
   254 => (x"e9",x"c0",x"86",x"c4"),
   255 => (x"e1",x"fa",x"1e",x"d4"),
   256 => (x"c0",x"86",x"c4",x"87"),
   257 => (x"1e",x"bf",x"f0",x"e7"),
   258 => (x"1e",x"c0",x"f0",x"c0"),
   259 => (x"c8",x"87",x"d3",x"fa"),
   260 => (x"e0",x"ef",x"c3",x"86"),
   261 => (x"bf",x"c8",x"ff",x"48"),
   262 => (x"48",x"a6",x"c8",x"78"),
   263 => (x"e7",x"c0",x"78",x"c1"),
   264 => (x"c0",x"48",x"bf",x"f0"),
   265 => (x"c8",x"06",x"a8",x"b7"),
   266 => (x"a6",x"cc",x"87",x"f5"),
   267 => (x"58",x"a6",x"d4",x"48"),
   268 => (x"a6",x"dc",x"80",x"c8"),
   269 => (x"48",x"a6",x"dc",x"58"),
   270 => (x"c1",x"58",x"a6",x"c8"),
   271 => (x"c1",x"48",x"c0",x"d0"),
   272 => (x"cf",x"c1",x"50",x"c1"),
   273 => (x"78",x"c0",x"48",x"fc"),
   274 => (x"97",x"c0",x"d0",x"c1"),
   275 => (x"c1",x"c1",x"49",x"bf"),
   276 => (x"c5",x"c0",x"02",x"a9"),
   277 => (x"c0",x"7e",x"c0",x"87"),
   278 => (x"7e",x"c1",x"87",x"c2"),
   279 => (x"bf",x"fc",x"cf",x"c1"),
   280 => (x"c1",x"b0",x"6e",x"48"),
   281 => (x"c1",x"58",x"c0",x"d0"),
   282 => (x"c1",x"48",x"c4",x"d0"),
   283 => (x"a6",x"dc",x"50",x"c2"),
   284 => (x"c4",x"78",x"c2",x"48"),
   285 => (x"c3",x"78",x"c3",x"80"),
   286 => (x"c0",x"49",x"f8",x"f1"),
   287 => (x"20",x"48",x"f8",x"e9"),
   288 => (x"20",x"41",x"20",x"41"),
   289 => (x"20",x"41",x"20",x"41"),
   290 => (x"20",x"41",x"20",x"41"),
   291 => (x"10",x"51",x"10",x"41"),
   292 => (x"d4",x"51",x"10",x"51"),
   293 => (x"78",x"c1",x"48",x"a6"),
   294 => (x"1e",x"f8",x"f1",x"c3"),
   295 => (x"1e",x"d8",x"f1",x"c3"),
   296 => (x"87",x"ca",x"fb",x"c0"),
   297 => (x"98",x"70",x"86",x"c8"),
   298 => (x"87",x"c5",x"c0",x"05"),
   299 => (x"c2",x"c0",x"49",x"c1"),
   300 => (x"c1",x"49",x"c0",x"87"),
   301 => (x"dc",x"59",x"c0",x"d0"),
   302 => (x"b7",x"c3",x"48",x"66"),
   303 => (x"ee",x"c0",x"03",x"a8"),
   304 => (x"49",x"66",x"dc",x"87"),
   305 => (x"48",x"71",x"91",x"c5"),
   306 => (x"a6",x"d0",x"88",x"c3"),
   307 => (x"1e",x"66",x"d0",x"58"),
   308 => (x"e4",x"c0",x"1e",x"c3"),
   309 => (x"f7",x"c0",x"1e",x"66"),
   310 => (x"86",x"cc",x"87",x"c1"),
   311 => (x"c1",x"48",x"66",x"dc"),
   312 => (x"a6",x"e0",x"c0",x"80"),
   313 => (x"48",x"66",x"dc",x"58"),
   314 => (x"04",x"a8",x"b7",x"c3"),
   315 => (x"cc",x"87",x"d2",x"ff"),
   316 => (x"e0",x"c0",x"1e",x"66"),
   317 => (x"d3",x"c1",x"1e",x"66"),
   318 => (x"d0",x"c1",x"1e",x"d0"),
   319 => (x"f6",x"c0",x"1e",x"c8"),
   320 => (x"86",x"d0",x"87",x"eb"),
   321 => (x"bf",x"f0",x"cf",x"c1"),
   322 => (x"f0",x"cf",x"c1",x"4c"),
   323 => (x"72",x"4b",x"bf",x"bf"),
   324 => (x"c1",x"49",x"73",x"1e"),
   325 => (x"48",x"bf",x"f0",x"cf"),
   326 => (x"4a",x"a1",x"f0",x"c0"),
   327 => (x"aa",x"71",x"41",x"20"),
   328 => (x"87",x"f8",x"ff",x"05"),
   329 => (x"a4",x"c8",x"4a",x"26"),
   330 => (x"49",x"a4",x"cc",x"7e"),
   331 => (x"a3",x"cc",x"79",x"c5"),
   332 => (x"6c",x"7d",x"69",x"4d"),
   333 => (x"d2",x"1e",x"73",x"7b"),
   334 => (x"86",x"c4",x"87",x"c9"),
   335 => (x"69",x"49",x"a3",x"c4"),
   336 => (x"87",x"e6",x"c0",x"05"),
   337 => (x"c6",x"49",x"a3",x"c8"),
   338 => (x"c4",x"1e",x"71",x"7d"),
   339 => (x"c0",x"1e",x"bf",x"66"),
   340 => (x"c8",x"87",x"ec",x"f3"),
   341 => (x"f0",x"cf",x"c1",x"86"),
   342 => (x"75",x"7b",x"bf",x"bf"),
   343 => (x"6d",x"1e",x"ca",x"1e"),
   344 => (x"f6",x"f4",x"c0",x"1e"),
   345 => (x"c0",x"86",x"cc",x"87"),
   346 => (x"49",x"6c",x"87",x"d9"),
   347 => (x"1e",x"72",x"1e",x"71"),
   348 => (x"c0",x"48",x"49",x"74"),
   349 => (x"20",x"4a",x"a1",x"f0"),
   350 => (x"05",x"aa",x"71",x"41"),
   351 => (x"26",x"87",x"f8",x"ff"),
   352 => (x"c1",x"49",x"26",x"4a"),
   353 => (x"c1",x"7e",x"97",x"c1"),
   354 => (x"bf",x"97",x"c4",x"d0"),
   355 => (x"b7",x"c1",x"c1",x"49"),
   356 => (x"e1",x"c1",x"04",x"a9"),
   357 => (x"4b",x"6e",x"97",x"87"),
   358 => (x"73",x"1e",x"c3",x"c1"),
   359 => (x"c0",x"1e",x"71",x"49"),
   360 => (x"c8",x"87",x"e9",x"f6"),
   361 => (x"a8",x"66",x"d4",x"86"),
   362 => (x"87",x"f9",x"c0",x"05"),
   363 => (x"c0",x"1e",x"66",x"d8"),
   364 => (x"ca",x"f2",x"c0",x"1e"),
   365 => (x"71",x"86",x"c8",x"87"),
   366 => (x"f8",x"f1",x"c3",x"1e"),
   367 => (x"d8",x"e9",x"c0",x"49"),
   368 => (x"20",x"41",x"20",x"48"),
   369 => (x"20",x"41",x"20",x"41"),
   370 => (x"20",x"41",x"20",x"41"),
   371 => (x"10",x"41",x"20",x"41"),
   372 => (x"10",x"51",x"10",x"51"),
   373 => (x"c0",x"49",x"26",x"51"),
   374 => (x"c8",x"48",x"a6",x"e0"),
   375 => (x"cf",x"c1",x"78",x"66"),
   376 => (x"66",x"c8",x"48",x"f8"),
   377 => (x"73",x"83",x"c1",x"78"),
   378 => (x"c4",x"d0",x"c1",x"4a"),
   379 => (x"71",x"49",x"bf",x"97"),
   380 => (x"fe",x"06",x"aa",x"b7"),
   381 => (x"e0",x"c0",x"87",x"e2"),
   382 => (x"66",x"dc",x"48",x"66"),
   383 => (x"a6",x"e4",x"c0",x"90"),
   384 => (x"72",x"1e",x"71",x"58"),
   385 => (x"66",x"e8",x"c0",x"1e"),
   386 => (x"4a",x"66",x"d4",x"49"),
   387 => (x"26",x"87",x"f4",x"f3"),
   388 => (x"c0",x"49",x"26",x"4a"),
   389 => (x"c0",x"58",x"a6",x"e0"),
   390 => (x"cc",x"49",x"66",x"e0"),
   391 => (x"91",x"c7",x"89",x"66"),
   392 => (x"66",x"dc",x"48",x"71"),
   393 => (x"a6",x"e4",x"c0",x"88"),
   394 => (x"bf",x"66",x"c4",x"58"),
   395 => (x"c1",x"82",x"ca",x"4a"),
   396 => (x"bf",x"97",x"c0",x"d0"),
   397 => (x"a9",x"c1",x"c1",x"49"),
   398 => (x"87",x"ce",x"c0",x"05"),
   399 => (x"48",x"72",x"8a",x"c1"),
   400 => (x"bf",x"f8",x"cf",x"c1"),
   401 => (x"08",x"66",x"c4",x"88"),
   402 => (x"66",x"c8",x"08",x"78"),
   403 => (x"cc",x"80",x"c1",x"48"),
   404 => (x"66",x"c8",x"58",x"a6"),
   405 => (x"f0",x"e7",x"c0",x"48"),
   406 => (x"06",x"a8",x"b7",x"bf"),
   407 => (x"c3",x"87",x"dc",x"f7"),
   408 => (x"ff",x"48",x"e4",x"ef"),
   409 => (x"c0",x"78",x"bf",x"c8"),
   410 => (x"f0",x"1e",x"f0",x"f0"),
   411 => (x"86",x"c4",x"87",x"f4"),
   412 => (x"1e",x"c0",x"f1",x"c0"),
   413 => (x"c4",x"87",x"eb",x"f0"),
   414 => (x"c4",x"f1",x"c0",x"86"),
   415 => (x"87",x"e2",x"f0",x"1e"),
   416 => (x"f1",x"c0",x"86",x"c4"),
   417 => (x"d9",x"f0",x"1e",x"fc"),
   418 => (x"c1",x"86",x"c4",x"87"),
   419 => (x"1e",x"bf",x"f8",x"cf"),
   420 => (x"1e",x"c0",x"f2",x"c0"),
   421 => (x"c8",x"87",x"cb",x"f0"),
   422 => (x"c0",x"1e",x"c5",x"86"),
   423 => (x"f0",x"1e",x"dc",x"f2"),
   424 => (x"86",x"c8",x"87",x"c0"),
   425 => (x"bf",x"fc",x"cf",x"c1"),
   426 => (x"f8",x"f2",x"c0",x"1e"),
   427 => (x"87",x"f2",x"ef",x"1e"),
   428 => (x"1e",x"c1",x"86",x"c8"),
   429 => (x"1e",x"d4",x"f3",x"c0"),
   430 => (x"c8",x"87",x"e7",x"ef"),
   431 => (x"c0",x"d0",x"c1",x"86"),
   432 => (x"71",x"49",x"bf",x"97"),
   433 => (x"f0",x"f3",x"c0",x"1e"),
   434 => (x"87",x"d6",x"ef",x"1e"),
   435 => (x"c1",x"c1",x"86",x"c8"),
   436 => (x"cc",x"f4",x"c0",x"1e"),
   437 => (x"87",x"ca",x"ef",x"1e"),
   438 => (x"d0",x"c1",x"86",x"c8"),
   439 => (x"49",x"bf",x"97",x"c4"),
   440 => (x"f4",x"c0",x"1e",x"71"),
   441 => (x"f9",x"ee",x"1e",x"e8"),
   442 => (x"c1",x"86",x"c8",x"87"),
   443 => (x"f5",x"c0",x"1e",x"c2"),
   444 => (x"ed",x"ee",x"1e",x"c4"),
   445 => (x"c1",x"86",x"c8",x"87"),
   446 => (x"1e",x"bf",x"e8",x"d0"),
   447 => (x"1e",x"e0",x"f5",x"c0"),
   448 => (x"c8",x"87",x"df",x"ee"),
   449 => (x"c0",x"1e",x"c7",x"86"),
   450 => (x"ee",x"1e",x"fc",x"f5"),
   451 => (x"86",x"c8",x"87",x"d4"),
   452 => (x"bf",x"ec",x"ec",x"c1"),
   453 => (x"d8",x"f6",x"c0",x"1e"),
   454 => (x"87",x"c6",x"ee",x"1e"),
   455 => (x"f6",x"c0",x"86",x"c8"),
   456 => (x"fd",x"ed",x"1e",x"f4"),
   457 => (x"c0",x"86",x"c4",x"87"),
   458 => (x"ed",x"1e",x"e0",x"f7"),
   459 => (x"86",x"c4",x"87",x"f4"),
   460 => (x"bf",x"f0",x"cf",x"c1"),
   461 => (x"f7",x"c0",x"1e",x"bf"),
   462 => (x"e5",x"ed",x"1e",x"ec"),
   463 => (x"c0",x"86",x"c8",x"87"),
   464 => (x"ed",x"1e",x"c8",x"f8"),
   465 => (x"86",x"c4",x"87",x"dc"),
   466 => (x"bf",x"f0",x"cf",x"c1"),
   467 => (x"69",x"81",x"c4",x"49"),
   468 => (x"fc",x"f8",x"c0",x"1e"),
   469 => (x"87",x"ca",x"ed",x"1e"),
   470 => (x"1e",x"c0",x"86",x"c8"),
   471 => (x"1e",x"d8",x"f9",x"c0"),
   472 => (x"c8",x"87",x"ff",x"ec"),
   473 => (x"f0",x"cf",x"c1",x"86"),
   474 => (x"81",x"c8",x"49",x"bf"),
   475 => (x"f9",x"c0",x"1e",x"69"),
   476 => (x"ed",x"ec",x"1e",x"f4"),
   477 => (x"c2",x"86",x"c8",x"87"),
   478 => (x"d0",x"fa",x"c0",x"1e"),
   479 => (x"87",x"e2",x"ec",x"1e"),
   480 => (x"cf",x"c1",x"86",x"c8"),
   481 => (x"cc",x"49",x"bf",x"f0"),
   482 => (x"c0",x"1e",x"69",x"81"),
   483 => (x"ec",x"1e",x"ec",x"fa"),
   484 => (x"86",x"c8",x"87",x"d0"),
   485 => (x"fb",x"c0",x"1e",x"d1"),
   486 => (x"c5",x"ec",x"1e",x"c8"),
   487 => (x"c1",x"86",x"c8",x"87"),
   488 => (x"49",x"bf",x"f0",x"cf"),
   489 => (x"1e",x"71",x"81",x"d0"),
   490 => (x"1e",x"e4",x"fb",x"c0"),
   491 => (x"c8",x"87",x"f3",x"eb"),
   492 => (x"c0",x"fc",x"c0",x"86"),
   493 => (x"87",x"ea",x"eb",x"1e"),
   494 => (x"fc",x"c0",x"86",x"c4"),
   495 => (x"e1",x"eb",x"1e",x"f8"),
   496 => (x"c1",x"86",x"c4",x"87"),
   497 => (x"bf",x"bf",x"f4",x"cf"),
   498 => (x"cc",x"fd",x"c0",x"1e"),
   499 => (x"87",x"d2",x"eb",x"1e"),
   500 => (x"fd",x"c0",x"86",x"c8"),
   501 => (x"c9",x"eb",x"1e",x"e8"),
   502 => (x"c1",x"86",x"c4",x"87"),
   503 => (x"49",x"bf",x"f4",x"cf"),
   504 => (x"1e",x"69",x"81",x"c4"),
   505 => (x"1e",x"e8",x"fe",x"c0"),
   506 => (x"c8",x"87",x"f7",x"ea"),
   507 => (x"c0",x"1e",x"c0",x"86"),
   508 => (x"ea",x"1e",x"c4",x"ff"),
   509 => (x"86",x"c8",x"87",x"ec"),
   510 => (x"bf",x"f4",x"cf",x"c1"),
   511 => (x"69",x"81",x"c8",x"49"),
   512 => (x"e0",x"ff",x"c0",x"1e"),
   513 => (x"87",x"da",x"ea",x"1e"),
   514 => (x"1e",x"c1",x"86",x"c8"),
   515 => (x"1e",x"fc",x"ff",x"c0"),
   516 => (x"c8",x"87",x"cf",x"ea"),
   517 => (x"f4",x"cf",x"c1",x"86"),
   518 => (x"81",x"cc",x"49",x"bf"),
   519 => (x"c0",x"c1",x"1e",x"69"),
   520 => (x"fd",x"e9",x"1e",x"d8"),
   521 => (x"d2",x"86",x"c8",x"87"),
   522 => (x"f4",x"c0",x"c1",x"1e"),
   523 => (x"87",x"f2",x"e9",x"1e"),
   524 => (x"cf",x"c1",x"86",x"c8"),
   525 => (x"d0",x"49",x"bf",x"f4"),
   526 => (x"c1",x"1e",x"71",x"81"),
   527 => (x"e9",x"1e",x"d0",x"c1"),
   528 => (x"86",x"c8",x"87",x"e0"),
   529 => (x"1e",x"ec",x"c1",x"c1"),
   530 => (x"c4",x"87",x"d7",x"e9"),
   531 => (x"1e",x"66",x"dc",x"86"),
   532 => (x"1e",x"e4",x"c2",x"c1"),
   533 => (x"c8",x"87",x"cb",x"e9"),
   534 => (x"c1",x"1e",x"c5",x"86"),
   535 => (x"e9",x"1e",x"c0",x"c3"),
   536 => (x"86",x"c8",x"87",x"c0"),
   537 => (x"1e",x"66",x"e0",x"c0"),
   538 => (x"1e",x"dc",x"c3",x"c1"),
   539 => (x"c8",x"87",x"f3",x"e8"),
   540 => (x"c1",x"1e",x"cd",x"86"),
   541 => (x"e8",x"1e",x"f8",x"c3"),
   542 => (x"86",x"c8",x"87",x"e8"),
   543 => (x"c1",x"1e",x"66",x"cc"),
   544 => (x"e8",x"1e",x"d4",x"c4"),
   545 => (x"86",x"c8",x"87",x"dc"),
   546 => (x"c4",x"c1",x"1e",x"c7"),
   547 => (x"d1",x"e8",x"1e",x"f0"),
   548 => (x"d4",x"86",x"c8",x"87"),
   549 => (x"c5",x"c1",x"1e",x"66"),
   550 => (x"c5",x"e8",x"1e",x"cc"),
   551 => (x"c1",x"86",x"c8",x"87"),
   552 => (x"e8",x"c5",x"c1",x"1e"),
   553 => (x"87",x"fa",x"e7",x"1e"),
   554 => (x"f1",x"c3",x"86",x"c8"),
   555 => (x"c6",x"c1",x"1e",x"d8"),
   556 => (x"ed",x"e7",x"1e",x"c4"),
   557 => (x"c1",x"86",x"c8",x"87"),
   558 => (x"e7",x"1e",x"e0",x"c6"),
   559 => (x"86",x"c4",x"87",x"e4"),
   560 => (x"1e",x"f8",x"f1",x"c3"),
   561 => (x"1e",x"d8",x"c7",x"c1"),
   562 => (x"c8",x"87",x"d7",x"e7"),
   563 => (x"f4",x"c7",x"c1",x"86"),
   564 => (x"87",x"ce",x"e7",x"1e"),
   565 => (x"c8",x"c1",x"86",x"c4"),
   566 => (x"c5",x"e7",x"1e",x"ec"),
   567 => (x"c3",x"86",x"c4",x"87"),
   568 => (x"49",x"bf",x"e4",x"ef"),
   569 => (x"bf",x"e0",x"ef",x"c3"),
   570 => (x"ec",x"ef",x"c3",x"89"),
   571 => (x"c1",x"1e",x"71",x"59"),
   572 => (x"e6",x"1e",x"f0",x"c8"),
   573 => (x"86",x"c8",x"87",x"ec"),
   574 => (x"bf",x"e8",x"ef",x"c3"),
   575 => (x"b7",x"f8",x"c1",x"48"),
   576 => (x"db",x"c0",x"03",x"a8"),
   577 => (x"d8",x"ea",x"c0",x"87"),
   578 => (x"87",x"d6",x"e6",x"1e"),
   579 => (x"eb",x"c0",x"86",x"c4"),
   580 => (x"cd",x"e6",x"1e",x"d0"),
   581 => (x"c0",x"86",x"c4",x"87"),
   582 => (x"e6",x"1e",x"f0",x"eb"),
   583 => (x"86",x"c4",x"87",x"c4"),
   584 => (x"bf",x"e8",x"ef",x"c3"),
   585 => (x"cf",x"4a",x"71",x"49"),
   586 => (x"1e",x"71",x"92",x"e8"),
   587 => (x"49",x"72",x"1e",x"72"),
   588 => (x"bf",x"f0",x"e7",x"c0"),
   589 => (x"87",x"cb",x"e7",x"4a"),
   590 => (x"49",x"26",x"4a",x"26"),
   591 => (x"58",x"f0",x"ef",x"c3"),
   592 => (x"bf",x"f0",x"e7",x"c0"),
   593 => (x"cf",x"4b",x"72",x"4a"),
   594 => (x"1e",x"71",x"93",x"e8"),
   595 => (x"09",x"73",x"1e",x"72"),
   596 => (x"87",x"ef",x"e6",x"4a"),
   597 => (x"49",x"26",x"4a",x"26"),
   598 => (x"58",x"f4",x"ef",x"c3"),
   599 => (x"71",x"92",x"f9",x"c8"),
   600 => (x"72",x"1e",x"72",x"1e"),
   601 => (x"da",x"e6",x"4a",x"09"),
   602 => (x"26",x"4a",x"26",x"87"),
   603 => (x"f8",x"ef",x"c3",x"49"),
   604 => (x"f4",x"eb",x"c0",x"58"),
   605 => (x"87",x"ea",x"e4",x"1e"),
   606 => (x"ef",x"c3",x"86",x"c4"),
   607 => (x"c0",x"1e",x"bf",x"ec"),
   608 => (x"e4",x"1e",x"e4",x"ec"),
   609 => (x"86",x"c8",x"87",x"dc"),
   610 => (x"1e",x"ec",x"ec",x"c0"),
   611 => (x"c4",x"87",x"d3",x"e4"),
   612 => (x"f0",x"ef",x"c3",x"86"),
   613 => (x"ed",x"c0",x"1e",x"bf"),
   614 => (x"c5",x"e4",x"1e",x"dc"),
   615 => (x"c3",x"86",x"c8",x"87"),
   616 => (x"1e",x"bf",x"f4",x"ef"),
   617 => (x"1e",x"e4",x"ed",x"c0"),
   618 => (x"c8",x"87",x"f7",x"e3"),
   619 => (x"c4",x"ee",x"c0",x"86"),
   620 => (x"87",x"ee",x"e3",x"1e"),
   621 => (x"48",x"c0",x"86",x"c4"),
   622 => (x"26",x"8e",x"dc",x"ff"),
   623 => (x"26",x"4c",x"26",x"4d"),
   624 => (x"1e",x"4f",x"26",x"4b"),
   625 => (x"bf",x"f0",x"cf",x"c1"),
   626 => (x"c4",x"87",x"c9",x"02"),
   627 => (x"cf",x"c1",x"48",x"66"),
   628 => (x"78",x"bf",x"bf",x"f0"),
   629 => (x"bf",x"f0",x"cf",x"c1"),
   630 => (x"71",x"81",x"cc",x"49"),
   631 => (x"f8",x"cf",x"c1",x"1e"),
   632 => (x"1e",x"ca",x"1e",x"bf"),
   633 => (x"87",x"f3",x"e2",x"c0"),
   634 => (x"4f",x"26",x"86",x"cc"),
   635 => (x"00",x"00",x"00",x"00"),
   636 => (x"00",x"00",x"61",x"a8"),
   637 => (x"67",x"6f",x"72",x"50"),
   638 => (x"20",x"6d",x"61",x"72"),
   639 => (x"70",x"6d",x"6f",x"63"),
   640 => (x"64",x"65",x"6c",x"69"),
   641 => (x"74",x"69",x"77",x"20"),
   642 => (x"72",x"27",x"20",x"68"),
   643 => (x"73",x"69",x"67",x"65"),
   644 => (x"27",x"72",x"65",x"74"),
   645 => (x"74",x"74",x"61",x"20"),
   646 => (x"75",x"62",x"69",x"72"),
   647 => (x"00",x"0a",x"65",x"74"),
   648 => (x"00",x"00",x"00",x"0a"),
   649 => (x"67",x"6f",x"72",x"50"),
   650 => (x"20",x"6d",x"61",x"72"),
   651 => (x"70",x"6d",x"6f",x"63"),
   652 => (x"64",x"65",x"6c",x"69"),
   653 => (x"74",x"69",x"77",x"20"),
   654 => (x"74",x"75",x"6f",x"68"),
   655 => (x"65",x"72",x"27",x"20"),
   656 => (x"74",x"73",x"69",x"67"),
   657 => (x"20",x"27",x"72",x"65"),
   658 => (x"72",x"74",x"74",x"61"),
   659 => (x"74",x"75",x"62",x"69"),
   660 => (x"00",x"00",x"0a",x"65"),
   661 => (x"00",x"00",x"00",x"0a"),
   662 => (x"59",x"52",x"48",x"44"),
   663 => (x"4e",x"4f",x"54",x"53"),
   664 => (x"52",x"50",x"20",x"45"),
   665 => (x"41",x"52",x"47",x"4f"),
   666 => (x"33",x"20",x"2c",x"4d"),
   667 => (x"20",x"44",x"52",x"27"),
   668 => (x"49",x"52",x"54",x"53"),
   669 => (x"00",x"00",x"47",x"4e"),
   670 => (x"59",x"52",x"48",x"44"),
   671 => (x"4e",x"4f",x"54",x"53"),
   672 => (x"52",x"50",x"20",x"45"),
   673 => (x"41",x"52",x"47",x"4f"),
   674 => (x"32",x"20",x"2c",x"4d"),
   675 => (x"20",x"44",x"4e",x"27"),
   676 => (x"49",x"52",x"54",x"53"),
   677 => (x"00",x"00",x"47",x"4e"),
   678 => (x"73",x"61",x"65",x"4d"),
   679 => (x"64",x"65",x"72",x"75"),
   680 => (x"6d",x"69",x"74",x"20"),
   681 => (x"6f",x"74",x"20",x"65"),
   682 => (x"6d",x"73",x"20",x"6f"),
   683 => (x"20",x"6c",x"6c",x"61"),
   684 => (x"6f",x"20",x"6f",x"74"),
   685 => (x"69",x"61",x"74",x"62"),
   686 => (x"65",x"6d",x"20",x"6e"),
   687 => (x"6e",x"69",x"6e",x"61"),
   688 => (x"6c",x"75",x"66",x"67"),
   689 => (x"73",x"65",x"72",x"20"),
   690 => (x"73",x"74",x"6c",x"75"),
   691 => (x"00",x"00",x"00",x"0a"),
   692 => (x"61",x"65",x"6c",x"50"),
   693 => (x"69",x"20",x"65",x"73"),
   694 => (x"65",x"72",x"63",x"6e"),
   695 => (x"20",x"65",x"73",x"61"),
   696 => (x"62",x"6d",x"75",x"6e"),
   697 => (x"6f",x"20",x"72",x"65"),
   698 => (x"75",x"72",x"20",x"66"),
   699 => (x"00",x"0a",x"73",x"6e"),
   700 => (x"00",x"00",x"00",x"0a"),
   701 => (x"72",x"63",x"69",x"4d"),
   702 => (x"63",x"65",x"73",x"6f"),
   703 => (x"73",x"64",x"6e",x"6f"),
   704 => (x"72",x"6f",x"66",x"20"),
   705 => (x"65",x"6e",x"6f",x"20"),
   706 => (x"6e",x"75",x"72",x"20"),
   707 => (x"72",x"68",x"74",x"20"),
   708 => (x"68",x"67",x"75",x"6f"),
   709 => (x"72",x"68",x"44",x"20"),
   710 => (x"6f",x"74",x"73",x"79"),
   711 => (x"20",x"3a",x"65",x"6e"),
   712 => (x"00",x"00",x"00",x"00"),
   713 => (x"0a",x"20",x"64",x"25"),
   714 => (x"00",x"00",x"00",x"00"),
   715 => (x"79",x"72",x"68",x"44"),
   716 => (x"6e",x"6f",x"74",x"73"),
   717 => (x"70",x"20",x"73",x"65"),
   718 => (x"53",x"20",x"72",x"65"),
   719 => (x"6e",x"6f",x"63",x"65"),
   720 => (x"20",x"20",x"3a",x"64"),
   721 => (x"20",x"20",x"20",x"20"),
   722 => (x"20",x"20",x"20",x"20"),
   723 => (x"20",x"20",x"20",x"20"),
   724 => (x"20",x"20",x"20",x"20"),
   725 => (x"20",x"20",x"20",x"20"),
   726 => (x"00",x"00",x"00",x"00"),
   727 => (x"0a",x"20",x"64",x"25"),
   728 => (x"00",x"00",x"00",x"00"),
   729 => (x"20",x"58",x"41",x"56"),
   730 => (x"53",x"50",x"49",x"4d"),
   731 => (x"74",x"61",x"72",x"20"),
   732 => (x"20",x"67",x"6e",x"69"),
   733 => (x"30",x"31",x"20",x"2a"),
   734 => (x"3d",x"20",x"30",x"30"),
   735 => (x"20",x"64",x"25",x"20"),
   736 => (x"00",x"00",x"00",x"0a"),
   737 => (x"00",x"00",x"00",x"0a"),
   738 => (x"59",x"52",x"48",x"44"),
   739 => (x"4e",x"4f",x"54",x"53"),
   740 => (x"52",x"50",x"20",x"45"),
   741 => (x"41",x"52",x"47",x"4f"),
   742 => (x"53",x"20",x"2c",x"4d"),
   743 => (x"20",x"45",x"4d",x"4f"),
   744 => (x"49",x"52",x"54",x"53"),
   745 => (x"00",x"00",x"47",x"4e"),
   746 => (x"59",x"52",x"48",x"44"),
   747 => (x"4e",x"4f",x"54",x"53"),
   748 => (x"52",x"50",x"20",x"45"),
   749 => (x"41",x"52",x"47",x"4f"),
   750 => (x"31",x"20",x"2c",x"4d"),
   751 => (x"20",x"54",x"53",x"27"),
   752 => (x"49",x"52",x"54",x"53"),
   753 => (x"00",x"00",x"47",x"4e"),
   754 => (x"00",x"00",x"00",x"0a"),
   755 => (x"79",x"72",x"68",x"44"),
   756 => (x"6e",x"6f",x"74",x"73"),
   757 => (x"65",x"42",x"20",x"65"),
   758 => (x"6d",x"68",x"63",x"6e"),
   759 => (x"2c",x"6b",x"72",x"61"),
   760 => (x"72",x"65",x"56",x"20"),
   761 => (x"6e",x"6f",x"69",x"73"),
   762 => (x"31",x"2e",x"32",x"20"),
   763 => (x"61",x"4c",x"28",x"20"),
   764 => (x"61",x"75",x"67",x"6e"),
   765 => (x"20",x"3a",x"65",x"67"),
   766 => (x"00",x"0a",x"29",x"43"),
   767 => (x"00",x"00",x"00",x"0a"),
   768 => (x"63",x"65",x"78",x"45"),
   769 => (x"6f",x"69",x"74",x"75"),
   770 => (x"74",x"73",x"20",x"6e"),
   771 => (x"73",x"74",x"72",x"61"),
   772 => (x"64",x"25",x"20",x"2c"),
   773 => (x"6e",x"75",x"72",x"20"),
   774 => (x"68",x"74",x"20",x"73"),
   775 => (x"67",x"75",x"6f",x"72"),
   776 => (x"68",x"44",x"20",x"68"),
   777 => (x"74",x"73",x"79",x"72"),
   778 => (x"0a",x"65",x"6e",x"6f"),
   779 => (x"00",x"00",x"00",x"00"),
   780 => (x"63",x"65",x"78",x"45"),
   781 => (x"6f",x"69",x"74",x"75"),
   782 => (x"6e",x"65",x"20",x"6e"),
   783 => (x"00",x"0a",x"73",x"64"),
   784 => (x"00",x"00",x"00",x"0a"),
   785 => (x"61",x"6e",x"69",x"46"),
   786 => (x"61",x"76",x"20",x"6c"),
   787 => (x"73",x"65",x"75",x"6c"),
   788 => (x"20",x"66",x"6f",x"20"),
   789 => (x"20",x"65",x"68",x"74"),
   790 => (x"69",x"72",x"61",x"76"),
   791 => (x"65",x"6c",x"62",x"61"),
   792 => (x"73",x"75",x"20",x"73"),
   793 => (x"69",x"20",x"64",x"65"),
   794 => (x"68",x"74",x"20",x"6e"),
   795 => (x"65",x"62",x"20",x"65"),
   796 => (x"6d",x"68",x"63",x"6e"),
   797 => (x"3a",x"6b",x"72",x"61"),
   798 => (x"00",x"00",x"00",x"0a"),
   799 => (x"00",x"00",x"00",x"0a"),
   800 => (x"5f",x"74",x"6e",x"49"),
   801 => (x"62",x"6f",x"6c",x"47"),
   802 => (x"20",x"20",x"20",x"3a"),
   803 => (x"20",x"20",x"20",x"20"),
   804 => (x"20",x"20",x"20",x"20"),
   805 => (x"0a",x"64",x"25",x"20"),
   806 => (x"00",x"00",x"00",x"00"),
   807 => (x"20",x"20",x"20",x"20"),
   808 => (x"20",x"20",x"20",x"20"),
   809 => (x"75",x"6f",x"68",x"73"),
   810 => (x"62",x"20",x"64",x"6c"),
   811 => (x"20",x"20",x"3a",x"65"),
   812 => (x"0a",x"64",x"25",x"20"),
   813 => (x"00",x"00",x"00",x"00"),
   814 => (x"6c",x"6f",x"6f",x"42"),
   815 => (x"6f",x"6c",x"47",x"5f"),
   816 => (x"20",x"20",x"3a",x"62"),
   817 => (x"20",x"20",x"20",x"20"),
   818 => (x"20",x"20",x"20",x"20"),
   819 => (x"0a",x"64",x"25",x"20"),
   820 => (x"00",x"00",x"00",x"00"),
   821 => (x"20",x"20",x"20",x"20"),
   822 => (x"20",x"20",x"20",x"20"),
   823 => (x"75",x"6f",x"68",x"73"),
   824 => (x"62",x"20",x"64",x"6c"),
   825 => (x"20",x"20",x"3a",x"65"),
   826 => (x"0a",x"64",x"25",x"20"),
   827 => (x"00",x"00",x"00",x"00"),
   828 => (x"31",x"5f",x"68",x"43"),
   829 => (x"6f",x"6c",x"47",x"5f"),
   830 => (x"20",x"20",x"3a",x"62"),
   831 => (x"20",x"20",x"20",x"20"),
   832 => (x"20",x"20",x"20",x"20"),
   833 => (x"0a",x"63",x"25",x"20"),
   834 => (x"00",x"00",x"00",x"00"),
   835 => (x"20",x"20",x"20",x"20"),
   836 => (x"20",x"20",x"20",x"20"),
   837 => (x"75",x"6f",x"68",x"73"),
   838 => (x"62",x"20",x"64",x"6c"),
   839 => (x"20",x"20",x"3a",x"65"),
   840 => (x"0a",x"63",x"25",x"20"),
   841 => (x"00",x"00",x"00",x"00"),
   842 => (x"32",x"5f",x"68",x"43"),
   843 => (x"6f",x"6c",x"47",x"5f"),
   844 => (x"20",x"20",x"3a",x"62"),
   845 => (x"20",x"20",x"20",x"20"),
   846 => (x"20",x"20",x"20",x"20"),
   847 => (x"0a",x"63",x"25",x"20"),
   848 => (x"00",x"00",x"00",x"00"),
   849 => (x"20",x"20",x"20",x"20"),
   850 => (x"20",x"20",x"20",x"20"),
   851 => (x"75",x"6f",x"68",x"73"),
   852 => (x"62",x"20",x"64",x"6c"),
   853 => (x"20",x"20",x"3a",x"65"),
   854 => (x"0a",x"63",x"25",x"20"),
   855 => (x"00",x"00",x"00",x"00"),
   856 => (x"5f",x"72",x"72",x"41"),
   857 => (x"6c",x"47",x"5f",x"31"),
   858 => (x"38",x"5b",x"62",x"6f"),
   859 => (x"20",x"20",x"3a",x"5d"),
   860 => (x"20",x"20",x"20",x"20"),
   861 => (x"0a",x"64",x"25",x"20"),
   862 => (x"00",x"00",x"00",x"00"),
   863 => (x"20",x"20",x"20",x"20"),
   864 => (x"20",x"20",x"20",x"20"),
   865 => (x"75",x"6f",x"68",x"73"),
   866 => (x"62",x"20",x"64",x"6c"),
   867 => (x"20",x"20",x"3a",x"65"),
   868 => (x"0a",x"64",x"25",x"20"),
   869 => (x"00",x"00",x"00",x"00"),
   870 => (x"5f",x"72",x"72",x"41"),
   871 => (x"6c",x"47",x"5f",x"32"),
   872 => (x"38",x"5b",x"62",x"6f"),
   873 => (x"5d",x"37",x"5b",x"5d"),
   874 => (x"20",x"20",x"20",x"3a"),
   875 => (x"0a",x"64",x"25",x"20"),
   876 => (x"00",x"00",x"00",x"00"),
   877 => (x"20",x"20",x"20",x"20"),
   878 => (x"20",x"20",x"20",x"20"),
   879 => (x"75",x"6f",x"68",x"73"),
   880 => (x"62",x"20",x"64",x"6c"),
   881 => (x"20",x"20",x"3a",x"65"),
   882 => (x"6d",x"75",x"4e",x"20"),
   883 => (x"5f",x"72",x"65",x"62"),
   884 => (x"52",x"5f",x"66",x"4f"),
   885 => (x"20",x"73",x"6e",x"75"),
   886 => (x"30",x"31",x"20",x"2b"),
   887 => (x"00",x"00",x"00",x"0a"),
   888 => (x"5f",x"72",x"74",x"50"),
   889 => (x"62",x"6f",x"6c",x"47"),
   890 => (x"00",x"0a",x"3e",x"2d"),
   891 => (x"74",x"50",x"20",x"20"),
   892 => (x"6f",x"43",x"5f",x"72"),
   893 => (x"20",x"3a",x"70",x"6d"),
   894 => (x"20",x"20",x"20",x"20"),
   895 => (x"20",x"20",x"20",x"20"),
   896 => (x"0a",x"64",x"25",x"20"),
   897 => (x"00",x"00",x"00",x"00"),
   898 => (x"20",x"20",x"20",x"20"),
   899 => (x"20",x"20",x"20",x"20"),
   900 => (x"75",x"6f",x"68",x"73"),
   901 => (x"62",x"20",x"64",x"6c"),
   902 => (x"20",x"20",x"3a",x"65"),
   903 => (x"6d",x"69",x"28",x"20"),
   904 => (x"6d",x"65",x"6c",x"70"),
   905 => (x"61",x"74",x"6e",x"65"),
   906 => (x"6e",x"6f",x"69",x"74"),
   907 => (x"70",x"65",x"64",x"2d"),
   908 => (x"65",x"64",x"6e",x"65"),
   909 => (x"0a",x"29",x"74",x"6e"),
   910 => (x"00",x"00",x"00",x"00"),
   911 => (x"69",x"44",x"20",x"20"),
   912 => (x"3a",x"72",x"63",x"73"),
   913 => (x"20",x"20",x"20",x"20"),
   914 => (x"20",x"20",x"20",x"20"),
   915 => (x"20",x"20",x"20",x"20"),
   916 => (x"0a",x"64",x"25",x"20"),
   917 => (x"00",x"00",x"00",x"00"),
   918 => (x"20",x"20",x"20",x"20"),
   919 => (x"20",x"20",x"20",x"20"),
   920 => (x"75",x"6f",x"68",x"73"),
   921 => (x"62",x"20",x"64",x"6c"),
   922 => (x"20",x"20",x"3a",x"65"),
   923 => (x"0a",x"64",x"25",x"20"),
   924 => (x"00",x"00",x"00",x"00"),
   925 => (x"6e",x"45",x"20",x"20"),
   926 => (x"43",x"5f",x"6d",x"75"),
   927 => (x"3a",x"70",x"6d",x"6f"),
   928 => (x"20",x"20",x"20",x"20"),
   929 => (x"20",x"20",x"20",x"20"),
   930 => (x"0a",x"64",x"25",x"20"),
   931 => (x"00",x"00",x"00",x"00"),
   932 => (x"20",x"20",x"20",x"20"),
   933 => (x"20",x"20",x"20",x"20"),
   934 => (x"75",x"6f",x"68",x"73"),
   935 => (x"62",x"20",x"64",x"6c"),
   936 => (x"20",x"20",x"3a",x"65"),
   937 => (x"0a",x"64",x"25",x"20"),
   938 => (x"00",x"00",x"00",x"00"),
   939 => (x"6e",x"49",x"20",x"20"),
   940 => (x"6f",x"43",x"5f",x"74"),
   941 => (x"20",x"3a",x"70",x"6d"),
   942 => (x"20",x"20",x"20",x"20"),
   943 => (x"20",x"20",x"20",x"20"),
   944 => (x"0a",x"64",x"25",x"20"),
   945 => (x"00",x"00",x"00",x"00"),
   946 => (x"20",x"20",x"20",x"20"),
   947 => (x"20",x"20",x"20",x"20"),
   948 => (x"75",x"6f",x"68",x"73"),
   949 => (x"62",x"20",x"64",x"6c"),
   950 => (x"20",x"20",x"3a",x"65"),
   951 => (x"0a",x"64",x"25",x"20"),
   952 => (x"00",x"00",x"00",x"00"),
   953 => (x"74",x"53",x"20",x"20"),
   954 => (x"6f",x"43",x"5f",x"72"),
   955 => (x"20",x"3a",x"70",x"6d"),
   956 => (x"20",x"20",x"20",x"20"),
   957 => (x"20",x"20",x"20",x"20"),
   958 => (x"0a",x"73",x"25",x"20"),
   959 => (x"00",x"00",x"00",x"00"),
   960 => (x"20",x"20",x"20",x"20"),
   961 => (x"20",x"20",x"20",x"20"),
   962 => (x"75",x"6f",x"68",x"73"),
   963 => (x"62",x"20",x"64",x"6c"),
   964 => (x"20",x"20",x"3a",x"65"),
   965 => (x"52",x"48",x"44",x"20"),
   966 => (x"4f",x"54",x"53",x"59"),
   967 => (x"50",x"20",x"45",x"4e"),
   968 => (x"52",x"47",x"4f",x"52"),
   969 => (x"20",x"2c",x"4d",x"41"),
   970 => (x"45",x"4d",x"4f",x"53"),
   971 => (x"52",x"54",x"53",x"20"),
   972 => (x"0a",x"47",x"4e",x"49"),
   973 => (x"00",x"00",x"00",x"00"),
   974 => (x"74",x"78",x"65",x"4e"),
   975 => (x"72",x"74",x"50",x"5f"),
   976 => (x"6f",x"6c",x"47",x"5f"),
   977 => (x"0a",x"3e",x"2d",x"62"),
   978 => (x"00",x"00",x"00",x"00"),
   979 => (x"74",x"50",x"20",x"20"),
   980 => (x"6f",x"43",x"5f",x"72"),
   981 => (x"20",x"3a",x"70",x"6d"),
   982 => (x"20",x"20",x"20",x"20"),
   983 => (x"20",x"20",x"20",x"20"),
   984 => (x"0a",x"64",x"25",x"20"),
   985 => (x"00",x"00",x"00",x"00"),
   986 => (x"20",x"20",x"20",x"20"),
   987 => (x"20",x"20",x"20",x"20"),
   988 => (x"75",x"6f",x"68",x"73"),
   989 => (x"62",x"20",x"64",x"6c"),
   990 => (x"20",x"20",x"3a",x"65"),
   991 => (x"6d",x"69",x"28",x"20"),
   992 => (x"6d",x"65",x"6c",x"70"),
   993 => (x"61",x"74",x"6e",x"65"),
   994 => (x"6e",x"6f",x"69",x"74"),
   995 => (x"70",x"65",x"64",x"2d"),
   996 => (x"65",x"64",x"6e",x"65"),
   997 => (x"2c",x"29",x"74",x"6e"),
   998 => (x"6d",x"61",x"73",x"20"),
   999 => (x"73",x"61",x"20",x"65"),
  1000 => (x"6f",x"62",x"61",x"20"),
  1001 => (x"00",x"0a",x"65",x"76"),
  1002 => (x"69",x"44",x"20",x"20"),
  1003 => (x"3a",x"72",x"63",x"73"),
  1004 => (x"20",x"20",x"20",x"20"),
  1005 => (x"20",x"20",x"20",x"20"),
  1006 => (x"20",x"20",x"20",x"20"),
  1007 => (x"0a",x"64",x"25",x"20"),
  1008 => (x"00",x"00",x"00",x"00"),
  1009 => (x"20",x"20",x"20",x"20"),
  1010 => (x"20",x"20",x"20",x"20"),
  1011 => (x"75",x"6f",x"68",x"73"),
  1012 => (x"62",x"20",x"64",x"6c"),
  1013 => (x"20",x"20",x"3a",x"65"),
  1014 => (x"0a",x"64",x"25",x"20"),
  1015 => (x"00",x"00",x"00",x"00"),
  1016 => (x"6e",x"45",x"20",x"20"),
  1017 => (x"43",x"5f",x"6d",x"75"),
  1018 => (x"3a",x"70",x"6d",x"6f"),
  1019 => (x"20",x"20",x"20",x"20"),
  1020 => (x"20",x"20",x"20",x"20"),
  1021 => (x"0a",x"64",x"25",x"20"),
  1022 => (x"00",x"00",x"00",x"00"),
  1023 => (x"20",x"20",x"20",x"20"),
  1024 => (x"20",x"20",x"20",x"20"),
  1025 => (x"75",x"6f",x"68",x"73"),
  1026 => (x"62",x"20",x"64",x"6c"),
  1027 => (x"20",x"20",x"3a",x"65"),
  1028 => (x"0a",x"64",x"25",x"20"),
  1029 => (x"00",x"00",x"00",x"00"),
  1030 => (x"6e",x"49",x"20",x"20"),
  1031 => (x"6f",x"43",x"5f",x"74"),
  1032 => (x"20",x"3a",x"70",x"6d"),
  1033 => (x"20",x"20",x"20",x"20"),
  1034 => (x"20",x"20",x"20",x"20"),
  1035 => (x"0a",x"64",x"25",x"20"),
  1036 => (x"00",x"00",x"00",x"00"),
  1037 => (x"20",x"20",x"20",x"20"),
  1038 => (x"20",x"20",x"20",x"20"),
  1039 => (x"75",x"6f",x"68",x"73"),
  1040 => (x"62",x"20",x"64",x"6c"),
  1041 => (x"20",x"20",x"3a",x"65"),
  1042 => (x"0a",x"64",x"25",x"20"),
  1043 => (x"00",x"00",x"00",x"00"),
  1044 => (x"74",x"53",x"20",x"20"),
  1045 => (x"6f",x"43",x"5f",x"72"),
  1046 => (x"20",x"3a",x"70",x"6d"),
  1047 => (x"20",x"20",x"20",x"20"),
  1048 => (x"20",x"20",x"20",x"20"),
  1049 => (x"0a",x"73",x"25",x"20"),
  1050 => (x"00",x"00",x"00",x"00"),
  1051 => (x"20",x"20",x"20",x"20"),
  1052 => (x"20",x"20",x"20",x"20"),
  1053 => (x"75",x"6f",x"68",x"73"),
  1054 => (x"62",x"20",x"64",x"6c"),
  1055 => (x"20",x"20",x"3a",x"65"),
  1056 => (x"52",x"48",x"44",x"20"),
  1057 => (x"4f",x"54",x"53",x"59"),
  1058 => (x"50",x"20",x"45",x"4e"),
  1059 => (x"52",x"47",x"4f",x"52"),
  1060 => (x"20",x"2c",x"4d",x"41"),
  1061 => (x"45",x"4d",x"4f",x"53"),
  1062 => (x"52",x"54",x"53",x"20"),
  1063 => (x"0a",x"47",x"4e",x"49"),
  1064 => (x"00",x"00",x"00",x"00"),
  1065 => (x"5f",x"74",x"6e",x"49"),
  1066 => (x"6f",x"4c",x"5f",x"31"),
  1067 => (x"20",x"20",x"3a",x"63"),
  1068 => (x"20",x"20",x"20",x"20"),
  1069 => (x"20",x"20",x"20",x"20"),
  1070 => (x"0a",x"64",x"25",x"20"),
  1071 => (x"00",x"00",x"00",x"00"),
  1072 => (x"20",x"20",x"20",x"20"),
  1073 => (x"20",x"20",x"20",x"20"),
  1074 => (x"75",x"6f",x"68",x"73"),
  1075 => (x"62",x"20",x"64",x"6c"),
  1076 => (x"20",x"20",x"3a",x"65"),
  1077 => (x"0a",x"64",x"25",x"20"),
  1078 => (x"00",x"00",x"00",x"00"),
  1079 => (x"5f",x"74",x"6e",x"49"),
  1080 => (x"6f",x"4c",x"5f",x"32"),
  1081 => (x"20",x"20",x"3a",x"63"),
  1082 => (x"20",x"20",x"20",x"20"),
  1083 => (x"20",x"20",x"20",x"20"),
  1084 => (x"0a",x"64",x"25",x"20"),
  1085 => (x"00",x"00",x"00",x"00"),
  1086 => (x"20",x"20",x"20",x"20"),
  1087 => (x"20",x"20",x"20",x"20"),
  1088 => (x"75",x"6f",x"68",x"73"),
  1089 => (x"62",x"20",x"64",x"6c"),
  1090 => (x"20",x"20",x"3a",x"65"),
  1091 => (x"0a",x"64",x"25",x"20"),
  1092 => (x"00",x"00",x"00",x"00"),
  1093 => (x"5f",x"74",x"6e",x"49"),
  1094 => (x"6f",x"4c",x"5f",x"33"),
  1095 => (x"20",x"20",x"3a",x"63"),
  1096 => (x"20",x"20",x"20",x"20"),
  1097 => (x"20",x"20",x"20",x"20"),
  1098 => (x"0a",x"64",x"25",x"20"),
  1099 => (x"00",x"00",x"00",x"00"),
  1100 => (x"20",x"20",x"20",x"20"),
  1101 => (x"20",x"20",x"20",x"20"),
  1102 => (x"75",x"6f",x"68",x"73"),
  1103 => (x"62",x"20",x"64",x"6c"),
  1104 => (x"20",x"20",x"3a",x"65"),
  1105 => (x"0a",x"64",x"25",x"20"),
  1106 => (x"00",x"00",x"00",x"00"),
  1107 => (x"6d",x"75",x"6e",x"45"),
  1108 => (x"63",x"6f",x"4c",x"5f"),
  1109 => (x"20",x"20",x"20",x"3a"),
  1110 => (x"20",x"20",x"20",x"20"),
  1111 => (x"20",x"20",x"20",x"20"),
  1112 => (x"0a",x"64",x"25",x"20"),
  1113 => (x"00",x"00",x"00",x"00"),
  1114 => (x"20",x"20",x"20",x"20"),
  1115 => (x"20",x"20",x"20",x"20"),
  1116 => (x"75",x"6f",x"68",x"73"),
  1117 => (x"62",x"20",x"64",x"6c"),
  1118 => (x"20",x"20",x"3a",x"65"),
  1119 => (x"0a",x"64",x"25",x"20"),
  1120 => (x"00",x"00",x"00",x"00"),
  1121 => (x"5f",x"72",x"74",x"53"),
  1122 => (x"6f",x"4c",x"5f",x"31"),
  1123 => (x"20",x"20",x"3a",x"63"),
  1124 => (x"20",x"20",x"20",x"20"),
  1125 => (x"20",x"20",x"20",x"20"),
  1126 => (x"0a",x"73",x"25",x"20"),
  1127 => (x"00",x"00",x"00",x"00"),
  1128 => (x"20",x"20",x"20",x"20"),
  1129 => (x"20",x"20",x"20",x"20"),
  1130 => (x"75",x"6f",x"68",x"73"),
  1131 => (x"62",x"20",x"64",x"6c"),
  1132 => (x"20",x"20",x"3a",x"65"),
  1133 => (x"52",x"48",x"44",x"20"),
  1134 => (x"4f",x"54",x"53",x"59"),
  1135 => (x"50",x"20",x"45",x"4e"),
  1136 => (x"52",x"47",x"4f",x"52"),
  1137 => (x"20",x"2c",x"4d",x"41"),
  1138 => (x"54",x"53",x"27",x"31"),
  1139 => (x"52",x"54",x"53",x"20"),
  1140 => (x"0a",x"47",x"4e",x"49"),
  1141 => (x"00",x"00",x"00",x"00"),
  1142 => (x"5f",x"72",x"74",x"53"),
  1143 => (x"6f",x"4c",x"5f",x"32"),
  1144 => (x"20",x"20",x"3a",x"63"),
  1145 => (x"20",x"20",x"20",x"20"),
  1146 => (x"20",x"20",x"20",x"20"),
  1147 => (x"0a",x"73",x"25",x"20"),
  1148 => (x"00",x"00",x"00",x"00"),
  1149 => (x"20",x"20",x"20",x"20"),
  1150 => (x"20",x"20",x"20",x"20"),
  1151 => (x"75",x"6f",x"68",x"73"),
  1152 => (x"62",x"20",x"64",x"6c"),
  1153 => (x"20",x"20",x"3a",x"65"),
  1154 => (x"52",x"48",x"44",x"20"),
  1155 => (x"4f",x"54",x"53",x"59"),
  1156 => (x"50",x"20",x"45",x"4e"),
  1157 => (x"52",x"47",x"4f",x"52"),
  1158 => (x"20",x"2c",x"4d",x"41"),
  1159 => (x"44",x"4e",x"27",x"32"),
  1160 => (x"52",x"54",x"53",x"20"),
  1161 => (x"0a",x"47",x"4e",x"49"),
  1162 => (x"00",x"00",x"00",x"00"),
  1163 => (x"00",x"00",x"00",x"0a"),
  1164 => (x"72",x"65",x"73",x"55"),
  1165 => (x"6d",x"69",x"74",x"20"),
  1166 => (x"25",x"20",x"3a",x"65"),
  1167 => (x"1e",x"00",x"0a",x"64"),
  1168 => (x"66",x"c8",x"1e",x"73"),
  1169 => (x"49",x"66",x"cc",x"4b"),
  1170 => (x"ab",x"c2",x"79",x"73"),
  1171 => (x"c1",x"87",x"c4",x"05"),
  1172 => (x"c0",x"87",x"c2",x"4a"),
  1173 => (x"05",x"9a",x"72",x"4a"),
  1174 => (x"79",x"c3",x"87",x"c2"),
  1175 => (x"d8",x"02",x"ab",x"c0"),
  1176 => (x"02",x"ab",x"c1",x"87"),
  1177 => (x"ab",x"c2",x"87",x"d7"),
  1178 => (x"87",x"e5",x"c0",x"02"),
  1179 => (x"c0",x"02",x"ab",x"c3"),
  1180 => (x"ab",x"c4",x"87",x"e5"),
  1181 => (x"de",x"87",x"de",x"02"),
  1182 => (x"da",x"79",x"c0",x"87"),
  1183 => (x"f8",x"cf",x"c1",x"87"),
  1184 => (x"e4",x"c1",x"48",x"bf"),
  1185 => (x"c4",x"06",x"a8",x"b7"),
  1186 => (x"ca",x"79",x"c0",x"87"),
  1187 => (x"c6",x"79",x"c3",x"87"),
  1188 => (x"c2",x"79",x"c1",x"87"),
  1189 => (x"26",x"79",x"c2",x"87"),
  1190 => (x"1e",x"4f",x"26",x"4b"),
  1191 => (x"c2",x"49",x"66",x"c4"),
  1192 => (x"48",x"66",x"c8",x"81"),
  1193 => (x"66",x"cc",x"80",x"71"),
  1194 => (x"26",x"08",x"78",x"08"),
  1195 => (x"1e",x"73",x"1e",x"4f"),
  1196 => (x"1e",x"75",x"1e",x"74"),
  1197 => (x"e4",x"c0",x"86",x"f4"),
  1198 => (x"84",x"c5",x"4c",x"66"),
  1199 => (x"90",x"c4",x"48",x"74"),
  1200 => (x"dc",x"58",x"a6",x"c8"),
  1201 => (x"66",x"c4",x"48",x"66"),
  1202 => (x"58",x"a6",x"c4",x"80"),
  1203 => (x"e8",x"c0",x"48",x"6e"),
  1204 => (x"a6",x"c8",x"78",x"66"),
  1205 => (x"78",x"a4",x"c1",x"48"),
  1206 => (x"dc",x"91",x"c4",x"49"),
  1207 => (x"e8",x"c0",x"81",x"66"),
  1208 => (x"a4",x"de",x"79",x"66"),
  1209 => (x"dc",x"91",x"c4",x"49"),
  1210 => (x"79",x"74",x"81",x"66"),
  1211 => (x"ac",x"b7",x"66",x"c8"),
  1212 => (x"87",x"e0",x"c0",x"01"),
  1213 => (x"c8",x"c3",x"49",x"74"),
  1214 => (x"66",x"e0",x"c0",x"91"),
  1215 => (x"71",x"4d",x"c4",x"81"),
  1216 => (x"82",x"66",x"c4",x"4a"),
  1217 => (x"74",x"4b",x"66",x"c8"),
  1218 => (x"74",x"83",x"c1",x"8b"),
  1219 => (x"c1",x"82",x"75",x"7a"),
  1220 => (x"87",x"f7",x"01",x"8b"),
  1221 => (x"c8",x"c3",x"4a",x"74"),
  1222 => (x"66",x"e0",x"c0",x"92"),
  1223 => (x"c1",x"49",x"74",x"82"),
  1224 => (x"72",x"91",x"c4",x"89"),
  1225 => (x"48",x"69",x"49",x"a1"),
  1226 => (x"79",x"70",x"80",x"c1"),
  1227 => (x"c3",x"49",x"a4",x"d4"),
  1228 => (x"e0",x"c0",x"91",x"c8"),
  1229 => (x"66",x"c4",x"81",x"66"),
  1230 => (x"79",x"bf",x"6e",x"81"),
  1231 => (x"48",x"f8",x"cf",x"c1"),
  1232 => (x"8e",x"f4",x"78",x"c5"),
  1233 => (x"4c",x"26",x"4d",x"26"),
  1234 => (x"4f",x"26",x"4b",x"26"),
  1235 => (x"97",x"1e",x"73",x"1e"),
  1236 => (x"73",x"4b",x"66",x"c8"),
  1237 => (x"66",x"cc",x"97",x"4a"),
  1238 => (x"aa",x"b7",x"71",x"49"),
  1239 => (x"c0",x"87",x"c4",x"02"),
  1240 => (x"c1",x"87",x"c7",x"48"),
  1241 => (x"5b",x"97",x"c4",x"d0"),
  1242 => (x"4b",x"26",x"48",x"c1"),
  1243 => (x"73",x"1e",x"4f",x"26"),
  1244 => (x"75",x"1e",x"74",x"1e"),
  1245 => (x"c2",x"86",x"f8",x"1e"),
  1246 => (x"49",x"66",x"dc",x"4d"),
  1247 => (x"66",x"d8",x"81",x"c1"),
  1248 => (x"a1",x"84",x"c2",x"4c"),
  1249 => (x"49",x"6b",x"97",x"4b"),
  1250 => (x"7e",x"97",x"6c",x"97"),
  1251 => (x"71",x"4a",x"6e",x"97"),
  1252 => (x"c7",x"02",x"aa",x"b7"),
  1253 => (x"48",x"a6",x"c4",x"87"),
  1254 => (x"87",x"cc",x"78",x"c0"),
  1255 => (x"48",x"c0",x"d0",x"c1"),
  1256 => (x"c4",x"50",x"6e",x"97"),
  1257 => (x"78",x"c1",x"48",x"a6"),
  1258 => (x"c4",x"05",x"66",x"c4"),
  1259 => (x"83",x"85",x"c1",x"87"),
  1260 => (x"ad",x"b7",x"c2",x"84"),
  1261 => (x"87",x"cd",x"ff",x"06"),
  1262 => (x"dc",x"4a",x"66",x"d8"),
  1263 => (x"fd",x"fe",x"49",x"66"),
  1264 => (x"b7",x"c0",x"87",x"f2"),
  1265 => (x"87",x"cb",x"06",x"a8"),
  1266 => (x"48",x"f8",x"cf",x"c1"),
  1267 => (x"c1",x"78",x"a5",x"c7"),
  1268 => (x"c0",x"87",x"c2",x"48"),
  1269 => (x"26",x"8e",x"f8",x"48"),
  1270 => (x"26",x"4c",x"26",x"4d"),
  1271 => (x"26",x"4f",x"26",x"4b"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
