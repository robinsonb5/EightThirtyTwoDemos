
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"c9",x"01"),
     1 => (x"cf",x"03",x"87",x"cc"),
     2 => (x"87",x"fd",x"00",x"87"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"36",x"27",x"4f",x"00"),
     5 => (x"4f",x"00",x"00",x"00"),
     6 => (x"0e",x"1e",x"18",x"0e"),
     7 => (x"00",x"00",x"44",x"27"),
     8 => (x"48",x"26",x"0f",x"00"),
     9 => (x"08",x"26",x"80",x"ff"),
    10 => (x"c0",x"c0",x"c2",x"4f"),
    11 => (x"17",x"36",x"27",x"4e"),
    12 => (x"00",x"0f",x"00",x"00"),
    13 => (x"f0",x"c1",x"87",x"fd"),
    14 => (x"43",x"27",x"4e",x"c0"),
    15 => (x"0f",x"00",x"00",x"00"),
    16 => (x"4f",x"87",x"fd",x"00"),
    17 => (x"0e",x"1e",x"18",x"0e"),
    18 => (x"80",x"ff",x"48",x"26"),
    19 => (x"1e",x"4f",x"08",x"26"),
    20 => (x"ff",x"1e",x"1e",x"72"),
    21 => (x"48",x"6a",x"4a",x"c0"),
    22 => (x"c4",x"98",x"c0",x"c4"),
    23 => (x"02",x"6e",x"58",x"a6"),
    24 => (x"cc",x"87",x"f3",x"ff"),
    25 => (x"66",x"cc",x"7a",x"66"),
    26 => (x"4a",x"26",x"26",x"48"),
    27 => (x"5e",x"0e",x"4f",x"26"),
    28 => (x"5d",x"5c",x"5b",x"5a"),
    29 => (x"4b",x"66",x"d4",x"0e"),
    30 => (x"4c",x"13",x"4d",x"c0"),
    31 => (x"c0",x"02",x"9c",x"74"),
    32 => (x"4a",x"74",x"87",x"d6"),
    33 => (x"4f",x"27",x"1e",x"72"),
    34 => (x"0f",x"00",x"00",x"00"),
    35 => (x"85",x"c1",x"86",x"c4"),
    36 => (x"9c",x"74",x"4c",x"13"),
    37 => (x"87",x"ea",x"ff",x"05"),
    38 => (x"4d",x"26",x"48",x"75"),
    39 => (x"4b",x"26",x"4c",x"26"),
    40 => (x"4f",x"26",x"4a",x"26"),
    41 => (x"5b",x"5a",x"5e",x"0e"),
    42 => (x"c8",x"0e",x"5d",x"5c"),
    43 => (x"66",x"e0",x"c0",x"8e"),
    44 => (x"4c",x"66",x"dc",x"4d"),
    45 => (x"00",x"1b",x"28",x"27"),
    46 => (x"49",x"76",x"4b",x"00"),
    47 => (x"00",x"19",x"92",x"27"),
    48 => (x"a6",x"c4",x"79",x"00"),
    49 => (x"c0",x"79",x"c0",x"49"),
    50 => (x"c0",x"03",x"ac",x"b7"),
    51 => (x"ed",x"c0",x"87",x"cd"),
    52 => (x"00",x"4f",x"27",x"1e"),
    53 => (x"c4",x"0f",x"00",x"00"),
    54 => (x"74",x"8c",x"0c",x"86"),
    55 => (x"c6",x"c0",x"05",x"9c"),
    56 => (x"53",x"f0",x"c0",x"87"),
    57 => (x"74",x"87",x"f6",x"c0"),
    58 => (x"f0",x"c0",x"02",x"9c"),
    59 => (x"72",x"49",x"74",x"87"),
    60 => (x"66",x"e8",x"c0",x"1e"),
    61 => (x"19",x"48",x"27",x"4a"),
    62 => (x"26",x"0f",x"00",x"00"),
    63 => (x"72",x"4a",x"71",x"4a"),
    64 => (x"12",x"82",x"6e",x"4a"),
    65 => (x"72",x"49",x"74",x"53"),
    66 => (x"66",x"e8",x"c0",x"1e"),
    67 => (x"19",x"48",x"27",x"4a"),
    68 => (x"26",x"0f",x"00",x"00"),
    69 => (x"74",x"4c",x"70",x"4a"),
    70 => (x"d0",x"ff",x"05",x"9c"),
    71 => (x"1b",x"28",x"27",x"87"),
    72 => (x"ab",x"b7",x"00",x"00"),
    73 => (x"87",x"d8",x"c0",x"02"),
    74 => (x"6b",x"97",x"8b",x"c1"),
    75 => (x"48",x"66",x"c4",x"55"),
    76 => (x"a6",x"c8",x"80",x"c1"),
    77 => (x"1b",x"28",x"27",x"58"),
    78 => (x"ab",x"b7",x"00",x"00"),
    79 => (x"87",x"e8",x"ff",x"05"),
    80 => (x"66",x"c4",x"55",x"c0"),
    81 => (x"26",x"86",x"c8",x"48"),
    82 => (x"26",x"4c",x"26",x"4d"),
    83 => (x"26",x"4a",x"26",x"4b"),
    84 => (x"5a",x"5e",x"0e",x"4f"),
    85 => (x"0e",x"5d",x"5c",x"5b"),
    86 => (x"76",x"4c",x"c0",x"1e"),
    87 => (x"dc",x"79",x"c0",x"49"),
    88 => (x"66",x"d8",x"4b",x"a6"),
    89 => (x"48",x"66",x"d8",x"4a"),
    90 => (x"a6",x"dc",x"80",x"c1"),
    91 => (x"c1",x"4d",x"12",x"58"),
    92 => (x"c0",x"c0",x"c0",x"c0"),
    93 => (x"b7",x"c0",x"c4",x"95"),
    94 => (x"9d",x"75",x"4d",x"95"),
    95 => (x"87",x"d2",x"c4",x"02"),
    96 => (x"d7",x"c3",x"02",x"6e"),
    97 => (x"c0",x"49",x"76",x"87"),
    98 => (x"c1",x"4a",x"75",x"79"),
    99 => (x"c2",x"02",x"ad",x"e3"),
   100 => (x"e4",x"c1",x"87",x"dd"),
   101 => (x"d8",x"c0",x"02",x"aa"),
   102 => (x"aa",x"ec",x"c1",x"87"),
   103 => (x"87",x"c8",x"c2",x"02"),
   104 => (x"02",x"aa",x"f3",x"c1"),
   105 => (x"c1",x"87",x"e8",x"c1"),
   106 => (x"c0",x"02",x"aa",x"f8"),
   107 => (x"d3",x"c2",x"87",x"f2"),
   108 => (x"27",x"1e",x"ca",x"87"),
   109 => (x"00",x"00",x"1b",x"78"),
   110 => (x"73",x"83",x"c4",x"1e"),
   111 => (x"6a",x"8a",x"c4",x"4a"),
   112 => (x"00",x"a4",x"27",x"1e"),
   113 => (x"cc",x"0f",x"00",x"00"),
   114 => (x"74",x"4a",x"70",x"86"),
   115 => (x"27",x"84",x"72",x"4c"),
   116 => (x"00",x"00",x"1b",x"78"),
   117 => (x"00",x"6e",x"27",x"1e"),
   118 => (x"c4",x"0f",x"00",x"00"),
   119 => (x"87",x"d4",x"c2",x"86"),
   120 => (x"78",x"27",x"1e",x"d0"),
   121 => (x"1e",x"00",x"00",x"1b"),
   122 => (x"4a",x"73",x"83",x"c4"),
   123 => (x"1e",x"6a",x"8a",x"c4"),
   124 => (x"00",x"00",x"a4",x"27"),
   125 => (x"86",x"cc",x"0f",x"00"),
   126 => (x"4c",x"74",x"4a",x"70"),
   127 => (x"78",x"27",x"84",x"72"),
   128 => (x"1e",x"00",x"00",x"1b"),
   129 => (x"00",x"00",x"6e",x"27"),
   130 => (x"86",x"c4",x"0f",x"00"),
   131 => (x"c4",x"87",x"e5",x"c1"),
   132 => (x"c4",x"4a",x"73",x"83"),
   133 => (x"27",x"1e",x"6a",x"8a"),
   134 => (x"00",x"00",x"00",x"6e"),
   135 => (x"70",x"86",x"c4",x"0f"),
   136 => (x"72",x"4c",x"74",x"4a"),
   137 => (x"87",x"cc",x"c1",x"84"),
   138 => (x"79",x"c1",x"49",x"76"),
   139 => (x"c4",x"87",x"c5",x"c1"),
   140 => (x"c4",x"4a",x"73",x"83"),
   141 => (x"27",x"1e",x"6a",x"8a"),
   142 => (x"00",x"00",x"00",x"4f"),
   143 => (x"c1",x"86",x"c4",x"0f"),
   144 => (x"87",x"f0",x"c0",x"84"),
   145 => (x"27",x"1e",x"e5",x"c0"),
   146 => (x"00",x"00",x"00",x"4f"),
   147 => (x"75",x"86",x"c4",x"0f"),
   148 => (x"00",x"4f",x"27",x"1e"),
   149 => (x"c4",x"0f",x"00",x"00"),
   150 => (x"87",x"d8",x"c0",x"86"),
   151 => (x"05",x"ad",x"e5",x"c0"),
   152 => (x"76",x"87",x"c7",x"c0"),
   153 => (x"c0",x"79",x"c1",x"49"),
   154 => (x"1e",x"75",x"87",x"ca"),
   155 => (x"00",x"00",x"4f",x"27"),
   156 => (x"86",x"c4",x"0f",x"00"),
   157 => (x"d8",x"4a",x"66",x"d8"),
   158 => (x"80",x"c1",x"48",x"66"),
   159 => (x"12",x"58",x"a6",x"dc"),
   160 => (x"c0",x"c0",x"c1",x"4d"),
   161 => (x"c4",x"95",x"c0",x"c0"),
   162 => (x"4d",x"95",x"b7",x"c0"),
   163 => (x"fb",x"05",x"9d",x"75"),
   164 => (x"48",x"74",x"87",x"ee"),
   165 => (x"26",x"4d",x"26",x"26"),
   166 => (x"26",x"4b",x"26",x"4c"),
   167 => (x"0e",x"4f",x"26",x"4a"),
   168 => (x"5c",x"5b",x"5a",x"5e"),
   169 => (x"8e",x"e4",x"c0",x"0e"),
   170 => (x"ff",x"4c",x"ff",x"c3"),
   171 => (x"7b",x"74",x"4b",x"d4"),
   172 => (x"9a",x"74",x"4a",x"6b"),
   173 => (x"48",x"6b",x"7b",x"74"),
   174 => (x"a6",x"c4",x"98",x"74"),
   175 => (x"c8",x"48",x"6e",x"58"),
   176 => (x"58",x"a6",x"c8",x"30"),
   177 => (x"72",x"49",x"a6",x"c8"),
   178 => (x"c4",x"4a",x"72",x"79"),
   179 => (x"7b",x"74",x"b2",x"66"),
   180 => (x"98",x"74",x"48",x"6b"),
   181 => (x"cc",x"58",x"a6",x"d0"),
   182 => (x"30",x"d0",x"48",x"66"),
   183 => (x"d4",x"58",x"a6",x"d4"),
   184 => (x"79",x"72",x"49",x"a6"),
   185 => (x"66",x"d0",x"4a",x"72"),
   186 => (x"6b",x"7b",x"74",x"b2"),
   187 => (x"dc",x"98",x"74",x"48"),
   188 => (x"66",x"d8",x"58",x"a6"),
   189 => (x"c0",x"30",x"d8",x"48"),
   190 => (x"c0",x"58",x"a6",x"e0"),
   191 => (x"72",x"49",x"a6",x"e0"),
   192 => (x"dc",x"4a",x"72",x"79"),
   193 => (x"48",x"72",x"b2",x"66"),
   194 => (x"26",x"86",x"e4",x"c0"),
   195 => (x"26",x"4b",x"26",x"4c"),
   196 => (x"0e",x"4f",x"26",x"4a"),
   197 => (x"5c",x"5b",x"5a",x"5e"),
   198 => (x"c3",x"8e",x"d8",x"0e"),
   199 => (x"d4",x"ff",x"4c",x"ff"),
   200 => (x"6b",x"7b",x"74",x"4b"),
   201 => (x"74",x"9a",x"74",x"4a"),
   202 => (x"6b",x"32",x"c8",x"7b"),
   203 => (x"c4",x"98",x"74",x"48"),
   204 => (x"a6",x"c4",x"58",x"a6"),
   205 => (x"72",x"79",x"72",x"49"),
   206 => (x"74",x"b2",x"6e",x"4a"),
   207 => (x"6b",x"32",x"c8",x"7b"),
   208 => (x"cc",x"98",x"74",x"48"),
   209 => (x"a6",x"cc",x"58",x"a6"),
   210 => (x"72",x"79",x"72",x"49"),
   211 => (x"b2",x"66",x"c8",x"4a"),
   212 => (x"32",x"c8",x"7b",x"74"),
   213 => (x"98",x"74",x"48",x"6b"),
   214 => (x"d4",x"58",x"a6",x"d4"),
   215 => (x"79",x"72",x"49",x"a6"),
   216 => (x"66",x"d0",x"4a",x"72"),
   217 => (x"d8",x"48",x"72",x"b2"),
   218 => (x"26",x"4c",x"26",x"86"),
   219 => (x"26",x"4a",x"26",x"4b"),
   220 => (x"5a",x"5e",x"0e",x"4f"),
   221 => (x"0e",x"5d",x"5c",x"5b"),
   222 => (x"d4",x"4d",x"d4",x"ff"),
   223 => (x"ff",x"c3",x"48",x"66"),
   224 => (x"27",x"7d",x"70",x"98"),
   225 => (x"00",x"00",x"1b",x"9c"),
   226 => (x"c8",x"c0",x"05",x"bf"),
   227 => (x"48",x"66",x"d8",x"87"),
   228 => (x"a6",x"dc",x"30",x"c9"),
   229 => (x"4a",x"66",x"d8",x"58"),
   230 => (x"48",x"72",x"2a",x"d8"),
   231 => (x"70",x"98",x"ff",x"c3"),
   232 => (x"4a",x"66",x"d8",x"7d"),
   233 => (x"48",x"72",x"2a",x"d0"),
   234 => (x"70",x"98",x"ff",x"c3"),
   235 => (x"4a",x"66",x"d8",x"7d"),
   236 => (x"48",x"72",x"2a",x"c8"),
   237 => (x"70",x"98",x"ff",x"c3"),
   238 => (x"48",x"66",x"d8",x"7d"),
   239 => (x"70",x"98",x"ff",x"c3"),
   240 => (x"4a",x"66",x"d4",x"7d"),
   241 => (x"48",x"72",x"2a",x"d0"),
   242 => (x"70",x"98",x"ff",x"c3"),
   243 => (x"c3",x"4c",x"6d",x"7d"),
   244 => (x"f0",x"c9",x"9c",x"ff"),
   245 => (x"ff",x"c3",x"4b",x"ff"),
   246 => (x"c0",x"05",x"ac",x"b7"),
   247 => (x"ff",x"c3",x"87",x"d8"),
   248 => (x"6d",x"7d",x"72",x"4a"),
   249 => (x"c1",x"9c",x"72",x"4c"),
   250 => (x"02",x"9b",x"73",x"8b"),
   251 => (x"72",x"87",x"c7",x"c0"),
   252 => (x"ff",x"02",x"ac",x"b7"),
   253 => (x"48",x"74",x"87",x"eb"),
   254 => (x"4c",x"26",x"4d",x"26"),
   255 => (x"4a",x"26",x"4b",x"26"),
   256 => (x"72",x"1e",x"4f",x"26"),
   257 => (x"ff",x"4a",x"c0",x"1e"),
   258 => (x"ff",x"c3",x"49",x"d4"),
   259 => (x"c3",x"82",x"c1",x"79"),
   260 => (x"04",x"aa",x"b7",x"c8"),
   261 => (x"26",x"87",x"f0",x"ff"),
   262 => (x"0e",x"4f",x"26",x"4a"),
   263 => (x"5c",x"5b",x"5a",x"5e"),
   264 => (x"ff",x"c0",x"0e",x"5d"),
   265 => (x"4d",x"f7",x"c1",x"f0"),
   266 => (x"c0",x"c0",x"c0",x"c1"),
   267 => (x"27",x"4b",x"c0",x"c0"),
   268 => (x"00",x"00",x"04",x"02"),
   269 => (x"df",x"f8",x"c4",x"0f"),
   270 => (x"75",x"1e",x"c0",x"4c"),
   271 => (x"03",x"71",x"27",x"1e"),
   272 => (x"c8",x"0f",x"00",x"00"),
   273 => (x"c1",x"4a",x"70",x"86"),
   274 => (x"c0",x"05",x"aa",x"b7"),
   275 => (x"d4",x"ff",x"87",x"ef"),
   276 => (x"79",x"ff",x"c3",x"49"),
   277 => (x"e1",x"c0",x"1e",x"73"),
   278 => (x"1e",x"e9",x"c1",x"f0"),
   279 => (x"00",x"03",x"71",x"27"),
   280 => (x"86",x"c8",x"0f",x"00"),
   281 => (x"9a",x"72",x"4a",x"70"),
   282 => (x"87",x"cb",x"c0",x"05"),
   283 => (x"c3",x"49",x"d4",x"ff"),
   284 => (x"48",x"c1",x"79",x"ff"),
   285 => (x"27",x"87",x"d0",x"c0"),
   286 => (x"00",x"00",x"04",x"02"),
   287 => (x"74",x"8c",x"c1",x"0f"),
   288 => (x"f4",x"fe",x"05",x"9c"),
   289 => (x"26",x"48",x"c0",x"87"),
   290 => (x"26",x"4c",x"26",x"4d"),
   291 => (x"26",x"4a",x"26",x"4b"),
   292 => (x"5a",x"5e",x"0e",x"4f"),
   293 => (x"c0",x"0e",x"5c",x"5b"),
   294 => (x"c1",x"c1",x"f0",x"ff"),
   295 => (x"49",x"d4",x"ff",x"4c"),
   296 => (x"27",x"79",x"ff",x"c3"),
   297 => (x"00",x"00",x"19",x"a3"),
   298 => (x"00",x"6e",x"27",x"1e"),
   299 => (x"c4",x"0f",x"00",x"00"),
   300 => (x"c0",x"4b",x"d3",x"86"),
   301 => (x"27",x"1e",x"74",x"1e"),
   302 => (x"00",x"00",x"03",x"71"),
   303 => (x"70",x"86",x"c8",x"0f"),
   304 => (x"05",x"9a",x"72",x"4a"),
   305 => (x"ff",x"87",x"cb",x"c0"),
   306 => (x"ff",x"c3",x"49",x"d4"),
   307 => (x"c0",x"48",x"c1",x"79"),
   308 => (x"02",x"27",x"87",x"d0"),
   309 => (x"0f",x"00",x"00",x"04"),
   310 => (x"9b",x"73",x"8b",x"c1"),
   311 => (x"87",x"d3",x"ff",x"05"),
   312 => (x"4c",x"26",x"48",x"c0"),
   313 => (x"4a",x"26",x"4b",x"26"),
   314 => (x"5e",x"0e",x"4f",x"26"),
   315 => (x"5d",x"5c",x"5b",x"5a"),
   316 => (x"ff",x"c3",x"1e",x"0e"),
   317 => (x"4c",x"d4",x"ff",x"4d"),
   318 => (x"00",x"04",x"02",x"27"),
   319 => (x"ea",x"c6",x"0f",x"00"),
   320 => (x"f0",x"e1",x"c0",x"1e"),
   321 => (x"27",x"1e",x"c8",x"c1"),
   322 => (x"00",x"00",x"03",x"71"),
   323 => (x"70",x"86",x"c8",x"0f"),
   324 => (x"27",x"1e",x"72",x"4a"),
   325 => (x"00",x"00",x"06",x"49"),
   326 => (x"01",x"51",x"27",x"1e"),
   327 => (x"c8",x"0f",x"00",x"00"),
   328 => (x"aa",x"b7",x"c1",x"86"),
   329 => (x"87",x"cb",x"c0",x"02"),
   330 => (x"00",x"04",x"91",x"27"),
   331 => (x"48",x"c0",x"0f",x"00"),
   332 => (x"27",x"87",x"c9",x"c3"),
   333 => (x"00",x"00",x"03",x"13"),
   334 => (x"cf",x"4a",x"70",x"0f"),
   335 => (x"c6",x"9a",x"ff",x"ff"),
   336 => (x"02",x"aa",x"b7",x"ea"),
   337 => (x"27",x"87",x"cb",x"c0"),
   338 => (x"00",x"00",x"04",x"91"),
   339 => (x"c2",x"48",x"c0",x"0f"),
   340 => (x"7c",x"75",x"87",x"ea"),
   341 => (x"f1",x"c0",x"49",x"76"),
   342 => (x"04",x"1b",x"27",x"79"),
   343 => (x"70",x"0f",x"00",x"00"),
   344 => (x"02",x"9a",x"72",x"4a"),
   345 => (x"c0",x"87",x"eb",x"c1"),
   346 => (x"f0",x"ff",x"c0",x"1e"),
   347 => (x"27",x"1e",x"fa",x"c1"),
   348 => (x"00",x"00",x"03",x"71"),
   349 => (x"70",x"86",x"c8",x"0f"),
   350 => (x"05",x"9b",x"73",x"4b"),
   351 => (x"73",x"87",x"c3",x"c1"),
   352 => (x"06",x"07",x"27",x"1e"),
   353 => (x"27",x"1e",x"00",x"00"),
   354 => (x"00",x"00",x"01",x"51"),
   355 => (x"75",x"86",x"c8",x"0f"),
   356 => (x"75",x"4b",x"6c",x"7c"),
   357 => (x"27",x"1e",x"73",x"9b"),
   358 => (x"00",x"00",x"06",x"13"),
   359 => (x"01",x"51",x"27",x"1e"),
   360 => (x"c8",x"0f",x"00",x"00"),
   361 => (x"75",x"7c",x"75",x"86"),
   362 => (x"75",x"7c",x"75",x"7c"),
   363 => (x"c1",x"4a",x"73",x"7c"),
   364 => (x"9a",x"72",x"9a",x"c0"),
   365 => (x"87",x"c5",x"c0",x"02"),
   366 => (x"ff",x"c0",x"48",x"c1"),
   367 => (x"c0",x"48",x"c0",x"87"),
   368 => (x"1e",x"73",x"87",x"fa"),
   369 => (x"00",x"06",x"21",x"27"),
   370 => (x"51",x"27",x"1e",x"00"),
   371 => (x"0f",x"00",x"00",x"01"),
   372 => (x"49",x"6e",x"86",x"c8"),
   373 => (x"05",x"a9",x"b7",x"c2"),
   374 => (x"27",x"87",x"d3",x"c0"),
   375 => (x"00",x"00",x"06",x"2d"),
   376 => (x"01",x"51",x"27",x"1e"),
   377 => (x"c4",x"0f",x"00",x"00"),
   378 => (x"c0",x"48",x"c0",x"86"),
   379 => (x"48",x"6e",x"87",x"ce"),
   380 => (x"a6",x"c4",x"88",x"c1"),
   381 => (x"fd",x"05",x"6e",x"58"),
   382 => (x"48",x"c0",x"87",x"df"),
   383 => (x"26",x"4d",x"26",x"26"),
   384 => (x"26",x"4b",x"26",x"4c"),
   385 => (x"43",x"4f",x"26",x"4a"),
   386 => (x"38",x"35",x"44",x"4d"),
   387 => (x"0a",x"64",x"25",x"20"),
   388 => (x"43",x"00",x"20",x"20"),
   389 => (x"38",x"35",x"44",x"4d"),
   390 => (x"25",x"20",x"32",x"5f"),
   391 => (x"20",x"20",x"0a",x"64"),
   392 => (x"44",x"4d",x"43",x"00"),
   393 => (x"25",x"20",x"38",x"35"),
   394 => (x"20",x"20",x"0a",x"64"),
   395 => (x"48",x"44",x"53",x"00"),
   396 => (x"6e",x"49",x"20",x"43"),
   397 => (x"61",x"69",x"74",x"69"),
   398 => (x"61",x"7a",x"69",x"6c"),
   399 => (x"6e",x"6f",x"69",x"74"),
   400 => (x"72",x"72",x"65",x"20"),
   401 => (x"0a",x"21",x"72",x"6f"),
   402 => (x"64",x"6d",x"63",x"00"),
   403 => (x"44",x"4d",x"43",x"5f"),
   404 => (x"65",x"72",x"20",x"38"),
   405 => (x"6e",x"6f",x"70",x"73"),
   406 => (x"20",x"3a",x"65",x"73"),
   407 => (x"00",x"0a",x"64",x"25"),
   408 => (x"5b",x"5a",x"5e",x"0e"),
   409 => (x"1e",x"0e",x"5d",x"5c"),
   410 => (x"c8",x"4c",x"d0",x"ff"),
   411 => (x"27",x"4b",x"c0",x"c0"),
   412 => (x"00",x"00",x"1b",x"9c"),
   413 => (x"27",x"79",x"c1",x"49"),
   414 => (x"00",x"00",x"07",x"7d"),
   415 => (x"00",x"6e",x"27",x"1e"),
   416 => (x"c4",x"0f",x"00",x"00"),
   417 => (x"6c",x"4d",x"c7",x"86"),
   418 => (x"c4",x"98",x"73",x"48"),
   419 => (x"02",x"6e",x"58",x"a6"),
   420 => (x"6c",x"87",x"cc",x"c0"),
   421 => (x"c4",x"98",x"73",x"48"),
   422 => (x"05",x"6e",x"58",x"a6"),
   423 => (x"c0",x"87",x"f4",x"ff"),
   424 => (x"04",x"02",x"27",x"7c"),
   425 => (x"6c",x"0f",x"00",x"00"),
   426 => (x"c4",x"98",x"73",x"48"),
   427 => (x"02",x"6e",x"58",x"a6"),
   428 => (x"6c",x"87",x"cc",x"c0"),
   429 => (x"c4",x"98",x"73",x"48"),
   430 => (x"05",x"6e",x"58",x"a6"),
   431 => (x"c1",x"87",x"f4",x"ff"),
   432 => (x"c0",x"1e",x"c0",x"7c"),
   433 => (x"c0",x"c1",x"d0",x"e5"),
   434 => (x"03",x"71",x"27",x"1e"),
   435 => (x"c8",x"0f",x"00",x"00"),
   436 => (x"c1",x"4a",x"70",x"86"),
   437 => (x"c0",x"05",x"aa",x"b7"),
   438 => (x"4d",x"c1",x"87",x"c2"),
   439 => (x"05",x"ad",x"b7",x"c2"),
   440 => (x"27",x"87",x"d3",x"c0"),
   441 => (x"00",x"00",x"07",x"78"),
   442 => (x"00",x"6e",x"27",x"1e"),
   443 => (x"c4",x"0f",x"00",x"00"),
   444 => (x"c1",x"48",x"c0",x"86"),
   445 => (x"8d",x"c1",x"87",x"f7"),
   446 => (x"fe",x"05",x"9d",x"75"),
   447 => (x"ea",x"27",x"87",x"c9"),
   448 => (x"0f",x"00",x"00",x"04"),
   449 => (x"00",x"1b",x"a0",x"27"),
   450 => (x"9c",x"27",x"58",x"00"),
   451 => (x"bf",x"00",x"00",x"1b"),
   452 => (x"87",x"d0",x"c0",x"05"),
   453 => (x"ff",x"c0",x"1e",x"c1"),
   454 => (x"1e",x"d0",x"c1",x"f0"),
   455 => (x"00",x"03",x"71",x"27"),
   456 => (x"86",x"c8",x"0f",x"00"),
   457 => (x"c3",x"49",x"d4",x"ff"),
   458 => (x"13",x"27",x"79",x"ff"),
   459 => (x"0f",x"00",x"00",x"0a"),
   460 => (x"00",x"1b",x"a4",x"27"),
   461 => (x"a0",x"27",x"58",x"00"),
   462 => (x"bf",x"00",x"00",x"1b"),
   463 => (x"07",x"81",x"27",x"1e"),
   464 => (x"27",x"1e",x"00",x"00"),
   465 => (x"00",x"00",x"01",x"51"),
   466 => (x"6c",x"86",x"c8",x"0f"),
   467 => (x"c4",x"98",x"73",x"48"),
   468 => (x"02",x"6e",x"58",x"a6"),
   469 => (x"6c",x"87",x"cc",x"c0"),
   470 => (x"c4",x"98",x"73",x"48"),
   471 => (x"05",x"6e",x"58",x"a6"),
   472 => (x"c0",x"87",x"f4",x"ff"),
   473 => (x"49",x"d4",x"ff",x"7c"),
   474 => (x"c1",x"79",x"ff",x"c3"),
   475 => (x"4d",x"26",x"26",x"48"),
   476 => (x"4b",x"26",x"4c",x"26"),
   477 => (x"4f",x"26",x"4a",x"26"),
   478 => (x"52",x"52",x"45",x"49"),
   479 => (x"49",x"50",x"53",x"00"),
   480 => (x"20",x"44",x"53",x"00"),
   481 => (x"64",x"72",x"61",x"63"),
   482 => (x"7a",x"69",x"73",x"20"),
   483 => (x"73",x"69",x"20",x"65"),
   484 => (x"0a",x"64",x"25",x"20"),
   485 => (x"5a",x"5e",x"0e",x"00"),
   486 => (x"0e",x"5d",x"5c",x"5b"),
   487 => (x"4d",x"ff",x"c3",x"1e"),
   488 => (x"75",x"4c",x"d4",x"ff"),
   489 => (x"bf",x"d0",x"ff",x"7c"),
   490 => (x"c0",x"c0",x"c8",x"48"),
   491 => (x"58",x"a6",x"c4",x"98"),
   492 => (x"d2",x"c0",x"02",x"6e"),
   493 => (x"c0",x"c0",x"c8",x"87"),
   494 => (x"bf",x"d0",x"ff",x"4a"),
   495 => (x"c4",x"98",x"72",x"48"),
   496 => (x"05",x"6e",x"58",x"a6"),
   497 => (x"ff",x"87",x"f2",x"ff"),
   498 => (x"c1",x"c4",x"49",x"d0"),
   499 => (x"d8",x"7c",x"75",x"79"),
   500 => (x"ff",x"c0",x"1e",x"66"),
   501 => (x"1e",x"d8",x"c1",x"f0"),
   502 => (x"00",x"03",x"71",x"27"),
   503 => (x"86",x"c8",x"0f",x"00"),
   504 => (x"9a",x"72",x"4a",x"70"),
   505 => (x"87",x"d3",x"c0",x"02"),
   506 => (x"00",x"08",x"9d",x"27"),
   507 => (x"6e",x"27",x"1e",x"00"),
   508 => (x"0f",x"00",x"00",x"00"),
   509 => (x"48",x"c1",x"86",x"c4"),
   510 => (x"75",x"87",x"d7",x"c2"),
   511 => (x"7c",x"fe",x"c3",x"7c"),
   512 => (x"79",x"c0",x"49",x"76"),
   513 => (x"4a",x"bf",x"66",x"dc"),
   514 => (x"b7",x"d8",x"4b",x"72"),
   515 => (x"75",x"48",x"73",x"2b"),
   516 => (x"72",x"7c",x"70",x"98"),
   517 => (x"2b",x"b7",x"d0",x"4b"),
   518 => (x"98",x"75",x"48",x"73"),
   519 => (x"4b",x"72",x"7c",x"70"),
   520 => (x"73",x"2b",x"b7",x"c8"),
   521 => (x"70",x"98",x"75",x"48"),
   522 => (x"75",x"48",x"72",x"7c"),
   523 => (x"dc",x"7c",x"70",x"98"),
   524 => (x"80",x"c4",x"48",x"66"),
   525 => (x"58",x"a6",x"e0",x"c0"),
   526 => (x"80",x"c1",x"48",x"6e"),
   527 => (x"6e",x"58",x"a6",x"c4"),
   528 => (x"b7",x"c0",x"c2",x"49"),
   529 => (x"fb",x"fe",x"04",x"a9"),
   530 => (x"75",x"7c",x"75",x"87"),
   531 => (x"d8",x"7c",x"75",x"7c"),
   532 => (x"75",x"4b",x"e0",x"da"),
   533 => (x"75",x"4a",x"6c",x"7c"),
   534 => (x"05",x"9a",x"72",x"9a"),
   535 => (x"c1",x"87",x"c8",x"c0"),
   536 => (x"05",x"9b",x"73",x"8b"),
   537 => (x"75",x"87",x"ec",x"ff"),
   538 => (x"bf",x"d0",x"ff",x"7c"),
   539 => (x"c0",x"c0",x"c8",x"48"),
   540 => (x"58",x"a6",x"c4",x"98"),
   541 => (x"d2",x"c0",x"02",x"6e"),
   542 => (x"c0",x"c0",x"c8",x"87"),
   543 => (x"bf",x"d0",x"ff",x"4a"),
   544 => (x"c4",x"98",x"72",x"48"),
   545 => (x"05",x"6e",x"58",x"a6"),
   546 => (x"ff",x"87",x"f2",x"ff"),
   547 => (x"79",x"c0",x"49",x"d0"),
   548 => (x"26",x"26",x"48",x"c0"),
   549 => (x"26",x"4c",x"26",x"4d"),
   550 => (x"26",x"4a",x"26",x"4b"),
   551 => (x"69",x"72",x"57",x"4f"),
   552 => (x"66",x"20",x"65",x"74"),
   553 => (x"65",x"6c",x"69",x"61"),
   554 => (x"0e",x"00",x"0a",x"64"),
   555 => (x"5c",x"5b",x"5a",x"5e"),
   556 => (x"d8",x"1e",x"0e",x"5d"),
   557 => (x"66",x"dc",x"4c",x"66"),
   558 => (x"c0",x"49",x"76",x"4b"),
   559 => (x"cd",x"ee",x"c5",x"79"),
   560 => (x"d4",x"ff",x"4d",x"df"),
   561 => (x"79",x"ff",x"c3",x"49"),
   562 => (x"4a",x"bf",x"d4",x"ff"),
   563 => (x"c3",x"9a",x"ff",x"c3"),
   564 => (x"05",x"aa",x"b7",x"fe"),
   565 => (x"27",x"87",x"e5",x"c1"),
   566 => (x"00",x"00",x"1b",x"98"),
   567 => (x"c4",x"79",x"c0",x"49"),
   568 => (x"c0",x"04",x"ab",x"b7"),
   569 => (x"9f",x"27",x"87",x"e4"),
   570 => (x"0f",x"00",x"00",x"02"),
   571 => (x"7c",x"72",x"4a",x"70"),
   572 => (x"98",x"27",x"84",x"c4"),
   573 => (x"bf",x"00",x"00",x"1b"),
   574 => (x"27",x"80",x"72",x"48"),
   575 => (x"00",x"00",x"1b",x"9c"),
   576 => (x"c4",x"8b",x"c4",x"58"),
   577 => (x"ff",x"03",x"ab",x"b7"),
   578 => (x"b7",x"c0",x"87",x"dc"),
   579 => (x"e5",x"c0",x"06",x"ab"),
   580 => (x"4d",x"d4",x"ff",x"87"),
   581 => (x"6d",x"7d",x"ff",x"c3"),
   582 => (x"7c",x"97",x"72",x"4a"),
   583 => (x"98",x"27",x"84",x"c1"),
   584 => (x"bf",x"00",x"00",x"1b"),
   585 => (x"27",x"80",x"72",x"48"),
   586 => (x"00",x"00",x"1b",x"9c"),
   587 => (x"c0",x"8b",x"c1",x"58"),
   588 => (x"ff",x"01",x"ab",x"b7"),
   589 => (x"4d",x"c1",x"87",x"de"),
   590 => (x"79",x"c1",x"49",x"76"),
   591 => (x"9d",x"75",x"8d",x"c1"),
   592 => (x"87",x"fe",x"fd",x"05"),
   593 => (x"c3",x"49",x"d4",x"ff"),
   594 => (x"48",x"6e",x"79",x"ff"),
   595 => (x"26",x"4d",x"26",x"26"),
   596 => (x"26",x"4b",x"26",x"4c"),
   597 => (x"0e",x"4f",x"26",x"4a"),
   598 => (x"5c",x"5b",x"5a",x"5e"),
   599 => (x"ff",x"1e",x"0e",x"5d"),
   600 => (x"c0",x"c8",x"4b",x"d0"),
   601 => (x"4c",x"c0",x"4a",x"c0"),
   602 => (x"c3",x"49",x"d4",x"ff"),
   603 => (x"48",x"6b",x"79",x"ff"),
   604 => (x"a6",x"c4",x"98",x"72"),
   605 => (x"c0",x"02",x"6e",x"58"),
   606 => (x"48",x"6b",x"87",x"cc"),
   607 => (x"a6",x"c4",x"98",x"72"),
   608 => (x"ff",x"05",x"6e",x"58"),
   609 => (x"c1",x"c4",x"87",x"f4"),
   610 => (x"49",x"d4",x"ff",x"7b"),
   611 => (x"d8",x"79",x"ff",x"c3"),
   612 => (x"ff",x"c0",x"1e",x"66"),
   613 => (x"1e",x"d1",x"c1",x"f0"),
   614 => (x"00",x"03",x"71",x"27"),
   615 => (x"86",x"c8",x"0f",x"00"),
   616 => (x"9d",x"75",x"4d",x"70"),
   617 => (x"87",x"d6",x"c0",x"02"),
   618 => (x"66",x"dc",x"1e",x"75"),
   619 => (x"09",x"f3",x"27",x"1e"),
   620 => (x"27",x"1e",x"00",x"00"),
   621 => (x"00",x"00",x"01",x"51"),
   622 => (x"c0",x"86",x"cc",x"0f"),
   623 => (x"c0",x"c8",x"87",x"e8"),
   624 => (x"66",x"e0",x"c0",x"1e"),
   625 => (x"87",x"e3",x"fb",x"1e"),
   626 => (x"4c",x"70",x"86",x"c8"),
   627 => (x"98",x"72",x"48",x"6b"),
   628 => (x"6e",x"58",x"a6",x"c4"),
   629 => (x"87",x"cc",x"c0",x"02"),
   630 => (x"98",x"72",x"48",x"6b"),
   631 => (x"6e",x"58",x"a6",x"c4"),
   632 => (x"87",x"f4",x"ff",x"05"),
   633 => (x"48",x"74",x"7b",x"c0"),
   634 => (x"26",x"4d",x"26",x"26"),
   635 => (x"26",x"4b",x"26",x"4c"),
   636 => (x"52",x"4f",x"26",x"4a"),
   637 => (x"20",x"64",x"61",x"65"),
   638 => (x"6d",x"6d",x"6f",x"63"),
   639 => (x"20",x"64",x"6e",x"61"),
   640 => (x"6c",x"69",x"61",x"66"),
   641 => (x"61",x"20",x"64",x"65"),
   642 => (x"64",x"25",x"20",x"74"),
   643 => (x"64",x"25",x"28",x"20"),
   644 => (x"0e",x"00",x"0a",x"29"),
   645 => (x"5c",x"5b",x"5a",x"5e"),
   646 => (x"c0",x"1e",x"0e",x"5d"),
   647 => (x"f0",x"ff",x"c0",x"1e"),
   648 => (x"27",x"1e",x"c9",x"c1"),
   649 => (x"00",x"00",x"03",x"71"),
   650 => (x"d2",x"86",x"c8",x"0f"),
   651 => (x"1b",x"b0",x"27",x"1e"),
   652 => (x"f9",x"1e",x"00",x"00"),
   653 => (x"86",x"c8",x"87",x"f5"),
   654 => (x"85",x"c1",x"4d",x"c0"),
   655 => (x"04",x"ad",x"b7",x"d2"),
   656 => (x"27",x"87",x"f7",x"ff"),
   657 => (x"00",x"00",x"1b",x"b0"),
   658 => (x"c3",x"4a",x"bf",x"97"),
   659 => (x"c0",x"c1",x"9a",x"c0"),
   660 => (x"c0",x"05",x"aa",x"b7"),
   661 => (x"b7",x"27",x"87",x"f2"),
   662 => (x"97",x"00",x"00",x"1b"),
   663 => (x"32",x"d0",x"4a",x"bf"),
   664 => (x"00",x"1b",x"b8",x"27"),
   665 => (x"4b",x"bf",x"97",x"00"),
   666 => (x"4a",x"72",x"33",x"c8"),
   667 => (x"b9",x"27",x"b2",x"73"),
   668 => (x"97",x"00",x"00",x"1b"),
   669 => (x"4a",x"72",x"4b",x"bf"),
   670 => (x"ff",x"cf",x"b2",x"73"),
   671 => (x"72",x"9a",x"ff",x"ff"),
   672 => (x"ca",x"85",x"c1",x"4d"),
   673 => (x"87",x"cb",x"c3",x"35"),
   674 => (x"00",x"1b",x"b9",x"27"),
   675 => (x"4a",x"bf",x"97",x"00"),
   676 => (x"9a",x"c6",x"32",x"c1"),
   677 => (x"00",x"1b",x"ba",x"27"),
   678 => (x"4b",x"bf",x"97",x"00"),
   679 => (x"72",x"2b",x"b7",x"c7"),
   680 => (x"27",x"b2",x"73",x"4a"),
   681 => (x"00",x"00",x"1b",x"b5"),
   682 => (x"73",x"4b",x"bf",x"97"),
   683 => (x"c4",x"98",x"cf",x"48"),
   684 => (x"b6",x"27",x"58",x"a6"),
   685 => (x"97",x"00",x"00",x"1b"),
   686 => (x"9b",x"c3",x"4b",x"bf"),
   687 => (x"b7",x"27",x"33",x"ca"),
   688 => (x"97",x"00",x"00",x"1b"),
   689 => (x"34",x"c2",x"4c",x"bf"),
   690 => (x"b3",x"74",x"4b",x"73"),
   691 => (x"00",x"1b",x"b8",x"27"),
   692 => (x"4c",x"bf",x"97",x"00"),
   693 => (x"c6",x"9c",x"c0",x"c3"),
   694 => (x"4b",x"73",x"2c",x"b7"),
   695 => (x"1e",x"73",x"b3",x"74"),
   696 => (x"72",x"1e",x"66",x"c4"),
   697 => (x"0b",x"60",x"27",x"1e"),
   698 => (x"27",x"1e",x"00",x"00"),
   699 => (x"00",x"00",x"01",x"51"),
   700 => (x"c2",x"86",x"d0",x"0f"),
   701 => (x"72",x"48",x"c1",x"82"),
   702 => (x"72",x"4a",x"70",x"30"),
   703 => (x"0b",x"8d",x"27",x"1e"),
   704 => (x"27",x"1e",x"00",x"00"),
   705 => (x"00",x"00",x"01",x"51"),
   706 => (x"c1",x"86",x"c8",x"0f"),
   707 => (x"c4",x"30",x"6e",x"48"),
   708 => (x"83",x"c1",x"58",x"a6"),
   709 => (x"95",x"72",x"4d",x"73"),
   710 => (x"1e",x"75",x"1e",x"6e"),
   711 => (x"00",x"0b",x"96",x"27"),
   712 => (x"51",x"27",x"1e",x"00"),
   713 => (x"0f",x"00",x"00",x"01"),
   714 => (x"49",x"6e",x"86",x"cc"),
   715 => (x"a9",x"b7",x"c0",x"c8"),
   716 => (x"87",x"cf",x"c0",x"06"),
   717 => (x"35",x"c1",x"4a",x"6e"),
   718 => (x"c8",x"2a",x"b7",x"c1"),
   719 => (x"01",x"aa",x"b7",x"c0"),
   720 => (x"75",x"87",x"f3",x"ff"),
   721 => (x"0b",x"ac",x"27",x"1e"),
   722 => (x"27",x"1e",x"00",x"00"),
   723 => (x"00",x"00",x"01",x"51"),
   724 => (x"75",x"86",x"c8",x"0f"),
   725 => (x"4d",x"26",x"26",x"48"),
   726 => (x"4b",x"26",x"4c",x"26"),
   727 => (x"4f",x"26",x"4a",x"26"),
   728 => (x"69",x"73",x"5f",x"63"),
   729 => (x"6d",x"5f",x"65",x"7a"),
   730 => (x"3a",x"74",x"6c",x"75"),
   731 => (x"2c",x"64",x"25",x"20"),
   732 => (x"61",x"65",x"72",x"20"),
   733 => (x"6c",x"62",x"5f",x"64"),
   734 => (x"6e",x"65",x"6c",x"5f"),
   735 => (x"64",x"25",x"20",x"3a"),
   736 => (x"73",x"63",x"20",x"2c"),
   737 => (x"3a",x"65",x"7a",x"69"),
   738 => (x"0a",x"64",x"25",x"20"),
   739 => (x"6c",x"75",x"4d",x"00"),
   740 => (x"64",x"25",x"20",x"74"),
   741 => (x"64",x"25",x"00",x"0a"),
   742 => (x"6f",x"6c",x"62",x"20"),
   743 => (x"20",x"73",x"6b",x"63"),
   744 => (x"73",x"20",x"66",x"6f"),
   745 => (x"20",x"65",x"7a",x"69"),
   746 => (x"00",x"0a",x"64",x"25"),
   747 => (x"62",x"20",x"64",x"25"),
   748 => (x"6b",x"63",x"6f",x"6c"),
   749 => (x"66",x"6f",x"20",x"73"),
   750 => (x"32",x"31",x"35",x"20"),
   751 => (x"74",x"79",x"62",x"20"),
   752 => (x"00",x"0a",x"73",x"65"),
   753 => (x"5b",x"5a",x"5e",x"0e"),
   754 => (x"d4",x"0e",x"5d",x"5c"),
   755 => (x"4c",x"c0",x"4d",x"66"),
   756 => (x"c0",x"49",x"66",x"dc"),
   757 => (x"c0",x"06",x"a9",x"b7"),
   758 => (x"4b",x"15",x"87",x"fb"),
   759 => (x"c0",x"c0",x"c0",x"c1"),
   760 => (x"c0",x"c4",x"93",x"c0"),
   761 => (x"d8",x"4b",x"93",x"b7"),
   762 => (x"4a",x"bf",x"97",x"66"),
   763 => (x"c0",x"c0",x"c0",x"c1"),
   764 => (x"c0",x"c4",x"92",x"c0"),
   765 => (x"d8",x"4a",x"92",x"b7"),
   766 => (x"80",x"c1",x"48",x"66"),
   767 => (x"72",x"58",x"a6",x"dc"),
   768 => (x"c0",x"02",x"ab",x"b7"),
   769 => (x"48",x"c1",x"87",x"c5"),
   770 => (x"c1",x"87",x"cc",x"c0"),
   771 => (x"b7",x"66",x"dc",x"84"),
   772 => (x"c5",x"ff",x"04",x"ac"),
   773 => (x"26",x"48",x"c0",x"87"),
   774 => (x"26",x"4c",x"26",x"4d"),
   775 => (x"26",x"4a",x"26",x"4b"),
   776 => (x"5a",x"5e",x"0e",x"4f"),
   777 => (x"0e",x"5d",x"5c",x"5b"),
   778 => (x"00",x"1d",x"d8",x"27"),
   779 => (x"79",x"c0",x"49",x"00"),
   780 => (x"00",x"1a",x"7b",x"27"),
   781 => (x"6e",x"27",x"1e",x"00"),
   782 => (x"0f",x"00",x"00",x"00"),
   783 => (x"d0",x"27",x"86",x"c4"),
   784 => (x"1e",x"00",x"00",x"1b"),
   785 => (x"57",x"27",x"1e",x"c0"),
   786 => (x"0f",x"00",x"00",x"09"),
   787 => (x"4a",x"70",x"86",x"c8"),
   788 => (x"c0",x"05",x"9a",x"72"),
   789 => (x"a7",x"27",x"87",x"d3"),
   790 => (x"1e",x"00",x"00",x"19"),
   791 => (x"00",x"00",x"6e",x"27"),
   792 => (x"86",x"c4",x"0f",x"00"),
   793 => (x"d8",x"cf",x"48",x"c0"),
   794 => (x"1a",x"88",x"27",x"87"),
   795 => (x"27",x"1e",x"00",x"00"),
   796 => (x"00",x"00",x"00",x"6e"),
   797 => (x"c0",x"86",x"c4",x"0f"),
   798 => (x"1e",x"04",x"27",x"4c"),
   799 => (x"c1",x"49",x"00",x"00"),
   800 => (x"27",x"1e",x"c8",x"79"),
   801 => (x"00",x"00",x"1a",x"9f"),
   802 => (x"1c",x"06",x"27",x"1e"),
   803 => (x"27",x"1e",x"00",x"00"),
   804 => (x"00",x"00",x"0b",x"c4"),
   805 => (x"70",x"86",x"cc",x"0f"),
   806 => (x"05",x"9a",x"72",x"4a"),
   807 => (x"27",x"87",x"c8",x"c0"),
   808 => (x"00",x"00",x"1e",x"04"),
   809 => (x"c8",x"79",x"c0",x"49"),
   810 => (x"1a",x"a8",x"27",x"1e"),
   811 => (x"27",x"1e",x"00",x"00"),
   812 => (x"00",x"00",x"1c",x"22"),
   813 => (x"0b",x"c4",x"27",x"1e"),
   814 => (x"cc",x"0f",x"00",x"00"),
   815 => (x"72",x"4a",x"70",x"86"),
   816 => (x"c8",x"c0",x"05",x"9a"),
   817 => (x"1e",x"04",x"27",x"87"),
   818 => (x"c0",x"49",x"00",x"00"),
   819 => (x"1e",x"04",x"27",x"79"),
   820 => (x"1e",x"bf",x"00",x"00"),
   821 => (x"00",x"1a",x"b1",x"27"),
   822 => (x"51",x"27",x"1e",x"00"),
   823 => (x"0f",x"00",x"00",x"01"),
   824 => (x"04",x"27",x"86",x"c8"),
   825 => (x"bf",x"00",x"00",x"1e"),
   826 => (x"87",x"c0",x"c3",x"02"),
   827 => (x"00",x"1b",x"d0",x"27"),
   828 => (x"8e",x"27",x"4d",x"00"),
   829 => (x"4b",x"00",x"00",x"1d"),
   830 => (x"00",x"1d",x"ce",x"27"),
   831 => (x"4a",x"bf",x"9f",x"00"),
   832 => (x"ce",x"27",x"1e",x"72"),
   833 => (x"4a",x"00",x"00",x"1d"),
   834 => (x"00",x"1b",x"d0",x"27"),
   835 => (x"1e",x"72",x"8a",x"00"),
   836 => (x"c0",x"c8",x"1e",x"d0"),
   837 => (x"19",x"d9",x"27",x"1e"),
   838 => (x"27",x"1e",x"00",x"00"),
   839 => (x"00",x"00",x"01",x"51"),
   840 => (x"73",x"86",x"d4",x"0f"),
   841 => (x"6a",x"82",x"c8",x"4a"),
   842 => (x"1d",x"ce",x"27",x"4c"),
   843 => (x"bf",x"9f",x"00",x"00"),
   844 => (x"ea",x"d6",x"c5",x"4a"),
   845 => (x"c0",x"05",x"aa",x"b7"),
   846 => (x"4a",x"73",x"87",x"d3"),
   847 => (x"1e",x"6a",x"82",x"c8"),
   848 => (x"00",x"13",x"a2",x"27"),
   849 => (x"86",x"c4",x"0f",x"00"),
   850 => (x"e4",x"c0",x"4c",x"70"),
   851 => (x"c7",x"4a",x"75",x"87"),
   852 => (x"6a",x"9f",x"82",x"fe"),
   853 => (x"d5",x"e9",x"ca",x"4a"),
   854 => (x"c0",x"02",x"aa",x"b7"),
   855 => (x"bb",x"27",x"87",x"d3"),
   856 => (x"1e",x"00",x"00",x"19"),
   857 => (x"00",x"00",x"6e",x"27"),
   858 => (x"86",x"c4",x"0f",x"00"),
   859 => (x"d0",x"cb",x"48",x"c0"),
   860 => (x"27",x"1e",x"74",x"87"),
   861 => (x"00",x"00",x"1a",x"16"),
   862 => (x"01",x"51",x"27",x"1e"),
   863 => (x"c8",x"0f",x"00",x"00"),
   864 => (x"1b",x"d0",x"27",x"86"),
   865 => (x"74",x"1e",x"00",x"00"),
   866 => (x"09",x"57",x"27",x"1e"),
   867 => (x"c8",x"0f",x"00",x"00"),
   868 => (x"72",x"4a",x"70",x"86"),
   869 => (x"c5",x"c0",x"05",x"9a"),
   870 => (x"ca",x"48",x"c0",x"87"),
   871 => (x"2e",x"27",x"87",x"e3"),
   872 => (x"1e",x"00",x"00",x"1a"),
   873 => (x"00",x"00",x"6e",x"27"),
   874 => (x"86",x"c4",x"0f",x"00"),
   875 => (x"00",x"1a",x"c4",x"27"),
   876 => (x"51",x"27",x"1e",x"00"),
   877 => (x"0f",x"00",x"00",x"01"),
   878 => (x"1e",x"c8",x"86",x"c4"),
   879 => (x"00",x"1a",x"dc",x"27"),
   880 => (x"22",x"27",x"1e",x"00"),
   881 => (x"1e",x"00",x"00",x"1c"),
   882 => (x"00",x"0b",x"c4",x"27"),
   883 => (x"86",x"cc",x"0f",x"00"),
   884 => (x"9a",x"72",x"4a",x"70"),
   885 => (x"87",x"cb",x"c0",x"05"),
   886 => (x"00",x"1d",x"d8",x"27"),
   887 => (x"79",x"c1",x"49",x"00"),
   888 => (x"c8",x"87",x"f1",x"c0"),
   889 => (x"1a",x"e5",x"27",x"1e"),
   890 => (x"27",x"1e",x"00",x"00"),
   891 => (x"00",x"00",x"1c",x"06"),
   892 => (x"0b",x"c4",x"27",x"1e"),
   893 => (x"cc",x"0f",x"00",x"00"),
   894 => (x"72",x"4a",x"70",x"86"),
   895 => (x"d3",x"c0",x"02",x"9a"),
   896 => (x"1a",x"55",x"27",x"87"),
   897 => (x"27",x"1e",x"00",x"00"),
   898 => (x"00",x"00",x"01",x"51"),
   899 => (x"c0",x"86",x"c4",x"0f"),
   900 => (x"87",x"ed",x"c8",x"48"),
   901 => (x"00",x"1d",x"ce",x"27"),
   902 => (x"4a",x"bf",x"97",x"00"),
   903 => (x"aa",x"b7",x"d5",x"c1"),
   904 => (x"87",x"d0",x"c0",x"05"),
   905 => (x"00",x"1d",x"cf",x"27"),
   906 => (x"4a",x"bf",x"97",x"00"),
   907 => (x"aa",x"b7",x"ea",x"c2"),
   908 => (x"87",x"c5",x"c0",x"02"),
   909 => (x"c8",x"c8",x"48",x"c0"),
   910 => (x"1b",x"d0",x"27",x"87"),
   911 => (x"bf",x"97",x"00",x"00"),
   912 => (x"b7",x"e9",x"c3",x"4a"),
   913 => (x"d5",x"c0",x"02",x"aa"),
   914 => (x"1b",x"d0",x"27",x"87"),
   915 => (x"bf",x"97",x"00",x"00"),
   916 => (x"b7",x"eb",x"c3",x"4a"),
   917 => (x"c5",x"c0",x"02",x"aa"),
   918 => (x"c7",x"48",x"c0",x"87"),
   919 => (x"db",x"27",x"87",x"e3"),
   920 => (x"97",x"00",x"00",x"1b"),
   921 => (x"9a",x"72",x"4a",x"bf"),
   922 => (x"87",x"cf",x"c0",x"05"),
   923 => (x"00",x"1b",x"dc",x"27"),
   924 => (x"4a",x"bf",x"97",x"00"),
   925 => (x"02",x"aa",x"b7",x"c2"),
   926 => (x"c0",x"87",x"c5",x"c0"),
   927 => (x"87",x"c1",x"c7",x"48"),
   928 => (x"00",x"1b",x"dd",x"27"),
   929 => (x"48",x"bf",x"97",x"00"),
   930 => (x"00",x"1d",x"d4",x"27"),
   931 => (x"d0",x"27",x"58",x"00"),
   932 => (x"bf",x"00",x"00",x"1d"),
   933 => (x"c1",x"4b",x"72",x"4a"),
   934 => (x"1d",x"d4",x"27",x"8b"),
   935 => (x"73",x"49",x"00",x"00"),
   936 => (x"72",x"1e",x"73",x"79"),
   937 => (x"1a",x"ee",x"27",x"1e"),
   938 => (x"27",x"1e",x"00",x"00"),
   939 => (x"00",x"00",x"01",x"51"),
   940 => (x"27",x"86",x"cc",x"0f"),
   941 => (x"00",x"00",x"1b",x"de"),
   942 => (x"74",x"4a",x"bf",x"97"),
   943 => (x"1b",x"df",x"27",x"82"),
   944 => (x"bf",x"97",x"00",x"00"),
   945 => (x"73",x"33",x"c8",x"4b"),
   946 => (x"27",x"80",x"72",x"48"),
   947 => (x"00",x"00",x"1d",x"e8"),
   948 => (x"1b",x"e0",x"27",x"58"),
   949 => (x"bf",x"97",x"00",x"00"),
   950 => (x"1d",x"fc",x"27",x"48"),
   951 => (x"27",x"58",x"00",x"00"),
   952 => (x"00",x"00",x"1d",x"d8"),
   953 => (x"df",x"c3",x"02",x"bf"),
   954 => (x"27",x"1e",x"c8",x"87"),
   955 => (x"00",x"00",x"1a",x"72"),
   956 => (x"1c",x"22",x"27",x"1e"),
   957 => (x"27",x"1e",x"00",x"00"),
   958 => (x"00",x"00",x"0b",x"c4"),
   959 => (x"70",x"86",x"cc",x"0f"),
   960 => (x"02",x"9a",x"72",x"4a"),
   961 => (x"c0",x"87",x"c5",x"c0"),
   962 => (x"87",x"f5",x"c4",x"48"),
   963 => (x"00",x"1d",x"d0",x"27"),
   964 => (x"73",x"4b",x"bf",x"00"),
   965 => (x"27",x"30",x"c4",x"48"),
   966 => (x"00",x"00",x"1e",x"00"),
   967 => (x"1d",x"f4",x"27",x"58"),
   968 => (x"73",x"49",x"00",x"00"),
   969 => (x"1b",x"f5",x"27",x"79"),
   970 => (x"bf",x"97",x"00",x"00"),
   971 => (x"27",x"32",x"c8",x"4a"),
   972 => (x"00",x"00",x"1b",x"f4"),
   973 => (x"72",x"4c",x"bf",x"97"),
   974 => (x"27",x"82",x"74",x"4a"),
   975 => (x"00",x"00",x"1b",x"f6"),
   976 => (x"d0",x"4c",x"bf",x"97"),
   977 => (x"74",x"4a",x"72",x"34"),
   978 => (x"1b",x"f7",x"27",x"82"),
   979 => (x"bf",x"97",x"00",x"00"),
   980 => (x"72",x"34",x"d8",x"4c"),
   981 => (x"27",x"82",x"74",x"4a"),
   982 => (x"00",x"00",x"1e",x"00"),
   983 => (x"72",x"79",x"72",x"49"),
   984 => (x"1d",x"f8",x"27",x"4a"),
   985 => (x"92",x"bf",x"00",x"00"),
   986 => (x"e4",x"27",x"4a",x"72"),
   987 => (x"bf",x"00",x"00",x"1d"),
   988 => (x"1d",x"e8",x"27",x"82"),
   989 => (x"72",x"49",x"00",x"00"),
   990 => (x"1b",x"fd",x"27",x"79"),
   991 => (x"bf",x"97",x"00",x"00"),
   992 => (x"27",x"34",x"c8",x"4c"),
   993 => (x"00",x"00",x"1b",x"fc"),
   994 => (x"74",x"4d",x"bf",x"97"),
   995 => (x"27",x"84",x"75",x"4c"),
   996 => (x"00",x"00",x"1b",x"fe"),
   997 => (x"d0",x"4d",x"bf",x"97"),
   998 => (x"75",x"4c",x"74",x"35"),
   999 => (x"1b",x"ff",x"27",x"84"),
  1000 => (x"bf",x"97",x"00",x"00"),
  1001 => (x"d8",x"9d",x"cf",x"4d"),
  1002 => (x"75",x"4c",x"74",x"35"),
  1003 => (x"1d",x"ec",x"27",x"84"),
  1004 => (x"74",x"49",x"00",x"00"),
  1005 => (x"73",x"8c",x"c2",x"79"),
  1006 => (x"73",x"93",x"74",x"4b"),
  1007 => (x"27",x"80",x"72",x"48"),
  1008 => (x"00",x"00",x"1d",x"f4"),
  1009 => (x"87",x"f7",x"c1",x"58"),
  1010 => (x"00",x"1b",x"e2",x"27"),
  1011 => (x"4a",x"bf",x"97",x"00"),
  1012 => (x"e1",x"27",x"32",x"c8"),
  1013 => (x"97",x"00",x"00",x"1b"),
  1014 => (x"4a",x"72",x"4b",x"bf"),
  1015 => (x"fc",x"27",x"82",x"73"),
  1016 => (x"49",x"00",x"00",x"1d"),
  1017 => (x"32",x"c5",x"79",x"72"),
  1018 => (x"c9",x"82",x"ff",x"c7"),
  1019 => (x"1d",x"f4",x"27",x"2a"),
  1020 => (x"72",x"49",x"00",x"00"),
  1021 => (x"1b",x"e7",x"27",x"79"),
  1022 => (x"bf",x"97",x"00",x"00"),
  1023 => (x"27",x"33",x"c8",x"4b"),
  1024 => (x"00",x"00",x"1b",x"e6"),
  1025 => (x"73",x"4c",x"bf",x"97"),
  1026 => (x"27",x"83",x"74",x"4b"),
  1027 => (x"00",x"00",x"1e",x"00"),
  1028 => (x"73",x"79",x"73",x"49"),
  1029 => (x"1d",x"f8",x"27",x"4b"),
  1030 => (x"93",x"bf",x"00",x"00"),
  1031 => (x"e4",x"27",x"4b",x"73"),
  1032 => (x"bf",x"00",x"00",x"1d"),
  1033 => (x"1d",x"f0",x"27",x"83"),
  1034 => (x"73",x"49",x"00",x"00"),
  1035 => (x"1d",x"ec",x"27",x"79"),
  1036 => (x"c0",x"49",x"00",x"00"),
  1037 => (x"72",x"48",x"73",x"79"),
  1038 => (x"1d",x"ec",x"27",x"80"),
  1039 => (x"c1",x"58",x"00",x"00"),
  1040 => (x"26",x"4d",x"26",x"48"),
  1041 => (x"26",x"4b",x"26",x"4c"),
  1042 => (x"0e",x"4f",x"26",x"4a"),
  1043 => (x"5c",x"5b",x"5a",x"5e"),
  1044 => (x"d8",x"27",x"0e",x"5d"),
  1045 => (x"bf",x"00",x"00",x"1d"),
  1046 => (x"87",x"cf",x"c0",x"02"),
  1047 => (x"c7",x"4c",x"66",x"d4"),
  1048 => (x"66",x"d4",x"2c",x"b7"),
  1049 => (x"9b",x"ff",x"c1",x"4b"),
  1050 => (x"d4",x"87",x"cc",x"c0"),
  1051 => (x"b7",x"c8",x"4c",x"66"),
  1052 => (x"4b",x"66",x"d4",x"2c"),
  1053 => (x"27",x"9b",x"ff",x"c3"),
  1054 => (x"00",x"00",x"1b",x"d0"),
  1055 => (x"1d",x"e4",x"27",x"1e"),
  1056 => (x"4a",x"bf",x"00",x"00"),
  1057 => (x"1e",x"72",x"82",x"74"),
  1058 => (x"00",x"09",x"57",x"27"),
  1059 => (x"86",x"c8",x"0f",x"00"),
  1060 => (x"9a",x"72",x"4a",x"70"),
  1061 => (x"87",x"c5",x"c0",x"05"),
  1062 => (x"f2",x"c0",x"48",x"c0"),
  1063 => (x"1d",x"d8",x"27",x"87"),
  1064 => (x"02",x"bf",x"00",x"00"),
  1065 => (x"73",x"87",x"d7",x"c0"),
  1066 => (x"72",x"92",x"c4",x"4a"),
  1067 => (x"1b",x"d0",x"27",x"4a"),
  1068 => (x"6a",x"82",x"00",x"00"),
  1069 => (x"ff",x"ff",x"cf",x"4d"),
  1070 => (x"c0",x"9d",x"ff",x"ff"),
  1071 => (x"4a",x"73",x"87",x"cf"),
  1072 => (x"4a",x"72",x"92",x"c2"),
  1073 => (x"00",x"1b",x"d0",x"27"),
  1074 => (x"6a",x"9f",x"82",x"00"),
  1075 => (x"26",x"48",x"75",x"4d"),
  1076 => (x"26",x"4c",x"26",x"4d"),
  1077 => (x"26",x"4a",x"26",x"4b"),
  1078 => (x"5a",x"5e",x"0e",x"4f"),
  1079 => (x"0e",x"5d",x"5c",x"5b"),
  1080 => (x"ff",x"cf",x"8e",x"cc"),
  1081 => (x"4d",x"f8",x"ff",x"ff"),
  1082 => (x"49",x"76",x"4c",x"c0"),
  1083 => (x"00",x"1d",x"ec",x"27"),
  1084 => (x"c4",x"79",x"bf",x"00"),
  1085 => (x"f0",x"27",x"49",x"a6"),
  1086 => (x"bf",x"00",x"00",x"1d"),
  1087 => (x"1d",x"d8",x"27",x"79"),
  1088 => (x"02",x"bf",x"00",x"00"),
  1089 => (x"27",x"87",x"cc",x"c0"),
  1090 => (x"00",x"00",x"1d",x"d0"),
  1091 => (x"32",x"c4",x"4a",x"bf"),
  1092 => (x"27",x"87",x"c9",x"c0"),
  1093 => (x"00",x"00",x"1d",x"f4"),
  1094 => (x"32",x"c4",x"4a",x"bf"),
  1095 => (x"72",x"49",x"a6",x"c8"),
  1096 => (x"c8",x"4b",x"c0",x"79"),
  1097 => (x"a9",x"c0",x"49",x"66"),
  1098 => (x"87",x"c6",x"c3",x"06"),
  1099 => (x"9a",x"cf",x"4a",x"73"),
  1100 => (x"c0",x"05",x"9a",x"72"),
  1101 => (x"d0",x"27",x"87",x"e4"),
  1102 => (x"1e",x"00",x"00",x"1b"),
  1103 => (x"c8",x"4a",x"66",x"c8"),
  1104 => (x"80",x"c1",x"48",x"66"),
  1105 => (x"72",x"58",x"a6",x"cc"),
  1106 => (x"09",x"57",x"27",x"1e"),
  1107 => (x"c8",x"0f",x"00",x"00"),
  1108 => (x"1b",x"d0",x"27",x"86"),
  1109 => (x"c0",x"4c",x"00",x"00"),
  1110 => (x"e0",x"c0",x"87",x"c3"),
  1111 => (x"4a",x"6c",x"97",x"84"),
  1112 => (x"c2",x"02",x"9a",x"72"),
  1113 => (x"6c",x"97",x"87",x"c3"),
  1114 => (x"b7",x"e5",x"c3",x"4a"),
  1115 => (x"f8",x"c1",x"02",x"aa"),
  1116 => (x"cb",x"4a",x"74",x"87"),
  1117 => (x"4a",x"6a",x"97",x"82"),
  1118 => (x"9a",x"72",x"9a",x"d8"),
  1119 => (x"87",x"e9",x"c1",x"05"),
  1120 => (x"e8",x"c0",x"1e",x"cb"),
  1121 => (x"1e",x"74",x"1e",x"66"),
  1122 => (x"00",x"0b",x"c4",x"27"),
  1123 => (x"86",x"cc",x"0f",x"00"),
  1124 => (x"9a",x"72",x"4a",x"70"),
  1125 => (x"87",x"d1",x"c1",x"05"),
  1126 => (x"83",x"dc",x"4b",x"74"),
  1127 => (x"4a",x"66",x"e0",x"c0"),
  1128 => (x"7a",x"6b",x"82",x"c4"),
  1129 => (x"83",x"da",x"4b",x"74"),
  1130 => (x"4a",x"66",x"e0",x"c0"),
  1131 => (x"6b",x"9f",x"82",x"c8"),
  1132 => (x"72",x"7a",x"70",x"48"),
  1133 => (x"1d",x"d8",x"27",x"4d"),
  1134 => (x"02",x"bf",x"00",x"00"),
  1135 => (x"74",x"87",x"d5",x"c0"),
  1136 => (x"9f",x"82",x"d4",x"4a"),
  1137 => (x"ff",x"c0",x"4a",x"6a"),
  1138 => (x"48",x"72",x"9a",x"ff"),
  1139 => (x"a6",x"c4",x"30",x"d0"),
  1140 => (x"87",x"c4",x"c0",x"58"),
  1141 => (x"79",x"c0",x"49",x"76"),
  1142 => (x"80",x"6d",x"48",x"6e"),
  1143 => (x"e0",x"c0",x"7d",x"70"),
  1144 => (x"79",x"c0",x"49",x"66"),
  1145 => (x"ce",x"c1",x"48",x"c1"),
  1146 => (x"c8",x"83",x"c1",x"87"),
  1147 => (x"fc",x"04",x"ab",x"66"),
  1148 => (x"ff",x"cf",x"87",x"fa"),
  1149 => (x"4d",x"f8",x"ff",x"ff"),
  1150 => (x"00",x"1d",x"d8",x"27"),
  1151 => (x"c0",x"02",x"bf",x"00"),
  1152 => (x"1e",x"6e",x"87",x"f3"),
  1153 => (x"00",x"10",x"4b",x"27"),
  1154 => (x"86",x"c4",x"0f",x"00"),
  1155 => (x"6e",x"58",x"a6",x"c4"),
  1156 => (x"75",x"9a",x"75",x"4a"),
  1157 => (x"dc",x"c0",x"02",x"aa"),
  1158 => (x"c2",x"4a",x"6e",x"87"),
  1159 => (x"27",x"4a",x"72",x"8a"),
  1160 => (x"00",x"00",x"1d",x"d0"),
  1161 => (x"e8",x"27",x"92",x"bf"),
  1162 => (x"bf",x"00",x"00",x"1d"),
  1163 => (x"c8",x"80",x"72",x"48"),
  1164 => (x"ec",x"fb",x"58",x"a6"),
  1165 => (x"cf",x"48",x"c0",x"87"),
  1166 => (x"f8",x"ff",x"ff",x"ff"),
  1167 => (x"26",x"86",x"cc",x"4d"),
  1168 => (x"26",x"4c",x"26",x"4d"),
  1169 => (x"26",x"4a",x"26",x"4b"),
  1170 => (x"5a",x"5e",x"0e",x"4f"),
  1171 => (x"66",x"cc",x"0e",x"5b"),
  1172 => (x"82",x"c1",x"4a",x"bf"),
  1173 => (x"72",x"49",x"66",x"cc"),
  1174 => (x"27",x"4a",x"72",x"79"),
  1175 => (x"00",x"00",x"1d",x"d4"),
  1176 => (x"9a",x"72",x"9a",x"bf"),
  1177 => (x"87",x"d3",x"c0",x"05"),
  1178 => (x"c8",x"4a",x"66",x"cc"),
  1179 => (x"27",x"1e",x"6a",x"82"),
  1180 => (x"00",x"00",x"10",x"4b"),
  1181 => (x"70",x"86",x"c4",x"0f"),
  1182 => (x"c1",x"7a",x"73",x"4b"),
  1183 => (x"26",x"4b",x"26",x"48"),
  1184 => (x"0e",x"4f",x"26",x"4a"),
  1185 => (x"0e",x"5b",x"5a",x"5e"),
  1186 => (x"00",x"1d",x"e8",x"27"),
  1187 => (x"cc",x"4a",x"bf",x"00"),
  1188 => (x"83",x"c8",x"4b",x"66"),
  1189 => (x"8b",x"c2",x"4b",x"6b"),
  1190 => (x"d0",x"27",x"4b",x"73"),
  1191 => (x"bf",x"00",x"00",x"1d"),
  1192 => (x"73",x"4a",x"72",x"93"),
  1193 => (x"1d",x"d4",x"27",x"82"),
  1194 => (x"4b",x"bf",x"00",x"00"),
  1195 => (x"9b",x"bf",x"66",x"cc"),
  1196 => (x"82",x"73",x"4a",x"72"),
  1197 => (x"72",x"1e",x"66",x"d0"),
  1198 => (x"09",x"57",x"27",x"1e"),
  1199 => (x"c8",x"0f",x"00",x"00"),
  1200 => (x"72",x"4a",x"70",x"86"),
  1201 => (x"c5",x"c0",x"05",x"9a"),
  1202 => (x"c0",x"48",x"c0",x"87"),
  1203 => (x"48",x"c1",x"87",x"c2"),
  1204 => (x"4a",x"26",x"4b",x"26"),
  1205 => (x"5e",x"0e",x"4f",x"26"),
  1206 => (x"5d",x"5c",x"5b",x"5a"),
  1207 => (x"4c",x"66",x"d8",x"0e"),
  1208 => (x"27",x"1e",x"66",x"d4"),
  1209 => (x"00",x"00",x"1e",x"08"),
  1210 => (x"10",x"d9",x"27",x"1e"),
  1211 => (x"c8",x"0f",x"00",x"00"),
  1212 => (x"72",x"4a",x"70",x"86"),
  1213 => (x"df",x"c1",x"02",x"9a"),
  1214 => (x"1e",x"0c",x"27",x"87"),
  1215 => (x"4a",x"bf",x"00",x"00"),
  1216 => (x"c9",x"82",x"ff",x"c7"),
  1217 => (x"c0",x"4d",x"72",x"2a"),
  1218 => (x"13",x"7a",x"27",x"4b"),
  1219 => (x"27",x"1e",x"00",x"00"),
  1220 => (x"00",x"00",x"00",x"6e"),
  1221 => (x"c0",x"86",x"c4",x"0f"),
  1222 => (x"c1",x"06",x"ad",x"b7"),
  1223 => (x"1e",x"74",x"87",x"d0"),
  1224 => (x"00",x"1e",x"08",x"27"),
  1225 => (x"83",x"27",x"1e",x"00"),
  1226 => (x"0f",x"00",x"00",x"12"),
  1227 => (x"4a",x"70",x"86",x"c8"),
  1228 => (x"c0",x"05",x"9a",x"72"),
  1229 => (x"48",x"c0",x"87",x"c5"),
  1230 => (x"27",x"87",x"f5",x"c0"),
  1231 => (x"00",x"00",x"1e",x"08"),
  1232 => (x"12",x"49",x"27",x"1e"),
  1233 => (x"c4",x"0f",x"00",x"00"),
  1234 => (x"84",x"c0",x"c8",x"86"),
  1235 => (x"b7",x"75",x"83",x"c1"),
  1236 => (x"c9",x"ff",x"04",x"ab"),
  1237 => (x"87",x"d6",x"c0",x"87"),
  1238 => (x"27",x"1e",x"66",x"d4"),
  1239 => (x"00",x"00",x"13",x"93"),
  1240 => (x"01",x"51",x"27",x"1e"),
  1241 => (x"c8",x"0f",x"00",x"00"),
  1242 => (x"c0",x"48",x"c0",x"86"),
  1243 => (x"48",x"c1",x"87",x"c2"),
  1244 => (x"4c",x"26",x"4d",x"26"),
  1245 => (x"4a",x"26",x"4b",x"26"),
  1246 => (x"70",x"4f",x"4f",x"26"),
  1247 => (x"64",x"65",x"6e",x"65"),
  1248 => (x"6c",x"69",x"66",x"20"),
  1249 => (x"6c",x"20",x"2c",x"65"),
  1250 => (x"69",x"64",x"61",x"6f"),
  1251 => (x"2e",x"2e",x"67",x"6e"),
  1252 => (x"43",x"00",x"0a",x"2e"),
  1253 => (x"74",x"27",x"6e",x"61"),
  1254 => (x"65",x"70",x"6f",x"20"),
  1255 => (x"73",x"25",x"20",x"6e"),
  1256 => (x"5e",x"0e",x"00",x"0a"),
  1257 => (x"cc",x"0e",x"5b",x"5a"),
  1258 => (x"2a",x"d8",x"4a",x"66"),
  1259 => (x"cc",x"9a",x"ff",x"c3"),
  1260 => (x"2b",x"c8",x"4b",x"66"),
  1261 => (x"9b",x"c0",x"fc",x"cf"),
  1262 => (x"b2",x"73",x"4a",x"72"),
  1263 => (x"c8",x"4b",x"66",x"cc"),
  1264 => (x"f0",x"ff",x"c0",x"33"),
  1265 => (x"72",x"9b",x"c0",x"c0"),
  1266 => (x"cc",x"b2",x"73",x"4a"),
  1267 => (x"33",x"d8",x"4b",x"66"),
  1268 => (x"c0",x"c0",x"c0",x"ff"),
  1269 => (x"4a",x"72",x"9b",x"c0"),
  1270 => (x"48",x"72",x"b2",x"73"),
  1271 => (x"4a",x"26",x"4b",x"26"),
  1272 => (x"5e",x"0e",x"4f",x"26"),
  1273 => (x"cc",x"0e",x"5b",x"5a"),
  1274 => (x"2b",x"c8",x"4b",x"66"),
  1275 => (x"4b",x"9b",x"ff",x"c3"),
  1276 => (x"c8",x"4a",x"66",x"cc"),
  1277 => (x"c0",x"fc",x"cf",x"32"),
  1278 => (x"73",x"4a",x"72",x"9a"),
  1279 => (x"48",x"72",x"4a",x"b2"),
  1280 => (x"4a",x"26",x"4b",x"26"),
  1281 => (x"5e",x"0e",x"4f",x"26"),
  1282 => (x"cc",x"0e",x"5b",x"5a"),
  1283 => (x"2a",x"d0",x"4a",x"66"),
  1284 => (x"9a",x"ff",x"ff",x"cf"),
  1285 => (x"4b",x"66",x"cc",x"4a"),
  1286 => (x"c0",x"f0",x"33",x"d0"),
  1287 => (x"4a",x"72",x"9b",x"c0"),
  1288 => (x"48",x"72",x"b2",x"73"),
  1289 => (x"4a",x"26",x"4b",x"26"),
  1290 => (x"ff",x"1e",x"4f",x"26"),
  1291 => (x"4f",x"26",x"87",x"fd"),
  1292 => (x"cc",x"1e",x"72",x"1e"),
  1293 => (x"df",x"c3",x"4a",x"66"),
  1294 => (x"8a",x"f7",x"c0",x"9a"),
  1295 => (x"03",x"aa",x"b7",x"c0"),
  1296 => (x"c0",x"87",x"c3",x"c0"),
  1297 => (x"66",x"c8",x"82",x"e7"),
  1298 => (x"cc",x"30",x"c4",x"48"),
  1299 => (x"66",x"c8",x"58",x"a6"),
  1300 => (x"cc",x"b0",x"72",x"48"),
  1301 => (x"66",x"c8",x"58",x"a6"),
  1302 => (x"26",x"4a",x"26",x"48"),
  1303 => (x"5a",x"5e",x"0e",x"4f"),
  1304 => (x"27",x"0e",x"5c",x"5b"),
  1305 => (x"00",x"00",x"1e",x"18"),
  1306 => (x"80",x"c1",x"48",x"bf"),
  1307 => (x"00",x"1e",x"1c",x"27"),
  1308 => (x"d0",x"97",x"58",x"00"),
  1309 => (x"c0",x"c1",x"4a",x"66"),
  1310 => (x"92",x"c0",x"c0",x"c0"),
  1311 => (x"92",x"b7",x"c0",x"c4"),
  1312 => (x"b7",x"d3",x"c1",x"4a"),
  1313 => (x"e9",x"c0",x"05",x"aa"),
  1314 => (x"1e",x"18",x"27",x"87"),
  1315 => (x"c0",x"49",x"00",x"00"),
  1316 => (x"1e",x"1c",x"27",x"79"),
  1317 => (x"c0",x"49",x"00",x"00"),
  1318 => (x"1e",x"24",x"27",x"79"),
  1319 => (x"c0",x"49",x"00",x"00"),
  1320 => (x"1e",x"28",x"27",x"79"),
  1321 => (x"c0",x"49",x"00",x"00"),
  1322 => (x"49",x"c0",x"ff",x"79"),
  1323 => (x"c9",x"79",x"d3",x"c1"),
  1324 => (x"18",x"27",x"87",x"f6"),
  1325 => (x"bf",x"00",x"00",x"1e"),
  1326 => (x"a9",x"b7",x"c1",x"49"),
  1327 => (x"87",x"db",x"c1",x"05"),
  1328 => (x"c1",x"49",x"c0",x"ff"),
  1329 => (x"d0",x"97",x"79",x"f4"),
  1330 => (x"c0",x"c1",x"4a",x"66"),
  1331 => (x"92",x"c0",x"c0",x"c0"),
  1332 => (x"92",x"b7",x"c0",x"c4"),
  1333 => (x"27",x"1e",x"72",x"4a"),
  1334 => (x"00",x"00",x"1e",x"28"),
  1335 => (x"30",x"27",x"1e",x"bf"),
  1336 => (x"0f",x"00",x"00",x"14"),
  1337 => (x"2c",x"27",x"86",x"c8"),
  1338 => (x"58",x"00",x"00",x"1e"),
  1339 => (x"00",x"1e",x"28",x"27"),
  1340 => (x"c3",x"4c",x"bf",x"00"),
  1341 => (x"c0",x"06",x"ac",x"b7"),
  1342 => (x"48",x"ca",x"87",x"c6"),
  1343 => (x"4c",x"70",x"88",x"74"),
  1344 => (x"82",x"c1",x"4a",x"74"),
  1345 => (x"30",x"c1",x"48",x"72"),
  1346 => (x"00",x"1e",x"24",x"27"),
  1347 => (x"48",x"74",x"58",x"00"),
  1348 => (x"ff",x"80",x"f0",x"c0"),
  1349 => (x"79",x"70",x"49",x"c0"),
  1350 => (x"27",x"87",x"cd",x"c8"),
  1351 => (x"00",x"00",x"1e",x"28"),
  1352 => (x"b7",x"c9",x"49",x"bf"),
  1353 => (x"ff",x"c7",x"01",x"a9"),
  1354 => (x"1e",x"28",x"27",x"87"),
  1355 => (x"49",x"bf",x"00",x"00"),
  1356 => (x"06",x"a9",x"b7",x"c0"),
  1357 => (x"27",x"87",x"f1",x"c7"),
  1358 => (x"00",x"00",x"1e",x"28"),
  1359 => (x"f0",x"c0",x"48",x"bf"),
  1360 => (x"49",x"c0",x"ff",x"80"),
  1361 => (x"18",x"27",x"79",x"70"),
  1362 => (x"bf",x"00",x"00",x"1e"),
  1363 => (x"a9",x"b7",x"c3",x"49"),
  1364 => (x"87",x"e9",x"c0",x"01"),
  1365 => (x"4a",x"66",x"d0",x"97"),
  1366 => (x"c0",x"c0",x"c0",x"c1"),
  1367 => (x"c0",x"c4",x"92",x"c0"),
  1368 => (x"72",x"4a",x"92",x"b7"),
  1369 => (x"1e",x"24",x"27",x"1e"),
  1370 => (x"1e",x"bf",x"00",x"00"),
  1371 => (x"00",x"14",x"30",x"27"),
  1372 => (x"86",x"c8",x"0f",x"00"),
  1373 => (x"00",x"1e",x"28",x"27"),
  1374 => (x"eb",x"c6",x"58",x"00"),
  1375 => (x"1e",x"20",x"27",x"87"),
  1376 => (x"4a",x"bf",x"00",x"00"),
  1377 => (x"18",x"27",x"82",x"c3"),
  1378 => (x"bf",x"00",x"00",x"1e"),
  1379 => (x"a9",x"b7",x"72",x"49"),
  1380 => (x"87",x"f1",x"c0",x"01"),
  1381 => (x"4a",x"66",x"d0",x"97"),
  1382 => (x"c0",x"c0",x"c0",x"c1"),
  1383 => (x"c0",x"c4",x"92",x"c0"),
  1384 => (x"72",x"4a",x"92",x"b7"),
  1385 => (x"1e",x"1c",x"27",x"1e"),
  1386 => (x"1e",x"bf",x"00",x"00"),
  1387 => (x"00",x"14",x"30",x"27"),
  1388 => (x"86",x"c8",x"0f",x"00"),
  1389 => (x"00",x"1e",x"20",x"27"),
  1390 => (x"2c",x"27",x"58",x"00"),
  1391 => (x"49",x"00",x"00",x"1e"),
  1392 => (x"e3",x"c5",x"79",x"c1"),
  1393 => (x"1e",x"28",x"27",x"87"),
  1394 => (x"49",x"bf",x"00",x"00"),
  1395 => (x"06",x"a9",x"b7",x"c0"),
  1396 => (x"27",x"87",x"d0",x"c3"),
  1397 => (x"00",x"00",x"1e",x"28"),
  1398 => (x"b7",x"c3",x"49",x"bf"),
  1399 => (x"c2",x"c3",x"01",x"a9"),
  1400 => (x"1e",x"24",x"27",x"87"),
  1401 => (x"4a",x"bf",x"00",x"00"),
  1402 => (x"82",x"c1",x"32",x"c1"),
  1403 => (x"00",x"1e",x"18",x"27"),
  1404 => (x"72",x"49",x"bf",x"00"),
  1405 => (x"c2",x"01",x"a9",x"b7"),
  1406 => (x"d0",x"97",x"87",x"c2"),
  1407 => (x"c0",x"c1",x"4a",x"66"),
  1408 => (x"92",x"c0",x"c0",x"c0"),
  1409 => (x"92",x"b7",x"c0",x"c4"),
  1410 => (x"27",x"1e",x"72",x"4a"),
  1411 => (x"00",x"00",x"1e",x"30"),
  1412 => (x"30",x"27",x"1e",x"bf"),
  1413 => (x"0f",x"00",x"00",x"14"),
  1414 => (x"34",x"27",x"86",x"c8"),
  1415 => (x"58",x"00",x"00",x"1e"),
  1416 => (x"00",x"1e",x"2c",x"27"),
  1417 => (x"c1",x"4a",x"bf",x"00"),
  1418 => (x"1e",x"2c",x"27",x"8a"),
  1419 => (x"72",x"49",x"00",x"00"),
  1420 => (x"aa",x"b7",x"c0",x"79"),
  1421 => (x"87",x"f0",x"c3",x"03"),
  1422 => (x"00",x"1e",x"1c",x"27"),
  1423 => (x"27",x"4a",x"bf",x"00"),
  1424 => (x"00",x"00",x"1e",x"30"),
  1425 => (x"27",x"52",x"bf",x"97"),
  1426 => (x"00",x"00",x"1e",x"1c"),
  1427 => (x"82",x"c1",x"4a",x"bf"),
  1428 => (x"00",x"1e",x"1c",x"27"),
  1429 => (x"79",x"72",x"49",x"00"),
  1430 => (x"00",x"1e",x"34",x"27"),
  1431 => (x"aa",x"b7",x"bf",x"00"),
  1432 => (x"87",x"cd",x"c0",x"06"),
  1433 => (x"00",x"1e",x"34",x"27"),
  1434 => (x"1c",x"27",x"49",x"00"),
  1435 => (x"bf",x"00",x"00",x"1e"),
  1436 => (x"1e",x"2c",x"27",x"79"),
  1437 => (x"c1",x"49",x"00",x"00"),
  1438 => (x"87",x"ec",x"c2",x"79"),
  1439 => (x"00",x"1e",x"2c",x"27"),
  1440 => (x"c2",x"05",x"bf",x"00"),
  1441 => (x"30",x"27",x"87",x"e2"),
  1442 => (x"bf",x"00",x"00",x"1e"),
  1443 => (x"27",x"33",x"c4",x"4b"),
  1444 => (x"00",x"00",x"1e",x"30"),
  1445 => (x"27",x"79",x"73",x"49"),
  1446 => (x"00",x"00",x"1e",x"1c"),
  1447 => (x"52",x"73",x"4a",x"bf"),
  1448 => (x"27",x"87",x"c5",x"c2"),
  1449 => (x"00",x"00",x"1e",x"28"),
  1450 => (x"b7",x"c7",x"49",x"bf"),
  1451 => (x"e8",x"c1",x"04",x"a9"),
  1452 => (x"fe",x"4b",x"c0",x"87"),
  1453 => (x"79",x"c1",x"49",x"f4"),
  1454 => (x"00",x"1e",x"1c",x"27"),
  1455 => (x"79",x"c0",x"49",x"00"),
  1456 => (x"00",x"1e",x"34",x"27"),
  1457 => (x"c0",x"49",x"bf",x"00"),
  1458 => (x"c0",x"06",x"a9",x"b7"),
  1459 => (x"1c",x"27",x"87",x"e5"),
  1460 => (x"bf",x"00",x"00",x"1e"),
  1461 => (x"1c",x"27",x"83",x"bf"),
  1462 => (x"bf",x"00",x"00",x"1e"),
  1463 => (x"27",x"82",x"c4",x"4a"),
  1464 => (x"00",x"00",x"1e",x"1c"),
  1465 => (x"27",x"79",x"72",x"49"),
  1466 => (x"00",x"00",x"1e",x"34"),
  1467 => (x"04",x"aa",x"b7",x"bf"),
  1468 => (x"73",x"87",x"db",x"ff"),
  1469 => (x"1e",x"34",x"27",x"1e"),
  1470 => (x"1e",x"bf",x"00",x"00"),
  1471 => (x"00",x"1b",x"12",x"27"),
  1472 => (x"51",x"27",x"1e",x"00"),
  1473 => (x"0f",x"00",x"00",x"01"),
  1474 => (x"c0",x"ff",x"86",x"cc"),
  1475 => (x"79",x"c2",x"c1",x"49"),
  1476 => (x"00",x"14",x"2a",x"27"),
  1477 => (x"cf",x"c0",x"0f",x"00"),
  1478 => (x"1e",x"28",x"27",x"87"),
  1479 => (x"48",x"bf",x"00",x"00"),
  1480 => (x"ff",x"80",x"f0",x"c0"),
  1481 => (x"79",x"70",x"49",x"c0"),
  1482 => (x"4b",x"26",x"4c",x"26"),
  1483 => (x"4f",x"26",x"4a",x"26"),
  1484 => (x"87",x"fd",x"ff",x"1e"),
  1485 => (x"5e",x"0e",x"4f",x"26"),
  1486 => (x"5d",x"5c",x"5b",x"5a"),
  1487 => (x"19",x"1e",x"27",x"0e"),
  1488 => (x"27",x"1e",x"00",x"00"),
  1489 => (x"00",x"00",x"00",x"6e"),
  1490 => (x"27",x"86",x"c4",x"0f"),
  1491 => (x"00",x"00",x"06",x"60"),
  1492 => (x"72",x"4a",x"70",x"0f"),
  1493 => (x"ce",x"c4",x"02",x"9a"),
  1494 => (x"18",x"fb",x"27",x"87"),
  1495 => (x"27",x"1e",x"00",x"00"),
  1496 => (x"00",x"00",x"00",x"6e"),
  1497 => (x"27",x"86",x"c4",x"0f"),
  1498 => (x"00",x"00",x"0c",x"21"),
  1499 => (x"1e",x"38",x"27",x"0f"),
  1500 => (x"27",x"1e",x"00",x"00"),
  1501 => (x"00",x"00",x"19",x"12"),
  1502 => (x"12",x"d6",x"27",x"1e"),
  1503 => (x"c8",x"0f",x"00",x"00"),
  1504 => (x"72",x"4a",x"70",x"86"),
  1505 => (x"d0",x"c3",x"02",x"9a"),
  1506 => (x"1e",x"38",x"27",x"87"),
  1507 => (x"27",x"4b",x"00",x"00"),
  1508 => (x"00",x"00",x"18",x"d0"),
  1509 => (x"00",x"6e",x"27",x"1e"),
  1510 => (x"c4",x"0f",x"00",x"00"),
  1511 => (x"13",x"4d",x"c0",x"86"),
  1512 => (x"c0",x"4a",x"74",x"4c"),
  1513 => (x"02",x"aa",x"b7",x"e0"),
  1514 => (x"74",x"87",x"ed",x"c1"),
  1515 => (x"49",x"c0",x"ff",x"48"),
  1516 => (x"4a",x"74",x"79",x"70"),
  1517 => (x"aa",x"b7",x"e3",x"c0"),
  1518 => (x"87",x"dc",x"c1",x"02"),
  1519 => (x"c7",x"c1",x"4a",x"74"),
  1520 => (x"c0",x"05",x"aa",x"b7"),
  1521 => (x"2a",x"27",x"87",x"c6"),
  1522 => (x"0f",x"00",x"00",x"14"),
  1523 => (x"b7",x"ca",x"4a",x"74"),
  1524 => (x"c6",x"c0",x"05",x"aa"),
  1525 => (x"17",x"30",x"27",x"87"),
  1526 => (x"74",x"0f",x"00",x"00"),
  1527 => (x"b7",x"cc",x"c1",x"4a"),
  1528 => (x"c6",x"c0",x"05",x"aa"),
  1529 => (x"1e",x"38",x"27",x"87"),
  1530 => (x"74",x"4b",x"00",x"00"),
  1531 => (x"9a",x"df",x"ff",x"4a"),
  1532 => (x"4c",x"72",x"8a",x"d0"),
  1533 => (x"f9",x"c0",x"4a",x"74"),
  1534 => (x"c0",x"04",x"aa",x"b7"),
  1535 => (x"4a",x"74",x"87",x"c6"),
  1536 => (x"4c",x"72",x"8a",x"d1"),
  1537 => (x"4a",x"74",x"35",x"c4"),
  1538 => (x"b5",x"72",x"4d",x"75"),
  1539 => (x"4a",x"74",x"4c",x"13"),
  1540 => (x"aa",x"b7",x"e0",x"c0"),
  1541 => (x"87",x"d3",x"fe",x"05"),
  1542 => (x"e3",x"c0",x"4a",x"74"),
  1543 => (x"c0",x"02",x"aa",x"b7"),
  1544 => (x"4a",x"13",x"87",x"e2"),
  1545 => (x"aa",x"b7",x"e0",x"c0"),
  1546 => (x"87",x"ca",x"c0",x"05"),
  1547 => (x"e0",x"c0",x"4a",x"13"),
  1548 => (x"ff",x"02",x"aa",x"b7"),
  1549 => (x"8b",x"c1",x"87",x"f6"),
  1550 => (x"1e",x"73",x"1e",x"75"),
  1551 => (x"00",x"12",x"d6",x"27"),
  1552 => (x"86",x"c8",x"0f",x"00"),
  1553 => (x"b7",x"ca",x"4a",x"13"),
  1554 => (x"d0",x"fd",x"02",x"aa"),
  1555 => (x"ca",x"4a",x"13",x"87"),
  1556 => (x"ff",x"05",x"aa",x"b7"),
  1557 => (x"c4",x"fd",x"87",x"f7"),
  1558 => (x"18",x"e2",x"27",x"87"),
  1559 => (x"27",x"1e",x"00",x"00"),
  1560 => (x"00",x"00",x"00",x"6e"),
  1561 => (x"27",x"86",x"c4",x"0f"),
  1562 => (x"00",x"00",x"19",x"34"),
  1563 => (x"00",x"6e",x"27",x"1e"),
  1564 => (x"c4",x"0f",x"00",x"00"),
  1565 => (x"1e",x"34",x"27",x"86"),
  1566 => (x"c0",x"49",x"00",x"00"),
  1567 => (x"c8",x"f4",x"c3",x"79"),
  1568 => (x"ee",x"c0",x"4d",x"ff"),
  1569 => (x"00",x"4f",x"27",x"1e"),
  1570 => (x"c4",x"0f",x"00",x"00"),
  1571 => (x"c3",x"4b",x"75",x"86"),
  1572 => (x"4d",x"c0",x"c9",x"f4"),
  1573 => (x"4c",x"bf",x"c0",x"ff"),
  1574 => (x"c0",x"c8",x"4a",x"74"),
  1575 => (x"02",x"9a",x"72",x"9a"),
  1576 => (x"74",x"87",x"d1",x"c0"),
  1577 => (x"9a",x"ff",x"c3",x"4a"),
  1578 => (x"5d",x"27",x"1e",x"72"),
  1579 => (x"0f",x"00",x"00",x"14"),
  1580 => (x"4b",x"75",x"86",x"c4"),
  1581 => (x"8b",x"c1",x"4a",x"73"),
  1582 => (x"ff",x"05",x"9a",x"72"),
  1583 => (x"f4",x"c3",x"87",x"d6"),
  1584 => (x"fe",x"4d",x"ff",x"c8"),
  1585 => (x"4d",x"26",x"87",x"fc"),
  1586 => (x"4b",x"26",x"4c",x"26"),
  1587 => (x"4f",x"26",x"4a",x"26"),
  1588 => (x"73",x"72",x"61",x"50"),
  1589 => (x"20",x"67",x"6e",x"69"),
  1590 => (x"69",x"6e",x"61",x"6d"),
  1591 => (x"74",x"73",x"65",x"66"),
  1592 => (x"6f",x"4c",x"00",x"0a"),
  1593 => (x"6e",x"69",x"64",x"61"),
  1594 => (x"61",x"6d",x"20",x"67"),
  1595 => (x"65",x"66",x"69",x"6e"),
  1596 => (x"66",x"20",x"74",x"73"),
  1597 => (x"65",x"6c",x"69",x"61"),
  1598 => (x"48",x"00",x"0a",x"64"),
  1599 => (x"69",x"74",x"6e",x"75"),
  1600 => (x"66",x"20",x"67",x"6e"),
  1601 => (x"70",x"20",x"72",x"6f"),
  1602 => (x"69",x"74",x"72",x"61"),
  1603 => (x"6e",x"6f",x"69",x"74"),
  1604 => (x"41",x"4d",x"00",x"0a"),
  1605 => (x"45",x"46",x"49",x"4e"),
  1606 => (x"53",x"4d",x"54",x"53"),
  1607 => (x"6e",x"49",x"00",x"54"),
  1608 => (x"61",x"69",x"74",x"69"),
  1609 => (x"69",x"7a",x"69",x"6c"),
  1610 => (x"53",x"20",x"67",x"6e"),
  1611 => (x"61",x"63",x"20",x"44"),
  1612 => (x"00",x"0a",x"64",x"72"),
  1613 => (x"74",x"6f",x"6f",x"42"),
  1614 => (x"20",x"67",x"6e",x"69"),
  1615 => (x"6d",x"6f",x"72",x"66"),
  1616 => (x"32",x"53",x"52",x"20"),
  1617 => (x"00",x"2e",x"32",x"33"),
  1618 => (x"72",x"1e",x"73",x"1e"),
  1619 => (x"87",x"d9",x"02",x"9a"),
  1620 => (x"4b",x"c1",x"48",x"c0"),
  1621 => (x"82",x"01",x"a9",x"72"),
  1622 => (x"87",x"f8",x"83",x"73"),
  1623 => (x"89",x"03",x"a9",x"72"),
  1624 => (x"c1",x"07",x"80",x"73"),
  1625 => (x"f3",x"05",x"2b",x"2a"),
  1626 => (x"26",x"4b",x"26",x"87"),
  1627 => (x"1e",x"75",x"1e",x"4f"),
  1628 => (x"a1",x"71",x"4d",x"c0"),
  1629 => (x"c1",x"b9",x"ff",x"04"),
  1630 => (x"72",x"07",x"bd",x"81"),
  1631 => (x"ba",x"ff",x"04",x"a2"),
  1632 => (x"07",x"bd",x"82",x"c1"),
  1633 => (x"9d",x"75",x"87",x"c2"),
  1634 => (x"c1",x"b8",x"ff",x"05"),
  1635 => (x"4d",x"25",x"07",x"80"),
  1636 => (x"31",x"30",x"4f",x"26"),
  1637 => (x"35",x"34",x"33",x"32"),
  1638 => (x"39",x"38",x"37",x"36"),
  1639 => (x"44",x"43",x"42",x"41"),
  1640 => (x"43",x"00",x"46",x"45"),
  1641 => (x"52",x"00",x"44",x"4d"),
  1642 => (x"20",x"64",x"61",x"65"),
  1643 => (x"4d",x"20",x"66",x"6f"),
  1644 => (x"66",x"20",x"52",x"42"),
  1645 => (x"65",x"6c",x"69",x"61"),
  1646 => (x"4e",x"00",x"0a",x"64"),
  1647 => (x"61",x"70",x"20",x"6f"),
  1648 => (x"74",x"69",x"74",x"72"),
  1649 => (x"20",x"6e",x"6f",x"69"),
  1650 => (x"6e",x"67",x"69",x"73"),
  1651 => (x"72",x"75",x"74",x"61"),
  1652 => (x"6f",x"66",x"20",x"65"),
  1653 => (x"0a",x"64",x"6e",x"75"),
  1654 => (x"52",x"42",x"4d",x"00"),
  1655 => (x"65",x"7a",x"69",x"73"),
  1656 => (x"64",x"25",x"20",x"3a"),
  1657 => (x"61",x"70",x"20",x"2c"),
  1658 => (x"74",x"69",x"74",x"72"),
  1659 => (x"73",x"6e",x"6f",x"69"),
  1660 => (x"3a",x"65",x"7a",x"69"),
  1661 => (x"2c",x"64",x"25",x"20"),
  1662 => (x"66",x"66",x"6f",x"20"),
  1663 => (x"20",x"74",x"65",x"73"),
  1664 => (x"73",x"20",x"66",x"6f"),
  1665 => (x"20",x"3a",x"67",x"69"),
  1666 => (x"20",x"2c",x"64",x"25"),
  1667 => (x"20",x"67",x"69",x"73"),
  1668 => (x"78",x"25",x"78",x"30"),
  1669 => (x"65",x"52",x"00",x"0a"),
  1670 => (x"6e",x"69",x"64",x"61"),
  1671 => (x"6f",x"62",x"20",x"67"),
  1672 => (x"73",x"20",x"74",x"6f"),
  1673 => (x"6f",x"74",x"63",x"65"),
  1674 => (x"64",x"25",x"20",x"72"),
  1675 => (x"65",x"52",x"00",x"0a"),
  1676 => (x"62",x"20",x"64",x"61"),
  1677 => (x"20",x"74",x"6f",x"6f"),
  1678 => (x"74",x"63",x"65",x"73"),
  1679 => (x"66",x"20",x"72",x"6f"),
  1680 => (x"20",x"6d",x"6f",x"72"),
  1681 => (x"73",x"72",x"69",x"66"),
  1682 => (x"61",x"70",x"20",x"74"),
  1683 => (x"74",x"69",x"74",x"72"),
  1684 => (x"0a",x"6e",x"6f",x"69"),
  1685 => (x"73",x"6e",x"55",x"00"),
  1686 => (x"6f",x"70",x"70",x"75"),
  1687 => (x"64",x"65",x"74",x"72"),
  1688 => (x"72",x"61",x"70",x"20"),
  1689 => (x"69",x"74",x"69",x"74"),
  1690 => (x"74",x"20",x"6e",x"6f"),
  1691 => (x"21",x"65",x"70",x"79"),
  1692 => (x"41",x"46",x"00",x"0d"),
  1693 => (x"20",x"32",x"33",x"54"),
  1694 => (x"52",x"00",x"20",x"20"),
  1695 => (x"69",x"64",x"61",x"65"),
  1696 => (x"4d",x"20",x"67",x"6e"),
  1697 => (x"00",x"0a",x"52",x"42"),
  1698 => (x"20",x"52",x"42",x"4d"),
  1699 => (x"63",x"63",x"75",x"73"),
  1700 => (x"66",x"73",x"73",x"65"),
  1701 => (x"79",x"6c",x"6c",x"75"),
  1702 => (x"61",x"65",x"72",x"20"),
  1703 => (x"46",x"00",x"0a",x"64"),
  1704 => (x"36",x"31",x"54",x"41"),
  1705 => (x"00",x"20",x"20",x"20"),
  1706 => (x"33",x"54",x"41",x"46"),
  1707 => (x"20",x"20",x"20",x"32"),
  1708 => (x"72",x"61",x"50",x"00"),
  1709 => (x"69",x"74",x"69",x"74"),
  1710 => (x"6f",x"63",x"6e",x"6f"),
  1711 => (x"20",x"74",x"6e",x"75"),
  1712 => (x"00",x"0a",x"64",x"25"),
  1713 => (x"74",x"6e",x"75",x"48"),
  1714 => (x"20",x"67",x"6e",x"69"),
  1715 => (x"20",x"72",x"6f",x"66"),
  1716 => (x"65",x"6c",x"69",x"66"),
  1717 => (x"74",x"73",x"79",x"73"),
  1718 => (x"00",x"0a",x"6d",x"65"),
  1719 => (x"33",x"54",x"41",x"46"),
  1720 => (x"20",x"20",x"20",x"32"),
  1721 => (x"54",x"41",x"46",x"00"),
  1722 => (x"20",x"20",x"36",x"31"),
  1723 => (x"6c",x"43",x"00",x"20"),
  1724 => (x"65",x"74",x"73",x"75"),
  1725 => (x"69",x"73",x"20",x"72"),
  1726 => (x"20",x"3a",x"65",x"7a"),
  1727 => (x"20",x"2c",x"64",x"25"),
  1728 => (x"73",x"75",x"6c",x"43"),
  1729 => (x"20",x"72",x"65",x"74"),
  1730 => (x"6b",x"73",x"61",x"6d"),
  1731 => (x"64",x"25",x"20",x"2c"),
  1732 => (x"68",x"43",x"00",x"0a"),
  1733 => (x"73",x"6b",x"63",x"65"),
  1734 => (x"74",x"20",x"6d",x"75"),
  1735 => (x"64",x"25",x"20",x"6f"),
  1736 => (x"64",x"25",x"20",x"3a"),
  1737 => (x"64",x"25",x"00",x"0a"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
