
package Toplevel_Config is
	constant Toplevel_UseSDRAM : boolean := true;
	constant Toplevel_UseUART : boolean := false;
	constant Toplevel_UseVGA : boolean := true;
	constant Toplevel_UseAudio : boolean := true;
	constant Toplevel_Frequency : integer := 100;
end package;
