package Board_Config is
	constant Board_HaveSDRAM : boolean := true;
	constant Board_SDRAM_Width : integer := 32;
	constant Board_SDRAM_RowBits : integer := 13;
	constant Board_SDRAM_ColBits : integer := 9;
	constant Board_VGA_Bits : integer := 4;
	constant Board_JTAG_Uart : boolean := false;
end package;

