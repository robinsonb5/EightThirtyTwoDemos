
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"3b",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"38"),
    10 => (x"20",x"00",x"27",x"4f"),
    11 => (x"27",x"4e",x"00",x"00"),
    12 => (x"00",x"00",x"04",x"0a"),
    13 => (x"87",x"fd",x"00",x"0f"),
    14 => (x"4f",x"87",x"fd",x"00"),
    15 => (x"ff",x"86",x"fc",x"1e"),
    16 => (x"48",x"69",x"49",x"c0"),
    17 => (x"c4",x"98",x"c0",x"c4"),
    18 => (x"02",x"6e",x"58",x"a6"),
    19 => (x"66",x"c8",x"87",x"f4"),
    20 => (x"8e",x"fc",x"48",x"79"),
    21 => (x"5e",x"0e",x"4f",x"26"),
    22 => (x"0e",x"5d",x"5c",x"5b"),
    23 => (x"c0",x"4b",x"66",x"d0"),
    24 => (x"c3",x"49",x"13",x"4c"),
    25 => (x"99",x"71",x"99",x"ff"),
    26 => (x"71",x"87",x"db",x"02"),
    27 => (x"4a",x"c0",x"ff",x"4d"),
    28 => (x"c0",x"c4",x"49",x"6a"),
    29 => (x"87",x"f8",x"02",x"99"),
    30 => (x"84",x"c1",x"7a",x"75"),
    31 => (x"ff",x"c3",x"49",x"13"),
    32 => (x"05",x"99",x"71",x"99"),
    33 => (x"48",x"74",x"87",x"e5"),
    34 => (x"4c",x"26",x"4d",x"26"),
    35 => (x"4f",x"26",x"4b",x"26"),
    36 => (x"5c",x"5b",x"5e",x"0e"),
    37 => (x"86",x"e4",x"0e",x"5d"),
    38 => (x"4d",x"66",x"f4",x"c0"),
    39 => (x"c0",x"48",x"a6",x"c4"),
    40 => (x"c0",x"80",x"c4",x"78"),
    41 => (x"66",x"ec",x"c0",x"78"),
    42 => (x"fe",x"4b",x"bf",x"97"),
    43 => (x"c0",x"bb",x"83",x"c0"),
    44 => (x"c1",x"48",x"66",x"ec"),
    45 => (x"a6",x"f0",x"c0",x"80"),
    46 => (x"02",x"9b",x"73",x"58"),
    47 => (x"c8",x"87",x"f7",x"c7"),
    48 => (x"c0",x"c7",x"02",x"66"),
    49 => (x"48",x"a6",x"d0",x"87"),
    50 => (x"80",x"f8",x"78",x"c0"),
    51 => (x"f0",x"c0",x"78",x"c0"),
    52 => (x"ea",x"c2",x"02",x"ab"),
    53 => (x"ab",x"e3",x"c1",x"87"),
    54 => (x"87",x"eb",x"c2",x"02"),
    55 => (x"02",x"ab",x"e4",x"c1"),
    56 => (x"c1",x"87",x"e2",x"c0"),
    57 => (x"c2",x"02",x"ab",x"ec"),
    58 => (x"f0",x"c1",x"87",x"d5"),
    59 => (x"87",x"dd",x"02",x"ab"),
    60 => (x"02",x"ab",x"f3",x"c1"),
    61 => (x"f5",x"c1",x"87",x"df"),
    62 => (x"87",x"c9",x"02",x"ab"),
    63 => (x"02",x"ab",x"f8",x"c1"),
    64 => (x"e7",x"c2",x"87",x"cb"),
    65 => (x"48",x"a6",x"d0",x"87"),
    66 => (x"c2",x"c3",x"78",x"ca"),
    67 => (x"48",x"a6",x"d0",x"87"),
    68 => (x"fa",x"c2",x"78",x"d0"),
    69 => (x"66",x"f0",x"c0",x"87"),
    70 => (x"c0",x"80",x"c4",x"48"),
    71 => (x"c0",x"58",x"a6",x"f4"),
    72 => (x"c4",x"49",x"66",x"f0"),
    73 => (x"69",x"48",x"76",x"89"),
    74 => (x"ff",x"80",x"d4",x"78"),
    75 => (x"bf",x"97",x"6e",x"78"),
    76 => (x"80",x"c0",x"fe",x"48"),
    77 => (x"58",x"a6",x"dc",x"b8"),
    78 => (x"80",x"c1",x"48",x"6e"),
    79 => (x"d0",x"58",x"a6",x"c4"),
    80 => (x"66",x"d8",x"5b",x"a6"),
    81 => (x"87",x"e8",x"c0",x"02"),
    82 => (x"6e",x"4c",x"66",x"d8"),
    83 => (x"48",x"66",x"d4",x"4b"),
    84 => (x"a6",x"d8",x"80",x"c1"),
    85 => (x"66",x"f8",x"c0",x"58"),
    86 => (x"75",x"1e",x"74",x"1e"),
    87 => (x"74",x"86",x"c8",x"0f"),
    88 => (x"87",x"cc",x"05",x"a8"),
    89 => (x"c0",x"fe",x"4c",x"13"),
    90 => (x"9c",x"74",x"bc",x"84"),
    91 => (x"87",x"dd",x"ff",x"05"),
    92 => (x"d4",x"4b",x"66",x"cc"),
    93 => (x"66",x"c4",x"48",x"66"),
    94 => (x"58",x"a6",x"c8",x"80"),
    95 => (x"c8",x"87",x"d0",x"c1"),
    96 => (x"78",x"c1",x"48",x"a6"),
    97 => (x"c0",x"87",x"c8",x"c1"),
    98 => (x"c0",x"1e",x"66",x"f8"),
    99 => (x"c4",x"48",x"66",x"f4"),
   100 => (x"a6",x"f8",x"c0",x"80"),
   101 => (x"66",x"f4",x"c0",x"58"),
   102 => (x"69",x"89",x"c4",x"49"),
   103 => (x"c8",x"0f",x"75",x"1e"),
   104 => (x"48",x"66",x"c4",x"86"),
   105 => (x"a6",x"c8",x"80",x"c1"),
   106 => (x"87",x"e3",x"c0",x"58"),
   107 => (x"02",x"ab",x"e5",x"c0"),
   108 => (x"f8",x"c0",x"87",x"cb"),
   109 => (x"e5",x"c0",x"1e",x"66"),
   110 => (x"c8",x"0f",x"75",x"1e"),
   111 => (x"66",x"f8",x"c0",x"86"),
   112 => (x"75",x"1e",x"73",x"1e"),
   113 => (x"c4",x"86",x"c8",x"0f"),
   114 => (x"80",x"c1",x"48",x"66"),
   115 => (x"d0",x"58",x"a6",x"c8"),
   116 => (x"c7",x"c3",x"02",x"66"),
   117 => (x"66",x"f0",x"c0",x"87"),
   118 => (x"c0",x"80",x"c4",x"48"),
   119 => (x"c0",x"58",x"a6",x"f4"),
   120 => (x"c4",x"49",x"66",x"f0"),
   121 => (x"69",x"48",x"76",x"89"),
   122 => (x"ab",x"e4",x"c1",x"78"),
   123 => (x"6e",x"87",x"d8",x"05"),
   124 => (x"a8",x"b7",x"c0",x"48"),
   125 => (x"c0",x"87",x"d0",x"03"),
   126 => (x"ff",x"f8",x"1e",x"ed"),
   127 => (x"6e",x"86",x"c4",x"87"),
   128 => (x"88",x"08",x"c0",x"48"),
   129 => (x"6e",x"58",x"a6",x"c4"),
   130 => (x"e4",x"d8",x"c1",x"4a"),
   131 => (x"48",x"a6",x"cc",x"4c"),
   132 => (x"05",x"6e",x"78",x"c0"),
   133 => (x"d8",x"c1",x"87",x"ce"),
   134 => (x"d8",x"c1",x"4c",x"e5"),
   135 => (x"f0",x"c0",x"48",x"e4"),
   136 => (x"87",x"eb",x"c0",x"50"),
   137 => (x"e6",x"c0",x"02",x"6e"),
   138 => (x"4b",x"66",x"d0",x"87"),
   139 => (x"49",x"72",x"1e",x"72"),
   140 => (x"d8",x"c5",x"4a",x"73"),
   141 => (x"cd",x"4a",x"26",x"87"),
   142 => (x"54",x"11",x"81",x"fc"),
   143 => (x"49",x"72",x"1e",x"71"),
   144 => (x"c8",x"c5",x"4a",x"73"),
   145 => (x"26",x"4a",x"70",x"87"),
   146 => (x"05",x"9a",x"72",x"49"),
   147 => (x"c1",x"87",x"dd",x"ff"),
   148 => (x"02",x"ac",x"e4",x"d8"),
   149 => (x"c0",x"87",x"e3",x"c0"),
   150 => (x"c1",x"1e",x"66",x"f8"),
   151 => (x"49",x"6c",x"97",x"8c"),
   152 => (x"b9",x"81",x"c0",x"fe"),
   153 => (x"0f",x"75",x"1e",x"71"),
   154 => (x"66",x"cc",x"86",x"c8"),
   155 => (x"d0",x"80",x"c1",x"48"),
   156 => (x"d8",x"c1",x"58",x"a6"),
   157 => (x"ff",x"05",x"ac",x"e4"),
   158 => (x"66",x"cc",x"87",x"dd"),
   159 => (x"80",x"66",x"c4",x"48"),
   160 => (x"d7",x"58",x"a6",x"c8"),
   161 => (x"ab",x"e5",x"c0",x"87"),
   162 => (x"c8",x"87",x"c7",x"05"),
   163 => (x"78",x"c1",x"48",x"a6"),
   164 => (x"f8",x"c0",x"87",x"ca"),
   165 => (x"1e",x"73",x"1e",x"66"),
   166 => (x"86",x"c8",x"0f",x"75"),
   167 => (x"97",x"66",x"ec",x"c0"),
   168 => (x"c0",x"fe",x"4b",x"bf"),
   169 => (x"ec",x"c0",x"bb",x"83"),
   170 => (x"80",x"c1",x"48",x"66"),
   171 => (x"58",x"a6",x"f0",x"c0"),
   172 => (x"f8",x"05",x"9b",x"73"),
   173 => (x"66",x"c4",x"87",x"c9"),
   174 => (x"26",x"8e",x"e4",x"48"),
   175 => (x"26",x"4c",x"26",x"4d"),
   176 => (x"1e",x"4f",x"26",x"4b"),
   177 => (x"fc",x"c0",x"1e",x"c0"),
   178 => (x"1e",x"66",x"d0",x"1e"),
   179 => (x"f6",x"1e",x"66",x"d0"),
   180 => (x"86",x"d0",x"87",x"fe"),
   181 => (x"c0",x"1e",x"4f",x"26"),
   182 => (x"1e",x"fc",x"c0",x"1e"),
   183 => (x"d0",x"1e",x"a6",x"d0"),
   184 => (x"eb",x"f6",x"1e",x"66"),
   185 => (x"26",x"86",x"d0",x"87"),
   186 => (x"86",x"f8",x"1e",x"4f"),
   187 => (x"66",x"cc",x"48",x"76"),
   188 => (x"ff",x"80",x"c4",x"78"),
   189 => (x"cd",x"1e",x"76",x"78"),
   190 => (x"a6",x"dc",x"1e",x"cc"),
   191 => (x"1e",x"66",x"dc",x"1e"),
   192 => (x"d0",x"87",x"cd",x"f6"),
   193 => (x"26",x"8e",x"f8",x"86"),
   194 => (x"86",x"f8",x"1e",x"4f"),
   195 => (x"66",x"cc",x"48",x"76"),
   196 => (x"d0",x"80",x"c4",x"78"),
   197 => (x"1e",x"76",x"78",x"66"),
   198 => (x"c0",x"1e",x"cc",x"cd"),
   199 => (x"c0",x"1e",x"a6",x"e0"),
   200 => (x"f5",x"1e",x"66",x"e0"),
   201 => (x"86",x"d0",x"87",x"ea"),
   202 => (x"4f",x"26",x"8e",x"f8"),
   203 => (x"76",x"86",x"f8",x"1e"),
   204 => (x"78",x"66",x"cc",x"48"),
   205 => (x"78",x"ff",x"80",x"c4"),
   206 => (x"cc",x"cd",x"1e",x"76"),
   207 => (x"1e",x"66",x"dc",x"1e"),
   208 => (x"f5",x"1e",x"66",x"dc"),
   209 => (x"86",x"d0",x"87",x"ca"),
   210 => (x"4f",x"26",x"8e",x"f8"),
   211 => (x"4a",x"66",x"c8",x"1e"),
   212 => (x"02",x"6a",x"82",x"c4"),
   213 => (x"6a",x"87",x"e0",x"c0"),
   214 => (x"70",x"88",x"c1",x"48"),
   215 => (x"bf",x"66",x"c8",x"7a"),
   216 => (x"c1",x"48",x"71",x"49"),
   217 => (x"08",x"66",x"c8",x"80"),
   218 => (x"c4",x"97",x"08",x"78"),
   219 => (x"ff",x"c3",x"51",x"66"),
   220 => (x"48",x"66",x"c4",x"98"),
   221 => (x"c0",x"87",x"c2",x"c0"),
   222 => (x"00",x"4f",x"26",x"48"),
   223 => (x"33",x"32",x"31",x"30"),
   224 => (x"37",x"36",x"35",x"34"),
   225 => (x"42",x"41",x"39",x"38"),
   226 => (x"46",x"45",x"44",x"43"),
   227 => (x"1e",x"73",x"1e",x"00"),
   228 => (x"c0",x"02",x"9a",x"72"),
   229 => (x"48",x"c0",x"87",x"e7"),
   230 => (x"a9",x"72",x"4b",x"c1"),
   231 => (x"72",x"87",x"d1",x"06"),
   232 => (x"87",x"c9",x"06",x"82"),
   233 => (x"a9",x"72",x"83",x"73"),
   234 => (x"c3",x"87",x"f4",x"01"),
   235 => (x"3a",x"b2",x"c1",x"87"),
   236 => (x"89",x"03",x"a9",x"72"),
   237 => (x"c1",x"07",x"80",x"73"),
   238 => (x"f3",x"05",x"2b",x"2a"),
   239 => (x"26",x"4b",x"26",x"87"),
   240 => (x"1e",x"75",x"1e",x"4f"),
   241 => (x"b7",x"71",x"4d",x"c4"),
   242 => (x"b9",x"ff",x"04",x"a1"),
   243 => (x"bd",x"c3",x"81",x"c1"),
   244 => (x"a2",x"b7",x"72",x"07"),
   245 => (x"c1",x"ba",x"ff",x"04"),
   246 => (x"07",x"bd",x"c1",x"82"),
   247 => (x"c1",x"87",x"ee",x"fe"),
   248 => (x"b8",x"ff",x"04",x"2d"),
   249 => (x"2d",x"07",x"80",x"c1"),
   250 => (x"c1",x"b9",x"ff",x"04"),
   251 => (x"4d",x"26",x"07",x"81"),
   252 => (x"72",x"1e",x"4f",x"26"),
   253 => (x"11",x"48",x"12",x"1e"),
   254 => (x"88",x"87",x"c4",x"02"),
   255 => (x"26",x"87",x"f6",x"02"),
   256 => (x"1e",x"4f",x"26",x"4a"),
   257 => (x"48",x"bf",x"c8",x"ff"),
   258 => (x"5e",x"0e",x"4f",x"26"),
   259 => (x"0e",x"5d",x"5c",x"5b"),
   260 => (x"c1",x"86",x"dc",x"ff"),
   261 => (x"c3",x"48",x"f8",x"d8"),
   262 => (x"c1",x"78",x"fc",x"f8"),
   263 => (x"c3",x"48",x"f4",x"d8"),
   264 => (x"48",x"78",x"ec",x"f9"),
   265 => (x"78",x"fc",x"f8",x"c3"),
   266 => (x"48",x"f0",x"f9",x"c3"),
   267 => (x"80",x"c4",x"78",x"c0"),
   268 => (x"f9",x"c3",x"78",x"c2"),
   269 => (x"e8",x"c0",x"48",x"f8"),
   270 => (x"c3",x"1e",x"71",x"78"),
   271 => (x"c0",x"49",x"fc",x"f9"),
   272 => (x"20",x"48",x"d0",x"f6"),
   273 => (x"20",x"41",x"20",x"41"),
   274 => (x"20",x"41",x"20",x"41"),
   275 => (x"20",x"41",x"20",x"41"),
   276 => (x"10",x"51",x"10",x"41"),
   277 => (x"26",x"51",x"10",x"51"),
   278 => (x"c3",x"1e",x"71",x"49"),
   279 => (x"c0",x"49",x"dc",x"fa"),
   280 => (x"20",x"48",x"f0",x"f6"),
   281 => (x"20",x"41",x"20",x"41"),
   282 => (x"20",x"41",x"20",x"41"),
   283 => (x"20",x"41",x"20",x"41"),
   284 => (x"10",x"51",x"10",x"41"),
   285 => (x"26",x"51",x"10",x"51"),
   286 => (x"f0",x"f5",x"c1",x"49"),
   287 => (x"c0",x"78",x"ca",x"48"),
   288 => (x"f9",x"1e",x"d0",x"f7"),
   289 => (x"86",x"c4",x"87",x"d0"),
   290 => (x"1e",x"d4",x"f7",x"c0"),
   291 => (x"c4",x"87",x"c7",x"f9"),
   292 => (x"c4",x"f8",x"c0",x"86"),
   293 => (x"87",x"fe",x"f8",x"1e"),
   294 => (x"ef",x"c0",x"86",x"c4"),
   295 => (x"d4",x"02",x"bf",x"f4"),
   296 => (x"fc",x"ef",x"c0",x"87"),
   297 => (x"87",x"ee",x"f8",x"1e"),
   298 => (x"f0",x"c0",x"86",x"c4"),
   299 => (x"e5",x"f8",x"1e",x"e8"),
   300 => (x"d2",x"86",x"c4",x"87"),
   301 => (x"ec",x"f0",x"c0",x"87"),
   302 => (x"87",x"da",x"f8",x"1e"),
   303 => (x"f1",x"c0",x"86",x"c4"),
   304 => (x"d1",x"f8",x"1e",x"dc"),
   305 => (x"c0",x"86",x"c4",x"87"),
   306 => (x"1e",x"bf",x"f8",x"ef"),
   307 => (x"1e",x"c8",x"f8",x"c0"),
   308 => (x"c8",x"87",x"c3",x"f8"),
   309 => (x"e4",x"f8",x"c3",x"86"),
   310 => (x"bf",x"c8",x"ff",x"48"),
   311 => (x"48",x"a6",x"c8",x"78"),
   312 => (x"ef",x"c0",x"78",x"c1"),
   313 => (x"c0",x"48",x"bf",x"f8"),
   314 => (x"c9",x"06",x"a8",x"b7"),
   315 => (x"a6",x"cc",x"87",x"dd"),
   316 => (x"58",x"a6",x"d4",x"48"),
   317 => (x"a6",x"dc",x"80",x"c8"),
   318 => (x"48",x"a6",x"dc",x"58"),
   319 => (x"c1",x"58",x"a6",x"c8"),
   320 => (x"c1",x"48",x"c4",x"d9"),
   321 => (x"d9",x"c1",x"50",x"c1"),
   322 => (x"78",x"c0",x"48",x"c0"),
   323 => (x"97",x"c4",x"d9",x"c1"),
   324 => (x"c0",x"fe",x"49",x"bf"),
   325 => (x"c1",x"c1",x"b9",x"81"),
   326 => (x"c7",x"c0",x"02",x"a9"),
   327 => (x"c0",x"48",x"76",x"87"),
   328 => (x"87",x"c4",x"c0",x"78"),
   329 => (x"78",x"c1",x"48",x"76"),
   330 => (x"bf",x"c0",x"d9",x"c1"),
   331 => (x"c1",x"b0",x"6e",x"48"),
   332 => (x"c1",x"58",x"c4",x"d9"),
   333 => (x"c1",x"48",x"c8",x"d9"),
   334 => (x"a6",x"dc",x"50",x"c2"),
   335 => (x"c4",x"78",x"c2",x"48"),
   336 => (x"c3",x"78",x"c3",x"80"),
   337 => (x"c0",x"49",x"fc",x"fa"),
   338 => (x"20",x"48",x"c0",x"f2"),
   339 => (x"20",x"41",x"20",x"41"),
   340 => (x"20",x"41",x"20",x"41"),
   341 => (x"20",x"41",x"20",x"41"),
   342 => (x"10",x"51",x"10",x"41"),
   343 => (x"d4",x"51",x"10",x"51"),
   344 => (x"78",x"c1",x"48",x"a6"),
   345 => (x"1e",x"fc",x"fa",x"c3"),
   346 => (x"1e",x"dc",x"fa",x"c3"),
   347 => (x"87",x"ed",x"c0",x"c1"),
   348 => (x"98",x"70",x"86",x"c8"),
   349 => (x"87",x"c5",x"c0",x"05"),
   350 => (x"c2",x"c0",x"49",x"c1"),
   351 => (x"c1",x"49",x"c0",x"87"),
   352 => (x"dc",x"59",x"c4",x"d9"),
   353 => (x"b7",x"c3",x"48",x"66"),
   354 => (x"ef",x"c0",x"03",x"a8"),
   355 => (x"49",x"66",x"dc",x"87"),
   356 => (x"71",x"91",x"b7",x"c5"),
   357 => (x"d0",x"88",x"c3",x"48"),
   358 => (x"66",x"d0",x"58",x"a6"),
   359 => (x"c0",x"1e",x"c3",x"1e"),
   360 => (x"c0",x"1e",x"66",x"e4"),
   361 => (x"cc",x"87",x"ce",x"fc"),
   362 => (x"48",x"66",x"dc",x"86"),
   363 => (x"e0",x"c0",x"80",x"c1"),
   364 => (x"66",x"dc",x"58",x"a6"),
   365 => (x"a8",x"b7",x"c3",x"48"),
   366 => (x"87",x"d1",x"ff",x"04"),
   367 => (x"c0",x"1e",x"66",x"cc"),
   368 => (x"c1",x"1e",x"66",x"e0"),
   369 => (x"c1",x"1e",x"d4",x"dc"),
   370 => (x"c0",x"1e",x"cc",x"d9"),
   371 => (x"d0",x"87",x"f8",x"fb"),
   372 => (x"f4",x"d8",x"c1",x"86"),
   373 => (x"d8",x"c1",x"4c",x"bf"),
   374 => (x"4b",x"bf",x"bf",x"f4"),
   375 => (x"49",x"73",x"1e",x"72"),
   376 => (x"bf",x"f4",x"d8",x"c1"),
   377 => (x"a1",x"f0",x"c0",x"48"),
   378 => (x"71",x"41",x"20",x"4a"),
   379 => (x"f8",x"ff",x"05",x"aa"),
   380 => (x"74",x"4a",x"26",x"87"),
   381 => (x"c4",x"80",x"c8",x"48"),
   382 => (x"49",x"74",x"58",x"a6"),
   383 => (x"79",x"c5",x"81",x"cc"),
   384 => (x"85",x"cc",x"4d",x"73"),
   385 => (x"7b",x"6c",x"7d",x"69"),
   386 => (x"fa",x"d6",x"1e",x"73"),
   387 => (x"73",x"86",x"c4",x"87"),
   388 => (x"69",x"81",x"c4",x"49"),
   389 => (x"87",x"e7",x"c0",x"05"),
   390 => (x"81",x"c8",x"49",x"73"),
   391 => (x"1e",x"71",x"7d",x"c6"),
   392 => (x"1e",x"bf",x"66",x"c4"),
   393 => (x"87",x"df",x"f8",x"c0"),
   394 => (x"d8",x"c1",x"86",x"c8"),
   395 => (x"7b",x"bf",x"bf",x"f4"),
   396 => (x"1e",x"ca",x"1e",x"75"),
   397 => (x"f9",x"c0",x"1e",x"6d"),
   398 => (x"86",x"cc",x"87",x"fb"),
   399 => (x"6c",x"87",x"d9",x"c0"),
   400 => (x"72",x"1e",x"71",x"49"),
   401 => (x"48",x"49",x"74",x"1e"),
   402 => (x"4a",x"a1",x"f0",x"c0"),
   403 => (x"aa",x"71",x"41",x"20"),
   404 => (x"87",x"f8",x"ff",x"05"),
   405 => (x"49",x"26",x"4a",x"26"),
   406 => (x"c1",x"c1",x"48",x"76"),
   407 => (x"c8",x"d9",x"c1",x"50"),
   408 => (x"fe",x"49",x"bf",x"97"),
   409 => (x"c1",x"b9",x"81",x"c0"),
   410 => (x"04",x"a9",x"b7",x"c1"),
   411 => (x"97",x"87",x"ed",x"c1"),
   412 => (x"c3",x"c1",x"4b",x"6e"),
   413 => (x"fe",x"49",x"73",x"1e"),
   414 => (x"71",x"b9",x"81",x"c0"),
   415 => (x"f1",x"fb",x"c0",x"1e"),
   416 => (x"d4",x"86",x"c8",x"87"),
   417 => (x"c0",x"05",x"a8",x"66"),
   418 => (x"66",x"d8",x"87",x"f9"),
   419 => (x"c0",x"1e",x"c0",x"1e"),
   420 => (x"c8",x"87",x"f4",x"f6"),
   421 => (x"c3",x"1e",x"71",x"86"),
   422 => (x"c0",x"49",x"fc",x"fa"),
   423 => (x"20",x"48",x"e0",x"f1"),
   424 => (x"20",x"41",x"20",x"41"),
   425 => (x"20",x"41",x"20",x"41"),
   426 => (x"20",x"41",x"20",x"41"),
   427 => (x"10",x"51",x"10",x"41"),
   428 => (x"26",x"51",x"10",x"51"),
   429 => (x"a6",x"e0",x"c0",x"49"),
   430 => (x"78",x"66",x"c8",x"48"),
   431 => (x"48",x"fc",x"d8",x"c1"),
   432 => (x"c1",x"78",x"66",x"c8"),
   433 => (x"fe",x"4a",x"73",x"83"),
   434 => (x"c1",x"ba",x"82",x"c0"),
   435 => (x"bf",x"97",x"c8",x"d9"),
   436 => (x"81",x"c0",x"fe",x"49"),
   437 => (x"aa",x"b7",x"71",x"b9"),
   438 => (x"87",x"d6",x"fe",x"06"),
   439 => (x"48",x"66",x"e0",x"c0"),
   440 => (x"90",x"b7",x"66",x"dc"),
   441 => (x"58",x"a6",x"e4",x"c0"),
   442 => (x"1e",x"72",x"1e",x"71"),
   443 => (x"49",x"66",x"e8",x"c0"),
   444 => (x"f3",x"4a",x"66",x"d4"),
   445 => (x"4a",x"26",x"87",x"cb"),
   446 => (x"e0",x"c0",x"49",x"26"),
   447 => (x"e0",x"c0",x"58",x"a6"),
   448 => (x"66",x"cc",x"49",x"66"),
   449 => (x"91",x"b7",x"c7",x"89"),
   450 => (x"66",x"dc",x"48",x"71"),
   451 => (x"a6",x"e4",x"c0",x"88"),
   452 => (x"bf",x"66",x"c4",x"58"),
   453 => (x"c1",x"82",x"ca",x"4a"),
   454 => (x"bf",x"97",x"c4",x"d9"),
   455 => (x"81",x"c0",x"fe",x"49"),
   456 => (x"a9",x"c1",x"c1",x"b9"),
   457 => (x"87",x"ce",x"c0",x"05"),
   458 => (x"48",x"72",x"8a",x"c1"),
   459 => (x"bf",x"fc",x"d8",x"c1"),
   460 => (x"08",x"66",x"c4",x"88"),
   461 => (x"66",x"c8",x"08",x"78"),
   462 => (x"cc",x"80",x"c1",x"48"),
   463 => (x"66",x"c8",x"58",x"a6"),
   464 => (x"f8",x"ef",x"c0",x"48"),
   465 => (x"06",x"a8",x"b7",x"bf"),
   466 => (x"c3",x"87",x"f4",x"f6"),
   467 => (x"ff",x"48",x"e8",x"f8"),
   468 => (x"c0",x"78",x"bf",x"c8"),
   469 => (x"ed",x"1e",x"f8",x"f8"),
   470 => (x"86",x"c4",x"87",x"fc"),
   471 => (x"1e",x"c8",x"f9",x"c0"),
   472 => (x"c4",x"87",x"f3",x"ed"),
   473 => (x"cc",x"f9",x"c0",x"86"),
   474 => (x"87",x"ea",x"ed",x"1e"),
   475 => (x"fa",x"c0",x"86",x"c4"),
   476 => (x"e1",x"ed",x"1e",x"c4"),
   477 => (x"c1",x"86",x"c4",x"87"),
   478 => (x"1e",x"bf",x"fc",x"d8"),
   479 => (x"1e",x"c8",x"fa",x"c0"),
   480 => (x"c8",x"87",x"d3",x"ed"),
   481 => (x"c0",x"1e",x"c5",x"86"),
   482 => (x"ed",x"1e",x"e4",x"fa"),
   483 => (x"86",x"c8",x"87",x"c8"),
   484 => (x"bf",x"c0",x"d9",x"c1"),
   485 => (x"c0",x"fb",x"c0",x"1e"),
   486 => (x"87",x"fa",x"ec",x"1e"),
   487 => (x"1e",x"c1",x"86",x"c8"),
   488 => (x"1e",x"dc",x"fb",x"c0"),
   489 => (x"c8",x"87",x"ef",x"ec"),
   490 => (x"c4",x"d9",x"c1",x"86"),
   491 => (x"fe",x"49",x"bf",x"97"),
   492 => (x"71",x"b9",x"81",x"c0"),
   493 => (x"f8",x"fb",x"c0",x"1e"),
   494 => (x"87",x"da",x"ec",x"1e"),
   495 => (x"c1",x"c1",x"86",x"c8"),
   496 => (x"d4",x"fc",x"c0",x"1e"),
   497 => (x"87",x"ce",x"ec",x"1e"),
   498 => (x"d9",x"c1",x"86",x"c8"),
   499 => (x"49",x"bf",x"97",x"c8"),
   500 => (x"b9",x"81",x"c0",x"fe"),
   501 => (x"fc",x"c0",x"1e",x"71"),
   502 => (x"f9",x"eb",x"1e",x"f0"),
   503 => (x"c1",x"86",x"c8",x"87"),
   504 => (x"fd",x"c0",x"1e",x"c2"),
   505 => (x"ed",x"eb",x"1e",x"cc"),
   506 => (x"c1",x"86",x"c8",x"87"),
   507 => (x"1e",x"bf",x"ec",x"d9"),
   508 => (x"1e",x"e8",x"fd",x"c0"),
   509 => (x"c8",x"87",x"df",x"eb"),
   510 => (x"c0",x"1e",x"c7",x"86"),
   511 => (x"eb",x"1e",x"c4",x"fe"),
   512 => (x"86",x"c8",x"87",x"d4"),
   513 => (x"bf",x"f0",x"f5",x"c1"),
   514 => (x"e0",x"fe",x"c0",x"1e"),
   515 => (x"87",x"c6",x"eb",x"1e"),
   516 => (x"fe",x"c0",x"86",x"c8"),
   517 => (x"fd",x"ea",x"1e",x"fc"),
   518 => (x"c0",x"86",x"c4",x"87"),
   519 => (x"ea",x"1e",x"e8",x"ff"),
   520 => (x"86",x"c4",x"87",x"f4"),
   521 => (x"bf",x"f4",x"d8",x"c1"),
   522 => (x"ff",x"c0",x"1e",x"bf"),
   523 => (x"e5",x"ea",x"1e",x"f4"),
   524 => (x"c1",x"86",x"c8",x"87"),
   525 => (x"ea",x"1e",x"d0",x"c0"),
   526 => (x"86",x"c4",x"87",x"dc"),
   527 => (x"bf",x"f4",x"d8",x"c1"),
   528 => (x"69",x"81",x"c4",x"49"),
   529 => (x"c4",x"c1",x"c1",x"1e"),
   530 => (x"87",x"ca",x"ea",x"1e"),
   531 => (x"1e",x"c0",x"86",x"c8"),
   532 => (x"1e",x"e0",x"c1",x"c1"),
   533 => (x"c8",x"87",x"ff",x"e9"),
   534 => (x"f4",x"d8",x"c1",x"86"),
   535 => (x"81",x"c8",x"49",x"bf"),
   536 => (x"c1",x"c1",x"1e",x"69"),
   537 => (x"ed",x"e9",x"1e",x"fc"),
   538 => (x"c2",x"86",x"c8",x"87"),
   539 => (x"d8",x"c2",x"c1",x"1e"),
   540 => (x"87",x"e2",x"e9",x"1e"),
   541 => (x"d8",x"c1",x"86",x"c8"),
   542 => (x"cc",x"49",x"bf",x"f4"),
   543 => (x"c1",x"1e",x"69",x"81"),
   544 => (x"e9",x"1e",x"f4",x"c2"),
   545 => (x"86",x"c8",x"87",x"d0"),
   546 => (x"c3",x"c1",x"1e",x"d1"),
   547 => (x"c5",x"e9",x"1e",x"d0"),
   548 => (x"c1",x"86",x"c8",x"87"),
   549 => (x"49",x"bf",x"f4",x"d8"),
   550 => (x"1e",x"71",x"81",x"d0"),
   551 => (x"1e",x"ec",x"c3",x"c1"),
   552 => (x"c8",x"87",x"f3",x"e8"),
   553 => (x"c8",x"c4",x"c1",x"86"),
   554 => (x"87",x"ea",x"e8",x"1e"),
   555 => (x"c5",x"c1",x"86",x"c4"),
   556 => (x"e1",x"e8",x"1e",x"c0"),
   557 => (x"c1",x"86",x"c4",x"87"),
   558 => (x"bf",x"bf",x"f8",x"d8"),
   559 => (x"d4",x"c5",x"c1",x"1e"),
   560 => (x"87",x"d2",x"e8",x"1e"),
   561 => (x"c5",x"c1",x"86",x"c8"),
   562 => (x"c9",x"e8",x"1e",x"f0"),
   563 => (x"c1",x"86",x"c4",x"87"),
   564 => (x"49",x"bf",x"f8",x"d8"),
   565 => (x"1e",x"69",x"81",x"c4"),
   566 => (x"1e",x"f0",x"c6",x"c1"),
   567 => (x"c8",x"87",x"f7",x"e7"),
   568 => (x"c1",x"1e",x"c0",x"86"),
   569 => (x"e7",x"1e",x"cc",x"c7"),
   570 => (x"86",x"c8",x"87",x"ec"),
   571 => (x"bf",x"f8",x"d8",x"c1"),
   572 => (x"69",x"81",x"c8",x"49"),
   573 => (x"e8",x"c7",x"c1",x"1e"),
   574 => (x"87",x"da",x"e7",x"1e"),
   575 => (x"1e",x"c1",x"86",x"c8"),
   576 => (x"1e",x"c4",x"c8",x"c1"),
   577 => (x"c8",x"87",x"cf",x"e7"),
   578 => (x"f8",x"d8",x"c1",x"86"),
   579 => (x"81",x"cc",x"49",x"bf"),
   580 => (x"c8",x"c1",x"1e",x"69"),
   581 => (x"fd",x"e6",x"1e",x"e0"),
   582 => (x"d2",x"86",x"c8",x"87"),
   583 => (x"fc",x"c8",x"c1",x"1e"),
   584 => (x"87",x"f2",x"e6",x"1e"),
   585 => (x"d8",x"c1",x"86",x"c8"),
   586 => (x"d0",x"49",x"bf",x"f8"),
   587 => (x"c1",x"1e",x"71",x"81"),
   588 => (x"e6",x"1e",x"d8",x"c9"),
   589 => (x"86",x"c8",x"87",x"e0"),
   590 => (x"1e",x"f4",x"c9",x"c1"),
   591 => (x"c4",x"87",x"d7",x"e6"),
   592 => (x"1e",x"66",x"dc",x"86"),
   593 => (x"1e",x"ec",x"ca",x"c1"),
   594 => (x"c8",x"87",x"cb",x"e6"),
   595 => (x"c1",x"1e",x"c5",x"86"),
   596 => (x"e6",x"1e",x"c8",x"cb"),
   597 => (x"86",x"c8",x"87",x"c0"),
   598 => (x"1e",x"66",x"e0",x"c0"),
   599 => (x"1e",x"e4",x"cb",x"c1"),
   600 => (x"c8",x"87",x"f3",x"e5"),
   601 => (x"c1",x"1e",x"cd",x"86"),
   602 => (x"e5",x"1e",x"c0",x"cc"),
   603 => (x"86",x"c8",x"87",x"e8"),
   604 => (x"c1",x"1e",x"66",x"cc"),
   605 => (x"e5",x"1e",x"dc",x"cc"),
   606 => (x"86",x"c8",x"87",x"dc"),
   607 => (x"cc",x"c1",x"1e",x"c7"),
   608 => (x"d1",x"e5",x"1e",x"f8"),
   609 => (x"d4",x"86",x"c8",x"87"),
   610 => (x"cd",x"c1",x"1e",x"66"),
   611 => (x"c5",x"e5",x"1e",x"d4"),
   612 => (x"c1",x"86",x"c8",x"87"),
   613 => (x"f0",x"cd",x"c1",x"1e"),
   614 => (x"87",x"fa",x"e4",x"1e"),
   615 => (x"fa",x"c3",x"86",x"c8"),
   616 => (x"ce",x"c1",x"1e",x"dc"),
   617 => (x"ed",x"e4",x"1e",x"cc"),
   618 => (x"c1",x"86",x"c8",x"87"),
   619 => (x"e4",x"1e",x"e8",x"ce"),
   620 => (x"86",x"c4",x"87",x"e4"),
   621 => (x"1e",x"fc",x"fa",x"c3"),
   622 => (x"1e",x"e0",x"cf",x"c1"),
   623 => (x"c8",x"87",x"d7",x"e4"),
   624 => (x"fc",x"cf",x"c1",x"86"),
   625 => (x"87",x"ce",x"e4",x"1e"),
   626 => (x"d0",x"c1",x"86",x"c4"),
   627 => (x"c5",x"e4",x"1e",x"f4"),
   628 => (x"c3",x"86",x"c4",x"87"),
   629 => (x"49",x"bf",x"e8",x"f8"),
   630 => (x"bf",x"e4",x"f8",x"c3"),
   631 => (x"f0",x"f8",x"c3",x"89"),
   632 => (x"c1",x"1e",x"71",x"59"),
   633 => (x"e3",x"1e",x"f8",x"d0"),
   634 => (x"86",x"c8",x"87",x"ec"),
   635 => (x"bf",x"ec",x"f8",x"c3"),
   636 => (x"b7",x"f8",x"c1",x"48"),
   637 => (x"db",x"c0",x"03",x"a8"),
   638 => (x"e0",x"f2",x"c0",x"87"),
   639 => (x"87",x"d6",x"e3",x"1e"),
   640 => (x"f3",x"c0",x"86",x"c4"),
   641 => (x"cd",x"e3",x"1e",x"d8"),
   642 => (x"c0",x"86",x"c4",x"87"),
   643 => (x"e3",x"1e",x"f8",x"f3"),
   644 => (x"86",x"c4",x"87",x"c4"),
   645 => (x"bf",x"ec",x"f8",x"c3"),
   646 => (x"cf",x"4a",x"71",x"49"),
   647 => (x"71",x"92",x"b7",x"e8"),
   648 => (x"72",x"1e",x"72",x"1e"),
   649 => (x"f8",x"ef",x"c0",x"49"),
   650 => (x"d4",x"e6",x"4a",x"bf"),
   651 => (x"26",x"4a",x"26",x"87"),
   652 => (x"f4",x"f8",x"c3",x"49"),
   653 => (x"f8",x"ef",x"c0",x"58"),
   654 => (x"4b",x"72",x"4a",x"bf"),
   655 => (x"93",x"b7",x"e8",x"cf"),
   656 => (x"1e",x"72",x"1e",x"71"),
   657 => (x"e5",x"4a",x"09",x"73"),
   658 => (x"4a",x"26",x"87",x"f7"),
   659 => (x"f8",x"c3",x"49",x"26"),
   660 => (x"f9",x"c8",x"58",x"f8"),
   661 => (x"1e",x"71",x"92",x"b7"),
   662 => (x"09",x"72",x"1e",x"72"),
   663 => (x"87",x"e1",x"e5",x"4a"),
   664 => (x"49",x"26",x"4a",x"26"),
   665 => (x"58",x"fc",x"f8",x"c3"),
   666 => (x"1e",x"fc",x"f3",x"c0"),
   667 => (x"c4",x"87",x"e7",x"e1"),
   668 => (x"f0",x"f8",x"c3",x"86"),
   669 => (x"f4",x"c0",x"1e",x"bf"),
   670 => (x"d9",x"e1",x"1e",x"ec"),
   671 => (x"c0",x"86",x"c8",x"87"),
   672 => (x"e1",x"1e",x"f4",x"f4"),
   673 => (x"86",x"c4",x"87",x"d0"),
   674 => (x"bf",x"f4",x"f8",x"c3"),
   675 => (x"e4",x"f5",x"c0",x"1e"),
   676 => (x"87",x"c2",x"e1",x"1e"),
   677 => (x"f8",x"c3",x"86",x"c8"),
   678 => (x"c0",x"1e",x"bf",x"f8"),
   679 => (x"e0",x"1e",x"ec",x"f5"),
   680 => (x"86",x"c8",x"87",x"f4"),
   681 => (x"1e",x"cc",x"f6",x"c0"),
   682 => (x"c4",x"87",x"eb",x"e0"),
   683 => (x"ff",x"48",x"c0",x"86"),
   684 => (x"4d",x"26",x"8e",x"dc"),
   685 => (x"4b",x"26",x"4c",x"26"),
   686 => (x"c1",x"1e",x"4f",x"26"),
   687 => (x"c1",x"48",x"c4",x"d9"),
   688 => (x"d9",x"c1",x"50",x"c1"),
   689 => (x"78",x"c0",x"48",x"c0"),
   690 => (x"c1",x"1e",x"4f",x"26"),
   691 => (x"bf",x"97",x"c4",x"d9"),
   692 => (x"81",x"c0",x"fe",x"49"),
   693 => (x"a9",x"c1",x"c1",x"b9"),
   694 => (x"87",x"c5",x"c0",x"02"),
   695 => (x"c2",x"c0",x"49",x"c0"),
   696 => (x"c1",x"49",x"c1",x"87"),
   697 => (x"48",x"bf",x"c0",x"d9"),
   698 => (x"d9",x"c1",x"b0",x"71"),
   699 => (x"d9",x"c1",x"58",x"c4"),
   700 => (x"c2",x"c1",x"48",x"c8"),
   701 => (x"0e",x"4f",x"26",x"50"),
   702 => (x"5d",x"5c",x"5b",x"5e"),
   703 => (x"d4",x"86",x"fc",x"0e"),
   704 => (x"4b",x"6d",x"4d",x"66"),
   705 => (x"d8",x"c1",x"49",x"73"),
   706 => (x"c0",x"48",x"bf",x"f4"),
   707 => (x"20",x"4a",x"a1",x"f0"),
   708 => (x"05",x"aa",x"71",x"41"),
   709 => (x"75",x"87",x"f8",x"ff"),
   710 => (x"c4",x"80",x"c8",x"48"),
   711 => (x"49",x"75",x"58",x"a6"),
   712 => (x"79",x"c5",x"81",x"cc"),
   713 => (x"84",x"cc",x"4c",x"73"),
   714 => (x"7b",x"6d",x"7c",x"c5"),
   715 => (x"bf",x"f4",x"d8",x"c1"),
   716 => (x"87",x"c6",x"c0",x"02"),
   717 => (x"bf",x"f4",x"d8",x"c1"),
   718 => (x"d8",x"c1",x"7b",x"bf"),
   719 => (x"cc",x"49",x"bf",x"f4"),
   720 => (x"c1",x"1e",x"71",x"81"),
   721 => (x"1e",x"bf",x"fc",x"d8"),
   722 => (x"e5",x"c0",x"1e",x"ca"),
   723 => (x"86",x"cc",x"87",x"e7"),
   724 => (x"81",x"c4",x"49",x"73"),
   725 => (x"e7",x"c0",x"05",x"69"),
   726 => (x"c8",x"49",x"73",x"87"),
   727 => (x"71",x"7c",x"c6",x"81"),
   728 => (x"bf",x"66",x"c4",x"1e"),
   729 => (x"de",x"e3",x"c0",x"1e"),
   730 => (x"c1",x"86",x"c8",x"87"),
   731 => (x"bf",x"bf",x"f4",x"d8"),
   732 => (x"ca",x"1e",x"74",x"7b"),
   733 => (x"c0",x"1e",x"6c",x"1e"),
   734 => (x"cc",x"87",x"fa",x"e4"),
   735 => (x"87",x"d5",x"c0",x"86"),
   736 => (x"1e",x"71",x"49",x"6d"),
   737 => (x"c0",x"48",x"49",x"75"),
   738 => (x"20",x"4a",x"a1",x"f0"),
   739 => (x"05",x"aa",x"71",x"41"),
   740 => (x"26",x"87",x"f8",x"ff"),
   741 => (x"26",x"8e",x"fc",x"49"),
   742 => (x"26",x"4c",x"26",x"4d"),
   743 => (x"1e",x"4f",x"26",x"4b"),
   744 => (x"4a",x"bf",x"66",x"c4"),
   745 => (x"d9",x"c1",x"82",x"ca"),
   746 => (x"49",x"bf",x"97",x"c4"),
   747 => (x"b9",x"81",x"c0",x"fe"),
   748 => (x"05",x"a9",x"c1",x"c1"),
   749 => (x"c1",x"87",x"ce",x"c0"),
   750 => (x"c1",x"48",x"72",x"8a"),
   751 => (x"88",x"bf",x"fc",x"d8"),
   752 => (x"78",x"08",x"66",x"c4"),
   753 => (x"1e",x"4f",x"26",x"08"),
   754 => (x"bf",x"f4",x"d8",x"c1"),
   755 => (x"87",x"c9",x"c0",x"02"),
   756 => (x"c1",x"48",x"66",x"c4"),
   757 => (x"bf",x"bf",x"f4",x"d8"),
   758 => (x"f4",x"d8",x"c1",x"78"),
   759 => (x"81",x"cc",x"49",x"bf"),
   760 => (x"d8",x"c1",x"1e",x"71"),
   761 => (x"ca",x"1e",x"bf",x"fc"),
   762 => (x"c8",x"e3",x"c0",x"1e"),
   763 => (x"26",x"86",x"cc",x"87"),
   764 => (x"00",x"00",x"00",x"4f"),
   765 => (x"00",x"00",x"00",x"00"),
   766 => (x"00",x"00",x"61",x"a8"),
   767 => (x"67",x"6f",x"72",x"50"),
   768 => (x"20",x"6d",x"61",x"72"),
   769 => (x"70",x"6d",x"6f",x"63"),
   770 => (x"64",x"65",x"6c",x"69"),
   771 => (x"74",x"69",x"77",x"20"),
   772 => (x"72",x"27",x"20",x"68"),
   773 => (x"73",x"69",x"67",x"65"),
   774 => (x"27",x"72",x"65",x"74"),
   775 => (x"74",x"74",x"61",x"20"),
   776 => (x"75",x"62",x"69",x"72"),
   777 => (x"00",x"0a",x"65",x"74"),
   778 => (x"00",x"00",x"00",x"0a"),
   779 => (x"67",x"6f",x"72",x"50"),
   780 => (x"20",x"6d",x"61",x"72"),
   781 => (x"70",x"6d",x"6f",x"63"),
   782 => (x"64",x"65",x"6c",x"69"),
   783 => (x"74",x"69",x"77",x"20"),
   784 => (x"74",x"75",x"6f",x"68"),
   785 => (x"65",x"72",x"27",x"20"),
   786 => (x"74",x"73",x"69",x"67"),
   787 => (x"20",x"27",x"72",x"65"),
   788 => (x"72",x"74",x"74",x"61"),
   789 => (x"74",x"75",x"62",x"69"),
   790 => (x"00",x"00",x"0a",x"65"),
   791 => (x"00",x"00",x"00",x"0a"),
   792 => (x"59",x"52",x"48",x"44"),
   793 => (x"4e",x"4f",x"54",x"53"),
   794 => (x"52",x"50",x"20",x"45"),
   795 => (x"41",x"52",x"47",x"4f"),
   796 => (x"33",x"20",x"2c",x"4d"),
   797 => (x"20",x"44",x"52",x"27"),
   798 => (x"49",x"52",x"54",x"53"),
   799 => (x"00",x"00",x"47",x"4e"),
   800 => (x"59",x"52",x"48",x"44"),
   801 => (x"4e",x"4f",x"54",x"53"),
   802 => (x"52",x"50",x"20",x"45"),
   803 => (x"41",x"52",x"47",x"4f"),
   804 => (x"32",x"20",x"2c",x"4d"),
   805 => (x"20",x"44",x"4e",x"27"),
   806 => (x"49",x"52",x"54",x"53"),
   807 => (x"00",x"00",x"47",x"4e"),
   808 => (x"73",x"61",x"65",x"4d"),
   809 => (x"64",x"65",x"72",x"75"),
   810 => (x"6d",x"69",x"74",x"20"),
   811 => (x"6f",x"74",x"20",x"65"),
   812 => (x"6d",x"73",x"20",x"6f"),
   813 => (x"20",x"6c",x"6c",x"61"),
   814 => (x"6f",x"20",x"6f",x"74"),
   815 => (x"69",x"61",x"74",x"62"),
   816 => (x"65",x"6d",x"20",x"6e"),
   817 => (x"6e",x"69",x"6e",x"61"),
   818 => (x"6c",x"75",x"66",x"67"),
   819 => (x"73",x"65",x"72",x"20"),
   820 => (x"73",x"74",x"6c",x"75"),
   821 => (x"00",x"00",x"00",x"0a"),
   822 => (x"61",x"65",x"6c",x"50"),
   823 => (x"69",x"20",x"65",x"73"),
   824 => (x"65",x"72",x"63",x"6e"),
   825 => (x"20",x"65",x"73",x"61"),
   826 => (x"62",x"6d",x"75",x"6e"),
   827 => (x"6f",x"20",x"72",x"65"),
   828 => (x"75",x"72",x"20",x"66"),
   829 => (x"00",x"0a",x"73",x"6e"),
   830 => (x"00",x"00",x"00",x"0a"),
   831 => (x"72",x"63",x"69",x"4d"),
   832 => (x"63",x"65",x"73",x"6f"),
   833 => (x"73",x"64",x"6e",x"6f"),
   834 => (x"72",x"6f",x"66",x"20"),
   835 => (x"65",x"6e",x"6f",x"20"),
   836 => (x"6e",x"75",x"72",x"20"),
   837 => (x"72",x"68",x"74",x"20"),
   838 => (x"68",x"67",x"75",x"6f"),
   839 => (x"72",x"68",x"44",x"20"),
   840 => (x"6f",x"74",x"73",x"79"),
   841 => (x"20",x"3a",x"65",x"6e"),
   842 => (x"00",x"00",x"00",x"00"),
   843 => (x"0a",x"20",x"64",x"25"),
   844 => (x"00",x"00",x"00",x"00"),
   845 => (x"79",x"72",x"68",x"44"),
   846 => (x"6e",x"6f",x"74",x"73"),
   847 => (x"70",x"20",x"73",x"65"),
   848 => (x"53",x"20",x"72",x"65"),
   849 => (x"6e",x"6f",x"63",x"65"),
   850 => (x"20",x"20",x"3a",x"64"),
   851 => (x"20",x"20",x"20",x"20"),
   852 => (x"20",x"20",x"20",x"20"),
   853 => (x"20",x"20",x"20",x"20"),
   854 => (x"20",x"20",x"20",x"20"),
   855 => (x"20",x"20",x"20",x"20"),
   856 => (x"00",x"00",x"00",x"00"),
   857 => (x"0a",x"20",x"64",x"25"),
   858 => (x"00",x"00",x"00",x"00"),
   859 => (x"20",x"58",x"41",x"56"),
   860 => (x"53",x"50",x"49",x"4d"),
   861 => (x"74",x"61",x"72",x"20"),
   862 => (x"20",x"67",x"6e",x"69"),
   863 => (x"30",x"31",x"20",x"2a"),
   864 => (x"3d",x"20",x"30",x"30"),
   865 => (x"20",x"64",x"25",x"20"),
   866 => (x"00",x"00",x"00",x"0a"),
   867 => (x"00",x"00",x"00",x"0a"),
   868 => (x"59",x"52",x"48",x"44"),
   869 => (x"4e",x"4f",x"54",x"53"),
   870 => (x"52",x"50",x"20",x"45"),
   871 => (x"41",x"52",x"47",x"4f"),
   872 => (x"53",x"20",x"2c",x"4d"),
   873 => (x"20",x"45",x"4d",x"4f"),
   874 => (x"49",x"52",x"54",x"53"),
   875 => (x"00",x"00",x"47",x"4e"),
   876 => (x"59",x"52",x"48",x"44"),
   877 => (x"4e",x"4f",x"54",x"53"),
   878 => (x"52",x"50",x"20",x"45"),
   879 => (x"41",x"52",x"47",x"4f"),
   880 => (x"31",x"20",x"2c",x"4d"),
   881 => (x"20",x"54",x"53",x"27"),
   882 => (x"49",x"52",x"54",x"53"),
   883 => (x"00",x"00",x"47",x"4e"),
   884 => (x"00",x"00",x"00",x"0a"),
   885 => (x"79",x"72",x"68",x"44"),
   886 => (x"6e",x"6f",x"74",x"73"),
   887 => (x"65",x"42",x"20",x"65"),
   888 => (x"6d",x"68",x"63",x"6e"),
   889 => (x"2c",x"6b",x"72",x"61"),
   890 => (x"72",x"65",x"56",x"20"),
   891 => (x"6e",x"6f",x"69",x"73"),
   892 => (x"31",x"2e",x"32",x"20"),
   893 => (x"61",x"4c",x"28",x"20"),
   894 => (x"61",x"75",x"67",x"6e"),
   895 => (x"20",x"3a",x"65",x"67"),
   896 => (x"00",x"0a",x"29",x"43"),
   897 => (x"00",x"00",x"00",x"0a"),
   898 => (x"63",x"65",x"78",x"45"),
   899 => (x"6f",x"69",x"74",x"75"),
   900 => (x"74",x"73",x"20",x"6e"),
   901 => (x"73",x"74",x"72",x"61"),
   902 => (x"64",x"25",x"20",x"2c"),
   903 => (x"6e",x"75",x"72",x"20"),
   904 => (x"68",x"74",x"20",x"73"),
   905 => (x"67",x"75",x"6f",x"72"),
   906 => (x"68",x"44",x"20",x"68"),
   907 => (x"74",x"73",x"79",x"72"),
   908 => (x"0a",x"65",x"6e",x"6f"),
   909 => (x"00",x"00",x"00",x"00"),
   910 => (x"63",x"65",x"78",x"45"),
   911 => (x"6f",x"69",x"74",x"75"),
   912 => (x"6e",x"65",x"20",x"6e"),
   913 => (x"00",x"0a",x"73",x"64"),
   914 => (x"00",x"00",x"00",x"0a"),
   915 => (x"61",x"6e",x"69",x"46"),
   916 => (x"61",x"76",x"20",x"6c"),
   917 => (x"73",x"65",x"75",x"6c"),
   918 => (x"20",x"66",x"6f",x"20"),
   919 => (x"20",x"65",x"68",x"74"),
   920 => (x"69",x"72",x"61",x"76"),
   921 => (x"65",x"6c",x"62",x"61"),
   922 => (x"73",x"75",x"20",x"73"),
   923 => (x"69",x"20",x"64",x"65"),
   924 => (x"68",x"74",x"20",x"6e"),
   925 => (x"65",x"62",x"20",x"65"),
   926 => (x"6d",x"68",x"63",x"6e"),
   927 => (x"3a",x"6b",x"72",x"61"),
   928 => (x"00",x"00",x"00",x"0a"),
   929 => (x"00",x"00",x"00",x"0a"),
   930 => (x"5f",x"74",x"6e",x"49"),
   931 => (x"62",x"6f",x"6c",x"47"),
   932 => (x"20",x"20",x"20",x"3a"),
   933 => (x"20",x"20",x"20",x"20"),
   934 => (x"20",x"20",x"20",x"20"),
   935 => (x"0a",x"64",x"25",x"20"),
   936 => (x"00",x"00",x"00",x"00"),
   937 => (x"20",x"20",x"20",x"20"),
   938 => (x"20",x"20",x"20",x"20"),
   939 => (x"75",x"6f",x"68",x"73"),
   940 => (x"62",x"20",x"64",x"6c"),
   941 => (x"20",x"20",x"3a",x"65"),
   942 => (x"0a",x"64",x"25",x"20"),
   943 => (x"00",x"00",x"00",x"00"),
   944 => (x"6c",x"6f",x"6f",x"42"),
   945 => (x"6f",x"6c",x"47",x"5f"),
   946 => (x"20",x"20",x"3a",x"62"),
   947 => (x"20",x"20",x"20",x"20"),
   948 => (x"20",x"20",x"20",x"20"),
   949 => (x"0a",x"64",x"25",x"20"),
   950 => (x"00",x"00",x"00",x"00"),
   951 => (x"20",x"20",x"20",x"20"),
   952 => (x"20",x"20",x"20",x"20"),
   953 => (x"75",x"6f",x"68",x"73"),
   954 => (x"62",x"20",x"64",x"6c"),
   955 => (x"20",x"20",x"3a",x"65"),
   956 => (x"0a",x"64",x"25",x"20"),
   957 => (x"00",x"00",x"00",x"00"),
   958 => (x"31",x"5f",x"68",x"43"),
   959 => (x"6f",x"6c",x"47",x"5f"),
   960 => (x"20",x"20",x"3a",x"62"),
   961 => (x"20",x"20",x"20",x"20"),
   962 => (x"20",x"20",x"20",x"20"),
   963 => (x"0a",x"63",x"25",x"20"),
   964 => (x"00",x"00",x"00",x"00"),
   965 => (x"20",x"20",x"20",x"20"),
   966 => (x"20",x"20",x"20",x"20"),
   967 => (x"75",x"6f",x"68",x"73"),
   968 => (x"62",x"20",x"64",x"6c"),
   969 => (x"20",x"20",x"3a",x"65"),
   970 => (x"0a",x"63",x"25",x"20"),
   971 => (x"00",x"00",x"00",x"00"),
   972 => (x"32",x"5f",x"68",x"43"),
   973 => (x"6f",x"6c",x"47",x"5f"),
   974 => (x"20",x"20",x"3a",x"62"),
   975 => (x"20",x"20",x"20",x"20"),
   976 => (x"20",x"20",x"20",x"20"),
   977 => (x"0a",x"63",x"25",x"20"),
   978 => (x"00",x"00",x"00",x"00"),
   979 => (x"20",x"20",x"20",x"20"),
   980 => (x"20",x"20",x"20",x"20"),
   981 => (x"75",x"6f",x"68",x"73"),
   982 => (x"62",x"20",x"64",x"6c"),
   983 => (x"20",x"20",x"3a",x"65"),
   984 => (x"0a",x"63",x"25",x"20"),
   985 => (x"00",x"00",x"00",x"00"),
   986 => (x"5f",x"72",x"72",x"41"),
   987 => (x"6c",x"47",x"5f",x"31"),
   988 => (x"38",x"5b",x"62",x"6f"),
   989 => (x"20",x"20",x"3a",x"5d"),
   990 => (x"20",x"20",x"20",x"20"),
   991 => (x"0a",x"64",x"25",x"20"),
   992 => (x"00",x"00",x"00",x"00"),
   993 => (x"20",x"20",x"20",x"20"),
   994 => (x"20",x"20",x"20",x"20"),
   995 => (x"75",x"6f",x"68",x"73"),
   996 => (x"62",x"20",x"64",x"6c"),
   997 => (x"20",x"20",x"3a",x"65"),
   998 => (x"0a",x"64",x"25",x"20"),
   999 => (x"00",x"00",x"00",x"00"),
  1000 => (x"5f",x"72",x"72",x"41"),
  1001 => (x"6c",x"47",x"5f",x"32"),
  1002 => (x"38",x"5b",x"62",x"6f"),
  1003 => (x"5d",x"37",x"5b",x"5d"),
  1004 => (x"20",x"20",x"20",x"3a"),
  1005 => (x"0a",x"64",x"25",x"20"),
  1006 => (x"00",x"00",x"00",x"00"),
  1007 => (x"20",x"20",x"20",x"20"),
  1008 => (x"20",x"20",x"20",x"20"),
  1009 => (x"75",x"6f",x"68",x"73"),
  1010 => (x"62",x"20",x"64",x"6c"),
  1011 => (x"20",x"20",x"3a",x"65"),
  1012 => (x"6d",x"75",x"4e",x"20"),
  1013 => (x"5f",x"72",x"65",x"62"),
  1014 => (x"52",x"5f",x"66",x"4f"),
  1015 => (x"20",x"73",x"6e",x"75"),
  1016 => (x"30",x"31",x"20",x"2b"),
  1017 => (x"00",x"00",x"00",x"0a"),
  1018 => (x"5f",x"72",x"74",x"50"),
  1019 => (x"62",x"6f",x"6c",x"47"),
  1020 => (x"00",x"0a",x"3e",x"2d"),
  1021 => (x"74",x"50",x"20",x"20"),
  1022 => (x"6f",x"43",x"5f",x"72"),
  1023 => (x"20",x"3a",x"70",x"6d"),
  1024 => (x"20",x"20",x"20",x"20"),
  1025 => (x"20",x"20",x"20",x"20"),
  1026 => (x"0a",x"64",x"25",x"20"),
  1027 => (x"00",x"00",x"00",x"00"),
  1028 => (x"20",x"20",x"20",x"20"),
  1029 => (x"20",x"20",x"20",x"20"),
  1030 => (x"75",x"6f",x"68",x"73"),
  1031 => (x"62",x"20",x"64",x"6c"),
  1032 => (x"20",x"20",x"3a",x"65"),
  1033 => (x"6d",x"69",x"28",x"20"),
  1034 => (x"6d",x"65",x"6c",x"70"),
  1035 => (x"61",x"74",x"6e",x"65"),
  1036 => (x"6e",x"6f",x"69",x"74"),
  1037 => (x"70",x"65",x"64",x"2d"),
  1038 => (x"65",x"64",x"6e",x"65"),
  1039 => (x"0a",x"29",x"74",x"6e"),
  1040 => (x"00",x"00",x"00",x"00"),
  1041 => (x"69",x"44",x"20",x"20"),
  1042 => (x"3a",x"72",x"63",x"73"),
  1043 => (x"20",x"20",x"20",x"20"),
  1044 => (x"20",x"20",x"20",x"20"),
  1045 => (x"20",x"20",x"20",x"20"),
  1046 => (x"0a",x"64",x"25",x"20"),
  1047 => (x"00",x"00",x"00",x"00"),
  1048 => (x"20",x"20",x"20",x"20"),
  1049 => (x"20",x"20",x"20",x"20"),
  1050 => (x"75",x"6f",x"68",x"73"),
  1051 => (x"62",x"20",x"64",x"6c"),
  1052 => (x"20",x"20",x"3a",x"65"),
  1053 => (x"0a",x"64",x"25",x"20"),
  1054 => (x"00",x"00",x"00",x"00"),
  1055 => (x"6e",x"45",x"20",x"20"),
  1056 => (x"43",x"5f",x"6d",x"75"),
  1057 => (x"3a",x"70",x"6d",x"6f"),
  1058 => (x"20",x"20",x"20",x"20"),
  1059 => (x"20",x"20",x"20",x"20"),
  1060 => (x"0a",x"64",x"25",x"20"),
  1061 => (x"00",x"00",x"00",x"00"),
  1062 => (x"20",x"20",x"20",x"20"),
  1063 => (x"20",x"20",x"20",x"20"),
  1064 => (x"75",x"6f",x"68",x"73"),
  1065 => (x"62",x"20",x"64",x"6c"),
  1066 => (x"20",x"20",x"3a",x"65"),
  1067 => (x"0a",x"64",x"25",x"20"),
  1068 => (x"00",x"00",x"00",x"00"),
  1069 => (x"6e",x"49",x"20",x"20"),
  1070 => (x"6f",x"43",x"5f",x"74"),
  1071 => (x"20",x"3a",x"70",x"6d"),
  1072 => (x"20",x"20",x"20",x"20"),
  1073 => (x"20",x"20",x"20",x"20"),
  1074 => (x"0a",x"64",x"25",x"20"),
  1075 => (x"00",x"00",x"00",x"00"),
  1076 => (x"20",x"20",x"20",x"20"),
  1077 => (x"20",x"20",x"20",x"20"),
  1078 => (x"75",x"6f",x"68",x"73"),
  1079 => (x"62",x"20",x"64",x"6c"),
  1080 => (x"20",x"20",x"3a",x"65"),
  1081 => (x"0a",x"64",x"25",x"20"),
  1082 => (x"00",x"00",x"00",x"00"),
  1083 => (x"74",x"53",x"20",x"20"),
  1084 => (x"6f",x"43",x"5f",x"72"),
  1085 => (x"20",x"3a",x"70",x"6d"),
  1086 => (x"20",x"20",x"20",x"20"),
  1087 => (x"20",x"20",x"20",x"20"),
  1088 => (x"0a",x"73",x"25",x"20"),
  1089 => (x"00",x"00",x"00",x"00"),
  1090 => (x"20",x"20",x"20",x"20"),
  1091 => (x"20",x"20",x"20",x"20"),
  1092 => (x"75",x"6f",x"68",x"73"),
  1093 => (x"62",x"20",x"64",x"6c"),
  1094 => (x"20",x"20",x"3a",x"65"),
  1095 => (x"52",x"48",x"44",x"20"),
  1096 => (x"4f",x"54",x"53",x"59"),
  1097 => (x"50",x"20",x"45",x"4e"),
  1098 => (x"52",x"47",x"4f",x"52"),
  1099 => (x"20",x"2c",x"4d",x"41"),
  1100 => (x"45",x"4d",x"4f",x"53"),
  1101 => (x"52",x"54",x"53",x"20"),
  1102 => (x"0a",x"47",x"4e",x"49"),
  1103 => (x"00",x"00",x"00",x"00"),
  1104 => (x"74",x"78",x"65",x"4e"),
  1105 => (x"72",x"74",x"50",x"5f"),
  1106 => (x"6f",x"6c",x"47",x"5f"),
  1107 => (x"0a",x"3e",x"2d",x"62"),
  1108 => (x"00",x"00",x"00",x"00"),
  1109 => (x"74",x"50",x"20",x"20"),
  1110 => (x"6f",x"43",x"5f",x"72"),
  1111 => (x"20",x"3a",x"70",x"6d"),
  1112 => (x"20",x"20",x"20",x"20"),
  1113 => (x"20",x"20",x"20",x"20"),
  1114 => (x"0a",x"64",x"25",x"20"),
  1115 => (x"00",x"00",x"00",x"00"),
  1116 => (x"20",x"20",x"20",x"20"),
  1117 => (x"20",x"20",x"20",x"20"),
  1118 => (x"75",x"6f",x"68",x"73"),
  1119 => (x"62",x"20",x"64",x"6c"),
  1120 => (x"20",x"20",x"3a",x"65"),
  1121 => (x"6d",x"69",x"28",x"20"),
  1122 => (x"6d",x"65",x"6c",x"70"),
  1123 => (x"61",x"74",x"6e",x"65"),
  1124 => (x"6e",x"6f",x"69",x"74"),
  1125 => (x"70",x"65",x"64",x"2d"),
  1126 => (x"65",x"64",x"6e",x"65"),
  1127 => (x"2c",x"29",x"74",x"6e"),
  1128 => (x"6d",x"61",x"73",x"20"),
  1129 => (x"73",x"61",x"20",x"65"),
  1130 => (x"6f",x"62",x"61",x"20"),
  1131 => (x"00",x"0a",x"65",x"76"),
  1132 => (x"69",x"44",x"20",x"20"),
  1133 => (x"3a",x"72",x"63",x"73"),
  1134 => (x"20",x"20",x"20",x"20"),
  1135 => (x"20",x"20",x"20",x"20"),
  1136 => (x"20",x"20",x"20",x"20"),
  1137 => (x"0a",x"64",x"25",x"20"),
  1138 => (x"00",x"00",x"00",x"00"),
  1139 => (x"20",x"20",x"20",x"20"),
  1140 => (x"20",x"20",x"20",x"20"),
  1141 => (x"75",x"6f",x"68",x"73"),
  1142 => (x"62",x"20",x"64",x"6c"),
  1143 => (x"20",x"20",x"3a",x"65"),
  1144 => (x"0a",x"64",x"25",x"20"),
  1145 => (x"00",x"00",x"00",x"00"),
  1146 => (x"6e",x"45",x"20",x"20"),
  1147 => (x"43",x"5f",x"6d",x"75"),
  1148 => (x"3a",x"70",x"6d",x"6f"),
  1149 => (x"20",x"20",x"20",x"20"),
  1150 => (x"20",x"20",x"20",x"20"),
  1151 => (x"0a",x"64",x"25",x"20"),
  1152 => (x"00",x"00",x"00",x"00"),
  1153 => (x"20",x"20",x"20",x"20"),
  1154 => (x"20",x"20",x"20",x"20"),
  1155 => (x"75",x"6f",x"68",x"73"),
  1156 => (x"62",x"20",x"64",x"6c"),
  1157 => (x"20",x"20",x"3a",x"65"),
  1158 => (x"0a",x"64",x"25",x"20"),
  1159 => (x"00",x"00",x"00",x"00"),
  1160 => (x"6e",x"49",x"20",x"20"),
  1161 => (x"6f",x"43",x"5f",x"74"),
  1162 => (x"20",x"3a",x"70",x"6d"),
  1163 => (x"20",x"20",x"20",x"20"),
  1164 => (x"20",x"20",x"20",x"20"),
  1165 => (x"0a",x"64",x"25",x"20"),
  1166 => (x"00",x"00",x"00",x"00"),
  1167 => (x"20",x"20",x"20",x"20"),
  1168 => (x"20",x"20",x"20",x"20"),
  1169 => (x"75",x"6f",x"68",x"73"),
  1170 => (x"62",x"20",x"64",x"6c"),
  1171 => (x"20",x"20",x"3a",x"65"),
  1172 => (x"0a",x"64",x"25",x"20"),
  1173 => (x"00",x"00",x"00",x"00"),
  1174 => (x"74",x"53",x"20",x"20"),
  1175 => (x"6f",x"43",x"5f",x"72"),
  1176 => (x"20",x"3a",x"70",x"6d"),
  1177 => (x"20",x"20",x"20",x"20"),
  1178 => (x"20",x"20",x"20",x"20"),
  1179 => (x"0a",x"73",x"25",x"20"),
  1180 => (x"00",x"00",x"00",x"00"),
  1181 => (x"20",x"20",x"20",x"20"),
  1182 => (x"20",x"20",x"20",x"20"),
  1183 => (x"75",x"6f",x"68",x"73"),
  1184 => (x"62",x"20",x"64",x"6c"),
  1185 => (x"20",x"20",x"3a",x"65"),
  1186 => (x"52",x"48",x"44",x"20"),
  1187 => (x"4f",x"54",x"53",x"59"),
  1188 => (x"50",x"20",x"45",x"4e"),
  1189 => (x"52",x"47",x"4f",x"52"),
  1190 => (x"20",x"2c",x"4d",x"41"),
  1191 => (x"45",x"4d",x"4f",x"53"),
  1192 => (x"52",x"54",x"53",x"20"),
  1193 => (x"0a",x"47",x"4e",x"49"),
  1194 => (x"00",x"00",x"00",x"00"),
  1195 => (x"5f",x"74",x"6e",x"49"),
  1196 => (x"6f",x"4c",x"5f",x"31"),
  1197 => (x"20",x"20",x"3a",x"63"),
  1198 => (x"20",x"20",x"20",x"20"),
  1199 => (x"20",x"20",x"20",x"20"),
  1200 => (x"0a",x"64",x"25",x"20"),
  1201 => (x"00",x"00",x"00",x"00"),
  1202 => (x"20",x"20",x"20",x"20"),
  1203 => (x"20",x"20",x"20",x"20"),
  1204 => (x"75",x"6f",x"68",x"73"),
  1205 => (x"62",x"20",x"64",x"6c"),
  1206 => (x"20",x"20",x"3a",x"65"),
  1207 => (x"0a",x"64",x"25",x"20"),
  1208 => (x"00",x"00",x"00",x"00"),
  1209 => (x"5f",x"74",x"6e",x"49"),
  1210 => (x"6f",x"4c",x"5f",x"32"),
  1211 => (x"20",x"20",x"3a",x"63"),
  1212 => (x"20",x"20",x"20",x"20"),
  1213 => (x"20",x"20",x"20",x"20"),
  1214 => (x"0a",x"64",x"25",x"20"),
  1215 => (x"00",x"00",x"00",x"00"),
  1216 => (x"20",x"20",x"20",x"20"),
  1217 => (x"20",x"20",x"20",x"20"),
  1218 => (x"75",x"6f",x"68",x"73"),
  1219 => (x"62",x"20",x"64",x"6c"),
  1220 => (x"20",x"20",x"3a",x"65"),
  1221 => (x"0a",x"64",x"25",x"20"),
  1222 => (x"00",x"00",x"00",x"00"),
  1223 => (x"5f",x"74",x"6e",x"49"),
  1224 => (x"6f",x"4c",x"5f",x"33"),
  1225 => (x"20",x"20",x"3a",x"63"),
  1226 => (x"20",x"20",x"20",x"20"),
  1227 => (x"20",x"20",x"20",x"20"),
  1228 => (x"0a",x"64",x"25",x"20"),
  1229 => (x"00",x"00",x"00",x"00"),
  1230 => (x"20",x"20",x"20",x"20"),
  1231 => (x"20",x"20",x"20",x"20"),
  1232 => (x"75",x"6f",x"68",x"73"),
  1233 => (x"62",x"20",x"64",x"6c"),
  1234 => (x"20",x"20",x"3a",x"65"),
  1235 => (x"0a",x"64",x"25",x"20"),
  1236 => (x"00",x"00",x"00",x"00"),
  1237 => (x"6d",x"75",x"6e",x"45"),
  1238 => (x"63",x"6f",x"4c",x"5f"),
  1239 => (x"20",x"20",x"20",x"3a"),
  1240 => (x"20",x"20",x"20",x"20"),
  1241 => (x"20",x"20",x"20",x"20"),
  1242 => (x"0a",x"64",x"25",x"20"),
  1243 => (x"00",x"00",x"00",x"00"),
  1244 => (x"20",x"20",x"20",x"20"),
  1245 => (x"20",x"20",x"20",x"20"),
  1246 => (x"75",x"6f",x"68",x"73"),
  1247 => (x"62",x"20",x"64",x"6c"),
  1248 => (x"20",x"20",x"3a",x"65"),
  1249 => (x"0a",x"64",x"25",x"20"),
  1250 => (x"00",x"00",x"00",x"00"),
  1251 => (x"5f",x"72",x"74",x"53"),
  1252 => (x"6f",x"4c",x"5f",x"31"),
  1253 => (x"20",x"20",x"3a",x"63"),
  1254 => (x"20",x"20",x"20",x"20"),
  1255 => (x"20",x"20",x"20",x"20"),
  1256 => (x"0a",x"73",x"25",x"20"),
  1257 => (x"00",x"00",x"00",x"00"),
  1258 => (x"20",x"20",x"20",x"20"),
  1259 => (x"20",x"20",x"20",x"20"),
  1260 => (x"75",x"6f",x"68",x"73"),
  1261 => (x"62",x"20",x"64",x"6c"),
  1262 => (x"20",x"20",x"3a",x"65"),
  1263 => (x"52",x"48",x"44",x"20"),
  1264 => (x"4f",x"54",x"53",x"59"),
  1265 => (x"50",x"20",x"45",x"4e"),
  1266 => (x"52",x"47",x"4f",x"52"),
  1267 => (x"20",x"2c",x"4d",x"41"),
  1268 => (x"54",x"53",x"27",x"31"),
  1269 => (x"52",x"54",x"53",x"20"),
  1270 => (x"0a",x"47",x"4e",x"49"),
  1271 => (x"00",x"00",x"00",x"00"),
  1272 => (x"5f",x"72",x"74",x"53"),
  1273 => (x"6f",x"4c",x"5f",x"32"),
  1274 => (x"20",x"20",x"3a",x"63"),
  1275 => (x"20",x"20",x"20",x"20"),
  1276 => (x"20",x"20",x"20",x"20"),
  1277 => (x"0a",x"73",x"25",x"20"),
  1278 => (x"00",x"00",x"00",x"00"),
  1279 => (x"20",x"20",x"20",x"20"),
  1280 => (x"20",x"20",x"20",x"20"),
  1281 => (x"75",x"6f",x"68",x"73"),
  1282 => (x"62",x"20",x"64",x"6c"),
  1283 => (x"20",x"20",x"3a",x"65"),
  1284 => (x"52",x"48",x"44",x"20"),
  1285 => (x"4f",x"54",x"53",x"59"),
  1286 => (x"50",x"20",x"45",x"4e"),
  1287 => (x"52",x"47",x"4f",x"52"),
  1288 => (x"20",x"2c",x"4d",x"41"),
  1289 => (x"44",x"4e",x"27",x"32"),
  1290 => (x"52",x"54",x"53",x"20"),
  1291 => (x"0a",x"47",x"4e",x"49"),
  1292 => (x"00",x"00",x"00",x"00"),
  1293 => (x"00",x"00",x"00",x"0a"),
  1294 => (x"72",x"65",x"73",x"55"),
  1295 => (x"6d",x"69",x"74",x"20"),
  1296 => (x"25",x"20",x"3a",x"65"),
  1297 => (x"0e",x"00",x"0a",x"64"),
  1298 => (x"c8",x"0e",x"5b",x"5e"),
  1299 => (x"66",x"cc",x"4b",x"66"),
  1300 => (x"c2",x"79",x"73",x"49"),
  1301 => (x"87",x"c4",x"05",x"ab"),
  1302 => (x"87",x"c2",x"4a",x"c1"),
  1303 => (x"9a",x"72",x"4a",x"c0"),
  1304 => (x"c3",x"87",x"c2",x"05"),
  1305 => (x"02",x"ab",x"c0",x"79"),
  1306 => (x"ab",x"c1",x"87",x"d8"),
  1307 => (x"c2",x"87",x"d7",x"02"),
  1308 => (x"e5",x"c0",x"02",x"ab"),
  1309 => (x"02",x"ab",x"c3",x"87"),
  1310 => (x"c4",x"87",x"e5",x"c0"),
  1311 => (x"87",x"de",x"02",x"ab"),
  1312 => (x"79",x"c0",x"87",x"de"),
  1313 => (x"d8",x"c1",x"87",x"da"),
  1314 => (x"c1",x"48",x"bf",x"fc"),
  1315 => (x"06",x"a8",x"b7",x"e4"),
  1316 => (x"79",x"c0",x"87",x"c4"),
  1317 => (x"79",x"c3",x"87",x"ca"),
  1318 => (x"79",x"c1",x"87",x"c6"),
  1319 => (x"79",x"c2",x"87",x"c2"),
  1320 => (x"4f",x"26",x"4b",x"26"),
  1321 => (x"48",x"66",x"c4",x"1e"),
  1322 => (x"c4",x"05",x"a8",x"c2"),
  1323 => (x"c2",x"48",x"c1",x"87"),
  1324 => (x"26",x"48",x"c0",x"87"),
  1325 => (x"66",x"c4",x"1e",x"4f"),
  1326 => (x"c8",x"81",x"c2",x"49"),
  1327 => (x"80",x"71",x"48",x"66"),
  1328 => (x"78",x"08",x"66",x"cc"),
  1329 => (x"0e",x"4f",x"26",x"08"),
  1330 => (x"5d",x"5c",x"5b",x"5e"),
  1331 => (x"c0",x"86",x"f4",x"0e"),
  1332 => (x"c5",x"4c",x"66",x"e4"),
  1333 => (x"c4",x"48",x"74",x"84"),
  1334 => (x"a6",x"c8",x"90",x"b7"),
  1335 => (x"48",x"66",x"dc",x"58"),
  1336 => (x"c4",x"80",x"66",x"c4"),
  1337 => (x"48",x"6e",x"58",x"a6"),
  1338 => (x"78",x"66",x"e8",x"c0"),
  1339 => (x"80",x"c1",x"48",x"74"),
  1340 => (x"c8",x"58",x"a6",x"cc"),
  1341 => (x"b7",x"c4",x"49",x"66"),
  1342 => (x"81",x"66",x"dc",x"91"),
  1343 => (x"79",x"66",x"e8",x"c0"),
  1344 => (x"81",x"de",x"49",x"74"),
  1345 => (x"dc",x"91",x"b7",x"c4"),
  1346 => (x"79",x"74",x"81",x"66"),
  1347 => (x"ac",x"b7",x"66",x"c8"),
  1348 => (x"87",x"e3",x"c0",x"01"),
  1349 => (x"c8",x"c3",x"49",x"74"),
  1350 => (x"e0",x"c0",x"91",x"b7"),
  1351 => (x"4d",x"c4",x"81",x"66"),
  1352 => (x"66",x"c4",x"4a",x"71"),
  1353 => (x"4b",x"66",x"c8",x"82"),
  1354 => (x"83",x"c1",x"8b",x"74"),
  1355 => (x"82",x"75",x"7a",x"74"),
  1356 => (x"9b",x"73",x"8b",x"c1"),
  1357 => (x"74",x"87",x"f5",x"01"),
  1358 => (x"b7",x"c8",x"c3",x"4a"),
  1359 => (x"66",x"e0",x"c0",x"92"),
  1360 => (x"c1",x"49",x"74",x"82"),
  1361 => (x"91",x"b7",x"c4",x"89"),
  1362 => (x"48",x"69",x"81",x"72"),
  1363 => (x"79",x"70",x"80",x"c1"),
  1364 => (x"81",x"d4",x"49",x"74"),
  1365 => (x"91",x"b7",x"c8",x"c3"),
  1366 => (x"81",x"66",x"e0",x"c0"),
  1367 => (x"6e",x"81",x"66",x"c4"),
  1368 => (x"d8",x"c1",x"79",x"bf"),
  1369 => (x"78",x"c5",x"48",x"fc"),
  1370 => (x"4d",x"26",x"8e",x"f4"),
  1371 => (x"4b",x"26",x"4c",x"26"),
  1372 => (x"5e",x"0e",x"4f",x"26"),
  1373 => (x"c8",x"97",x"0e",x"5b"),
  1374 => (x"4a",x"73",x"4b",x"66"),
  1375 => (x"ba",x"82",x"c0",x"fe"),
  1376 => (x"49",x"66",x"cc",x"97"),
  1377 => (x"b9",x"81",x"c0",x"fe"),
  1378 => (x"02",x"aa",x"b7",x"71"),
  1379 => (x"48",x"c0",x"87",x"c4"),
  1380 => (x"d9",x"c1",x"87",x"c7"),
  1381 => (x"c1",x"5b",x"97",x"c8"),
  1382 => (x"26",x"4b",x"26",x"48"),
  1383 => (x"5b",x"5e",x"0e",x"4f"),
  1384 => (x"f8",x"0e",x"5d",x"5c"),
  1385 => (x"dc",x"4d",x"c2",x"86"),
  1386 => (x"81",x"c1",x"49",x"66"),
  1387 => (x"c2",x"4c",x"66",x"d8"),
  1388 => (x"c2",x"4b",x"71",x"84"),
  1389 => (x"fe",x"49",x"13",x"83"),
  1390 => (x"c3",x"b9",x"81",x"c0"),
  1391 => (x"4a",x"14",x"99",x"ff"),
  1392 => (x"ba",x"82",x"c0",x"fe"),
  1393 => (x"5a",x"97",x"a6",x"c4"),
  1394 => (x"fe",x"4a",x"6e",x"97"),
  1395 => (x"fe",x"ba",x"82",x"c0"),
  1396 => (x"71",x"b9",x"81",x"c0"),
  1397 => (x"c7",x"02",x"aa",x"b7"),
  1398 => (x"48",x"a6",x"c4",x"87"),
  1399 => (x"87",x"cc",x"78",x"c0"),
  1400 => (x"48",x"c4",x"d9",x"c1"),
  1401 => (x"c4",x"50",x"6e",x"97"),
  1402 => (x"78",x"c1",x"48",x"a6"),
  1403 => (x"c2",x"05",x"66",x"c4"),
  1404 => (x"c2",x"85",x"c1",x"87"),
  1405 => (x"fe",x"06",x"ad",x"b7"),
  1406 => (x"66",x"d8",x"87",x"fb"),
  1407 => (x"49",x"66",x"dc",x"4a"),
  1408 => (x"87",x"ee",x"f7",x"fe"),
  1409 => (x"06",x"a8",x"b7",x"c0"),
  1410 => (x"48",x"75",x"87",x"cc"),
  1411 => (x"d9",x"c1",x"80",x"c7"),
  1412 => (x"48",x"c1",x"58",x"c0"),
  1413 => (x"48",x"c0",x"87",x"c2"),
  1414 => (x"4d",x"26",x"8e",x"f8"),
  1415 => (x"4b",x"26",x"4c",x"26"),
  1416 => (x"4b",x"26",x"4f",x"26"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
