
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"d7",x"01"),
     1 => (x"58",x"0e",x"87",x"da"),
     2 => (x"27",x"0e",x"59",x"5e"),
     3 => (x"00",x"00",x"00",x"43"),
     4 => (x"26",x"49",x"26",x"0f"),
     5 => (x"26",x"80",x"ff",x"48"),
     6 => (x"26",x"27",x"4f",x"08"),
     7 => (x"4f",x"00",x"00",x"00"),
     8 => (x"00",x"00",x"35",x"27"),
     9 => (x"b8",x"27",x"4f",x"00"),
    10 => (x"4e",x"00",x"00",x"42"),
    11 => (x"00",x"06",x"f9",x"27"),
    12 => (x"fd",x"00",x"0f",x"00"),
    13 => (x"c0",x"f0",x"c1",x"87"),
    14 => (x"00",x"42",x"27",x"4e"),
    15 => (x"00",x"0f",x"00",x"00"),
    16 => (x"4f",x"4f",x"87",x"fd"),
    17 => (x"1e",x"1e",x"72",x"1e"),
    18 => (x"6a",x"4a",x"c0",x"ff"),
    19 => (x"98",x"c0",x"c4",x"48"),
    20 => (x"6e",x"58",x"a6",x"c4"),
    21 => (x"87",x"f3",x"ff",x"02"),
    22 => (x"cc",x"7a",x"66",x"cc"),
    23 => (x"26",x"26",x"48",x"66"),
    24 => (x"0e",x"4f",x"26",x"4a"),
    25 => (x"5c",x"5b",x"5a",x"5e"),
    26 => (x"66",x"d4",x"0e",x"5d"),
    27 => (x"13",x"4d",x"c0",x"4b"),
    28 => (x"02",x"9c",x"74",x"4c"),
    29 => (x"74",x"87",x"d9",x"c0"),
    30 => (x"9a",x"ff",x"c3",x"4a"),
    31 => (x"44",x"27",x"1e",x"72"),
    32 => (x"0f",x"00",x"00",x"00"),
    33 => (x"85",x"c1",x"86",x"c4"),
    34 => (x"9c",x"74",x"4c",x"13"),
    35 => (x"87",x"e7",x"ff",x"05"),
    36 => (x"4d",x"26",x"48",x"75"),
    37 => (x"4b",x"26",x"4c",x"26"),
    38 => (x"4f",x"26",x"4a",x"26"),
    39 => (x"5b",x"5a",x"5e",x"0e"),
    40 => (x"1e",x"0e",x"5d",x"5c"),
    41 => (x"27",x"4c",x"66",x"d8"),
    42 => (x"00",x"00",x"18",x"00"),
    43 => (x"27",x"49",x"76",x"4b"),
    44 => (x"00",x"00",x"10",x"48"),
    45 => (x"74",x"4d",x"c0",x"79"),
    46 => (x"c6",x"c0",x"05",x"9c"),
    47 => (x"53",x"f0",x"c0",x"87"),
    48 => (x"74",x"87",x"f4",x"c0"),
    49 => (x"ee",x"c0",x"02",x"9c"),
    50 => (x"72",x"49",x"74",x"87"),
    51 => (x"66",x"e0",x"c0",x"1e"),
    52 => (x"06",x"7d",x"27",x"4a"),
    53 => (x"26",x"0f",x"00",x"00"),
    54 => (x"6e",x"4a",x"71",x"4a"),
    55 => (x"74",x"53",x"12",x"82"),
    56 => (x"c0",x"1e",x"72",x"49"),
    57 => (x"27",x"4a",x"66",x"e0"),
    58 => (x"00",x"00",x"06",x"7d"),
    59 => (x"70",x"4a",x"26",x"0f"),
    60 => (x"05",x"9c",x"74",x"4c"),
    61 => (x"27",x"87",x"d2",x"ff"),
    62 => (x"00",x"00",x"18",x"00"),
    63 => (x"ea",x"c0",x"02",x"ab"),
    64 => (x"66",x"e0",x"c0",x"87"),
    65 => (x"66",x"e4",x"c0",x"4c"),
    66 => (x"97",x"8b",x"c1",x"1e"),
    67 => (x"c0",x"c1",x"4a",x"6b"),
    68 => (x"92",x"c0",x"c0",x"c0"),
    69 => (x"92",x"b7",x"c0",x"c4"),
    70 => (x"74",x"1e",x"72",x"4a"),
    71 => (x"c1",x"86",x"c8",x"0f"),
    72 => (x"18",x"00",x"27",x"85"),
    73 => (x"05",x"ab",x"00",x"00"),
    74 => (x"75",x"87",x"da",x"ff"),
    75 => (x"4d",x"26",x"26",x"48"),
    76 => (x"4b",x"26",x"4c",x"26"),
    77 => (x"4f",x"26",x"4a",x"26"),
    78 => (x"5b",x"5a",x"5e",x"0e"),
    79 => (x"d4",x"0e",x"5d",x"5c"),
    80 => (x"4d",x"ff",x"4c",x"66"),
    81 => (x"c0",x"c1",x"4b",x"14"),
    82 => (x"93",x"c0",x"c0",x"c0"),
    83 => (x"93",x"b7",x"c0",x"c4"),
    84 => (x"02",x"9b",x"73",x"4b"),
    85 => (x"c1",x"87",x"e8",x"c0"),
    86 => (x"1e",x"66",x"dc",x"85"),
    87 => (x"e0",x"c0",x"1e",x"73"),
    88 => (x"86",x"c8",x"0f",x"66"),
    89 => (x"aa",x"73",x"4a",x"70"),
    90 => (x"87",x"d3",x"c0",x"05"),
    91 => (x"c0",x"c1",x"4b",x"14"),
    92 => (x"93",x"c0",x"c0",x"c0"),
    93 => (x"93",x"b7",x"c0",x"c4"),
    94 => (x"05",x"9b",x"73",x"4b"),
    95 => (x"75",x"87",x"d8",x"ff"),
    96 => (x"26",x"4d",x"26",x"48"),
    97 => (x"26",x"4b",x"26",x"4c"),
    98 => (x"0e",x"4f",x"26",x"4a"),
    99 => (x"5c",x"5b",x"5a",x"5e"),
   100 => (x"8e",x"cc",x"0e",x"5d"),
   101 => (x"4b",x"66",x"e8",x"c0"),
   102 => (x"a6",x"c4",x"4c",x"c0"),
   103 => (x"c0",x"79",x"c0",x"49"),
   104 => (x"bf",x"97",x"66",x"e0"),
   105 => (x"c0",x"c0",x"c1",x"4d"),
   106 => (x"c4",x"95",x"c0",x"c0"),
   107 => (x"4d",x"95",x"b7",x"c0"),
   108 => (x"48",x"66",x"e0",x"c0"),
   109 => (x"e4",x"c0",x"80",x"c1"),
   110 => (x"9d",x"75",x"58",x"a6"),
   111 => (x"87",x"ce",x"c5",x"02"),
   112 => (x"c4",x"02",x"66",x"c4"),
   113 => (x"a6",x"c8",x"87",x"ce"),
   114 => (x"c4",x"79",x"c0",x"49"),
   115 => (x"79",x"c0",x"49",x"a6"),
   116 => (x"f0",x"c0",x"4a",x"75"),
   117 => (x"e8",x"c1",x"02",x"ad"),
   118 => (x"aa",x"e3",x"c1",x"87"),
   119 => (x"87",x"e9",x"c1",x"02"),
   120 => (x"02",x"aa",x"e4",x"c1"),
   121 => (x"c1",x"87",x"e6",x"c0"),
   122 => (x"c1",x"02",x"aa",x"ec"),
   123 => (x"f0",x"c1",x"87",x"d3"),
   124 => (x"e0",x"c0",x"02",x"aa"),
   125 => (x"aa",x"f3",x"c1",x"87"),
   126 => (x"87",x"e1",x"c0",x"02"),
   127 => (x"02",x"aa",x"f5",x"c1"),
   128 => (x"c1",x"87",x"ca",x"c0"),
   129 => (x"c0",x"02",x"aa",x"f8"),
   130 => (x"db",x"c1",x"87",x"cb"),
   131 => (x"49",x"a6",x"c8",x"87"),
   132 => (x"ea",x"c1",x"79",x"ca"),
   133 => (x"49",x"a6",x"c8",x"87"),
   134 => (x"e2",x"c1",x"79",x"d0"),
   135 => (x"66",x"ec",x"c0",x"87"),
   136 => (x"c0",x"1e",x"73",x"1e"),
   137 => (x"c4",x"48",x"66",x"ec"),
   138 => (x"a6",x"f0",x"c0",x"80"),
   139 => (x"66",x"ec",x"c0",x"58"),
   140 => (x"6a",x"8a",x"c4",x"4a"),
   141 => (x"87",x"c0",x"fc",x"1e"),
   142 => (x"4a",x"70",x"86",x"cc"),
   143 => (x"fe",x"c0",x"84",x"72"),
   144 => (x"49",x"a6",x"c4",x"87"),
   145 => (x"f6",x"c0",x"79",x"c1"),
   146 => (x"66",x"ec",x"c0",x"87"),
   147 => (x"66",x"e8",x"c0",x"1e"),
   148 => (x"c0",x"80",x"c4",x"48"),
   149 => (x"c0",x"58",x"a6",x"ec"),
   150 => (x"c4",x"4a",x"66",x"e8"),
   151 => (x"73",x"1e",x"6a",x"8a"),
   152 => (x"c1",x"86",x"c8",x"0f"),
   153 => (x"87",x"d7",x"c0",x"84"),
   154 => (x"1e",x"66",x"ec",x"c0"),
   155 => (x"73",x"1e",x"e5",x"c0"),
   156 => (x"c0",x"86",x"c8",x"0f"),
   157 => (x"75",x"1e",x"66",x"ec"),
   158 => (x"c8",x"0f",x"73",x"1e"),
   159 => (x"c8",x"84",x"c1",x"86"),
   160 => (x"e8",x"c1",x"02",x"66"),
   161 => (x"66",x"e4",x"c0",x"87"),
   162 => (x"c0",x"80",x"c4",x"48"),
   163 => (x"c0",x"58",x"a6",x"e8"),
   164 => (x"c4",x"4a",x"66",x"e4"),
   165 => (x"6a",x"49",x"76",x"8a"),
   166 => (x"ad",x"e4",x"c1",x"79"),
   167 => (x"87",x"dc",x"c0",x"05"),
   168 => (x"b7",x"c0",x"49",x"6e"),
   169 => (x"d3",x"c0",x"03",x"a9"),
   170 => (x"1e",x"ed",x"c0",x"87"),
   171 => (x"00",x"00",x"44",x"27"),
   172 => (x"86",x"c4",x"0f",x"00"),
   173 => (x"08",x"c0",x"48",x"6e"),
   174 => (x"58",x"a6",x"c4",x"88"),
   175 => (x"1e",x"66",x"ec",x"c0"),
   176 => (x"66",x"d0",x"1e",x"73"),
   177 => (x"1e",x"66",x"cc",x"1e"),
   178 => (x"d0",x"87",x"d1",x"f7"),
   179 => (x"72",x"4a",x"70",x"86"),
   180 => (x"87",x"d9",x"c0",x"84"),
   181 => (x"05",x"ad",x"e5",x"c0"),
   182 => (x"c4",x"87",x"c8",x"c0"),
   183 => (x"79",x"c1",x"49",x"a6"),
   184 => (x"c0",x"87",x"ca",x"c0"),
   185 => (x"75",x"1e",x"66",x"ec"),
   186 => (x"c8",x"0f",x"73",x"1e"),
   187 => (x"66",x"e0",x"c0",x"86"),
   188 => (x"c1",x"4d",x"bf",x"97"),
   189 => (x"c0",x"c0",x"c0",x"c0"),
   190 => (x"b7",x"c0",x"c4",x"95"),
   191 => (x"e0",x"c0",x"4d",x"95"),
   192 => (x"80",x"c1",x"48",x"66"),
   193 => (x"58",x"a6",x"e4",x"c0"),
   194 => (x"fa",x"05",x"9d",x"75"),
   195 => (x"48",x"74",x"87",x"f2"),
   196 => (x"4d",x"26",x"86",x"cc"),
   197 => (x"4b",x"26",x"4c",x"26"),
   198 => (x"4f",x"26",x"4a",x"26"),
   199 => (x"c0",x"1e",x"72",x"1e"),
   200 => (x"00",x"44",x"27",x"1e"),
   201 => (x"d4",x"1e",x"00",x"00"),
   202 => (x"66",x"d4",x"1e",x"66"),
   203 => (x"01",x"8b",x"27",x"1e"),
   204 => (x"d0",x"0f",x"00",x"00"),
   205 => (x"72",x"4a",x"70",x"86"),
   206 => (x"26",x"4a",x"26",x"48"),
   207 => (x"1e",x"72",x"1e",x"4f"),
   208 => (x"c0",x"4a",x"a6",x"cc"),
   209 => (x"00",x"44",x"27",x"1e"),
   210 => (x"72",x"1e",x"00",x"00"),
   211 => (x"1e",x"66",x"d4",x"1e"),
   212 => (x"00",x"01",x"8b",x"27"),
   213 => (x"86",x"d0",x"0f",x"00"),
   214 => (x"48",x"72",x"4a",x"70"),
   215 => (x"4f",x"26",x"4a",x"26"),
   216 => (x"5b",x"5a",x"5e",x"0e"),
   217 => (x"4b",x"66",x"d0",x"0e"),
   218 => (x"c4",x"4a",x"66",x"d0"),
   219 => (x"c0",x"02",x"6a",x"82"),
   220 => (x"4a",x"73",x"87",x"dc"),
   221 => (x"48",x"6a",x"82",x"c4"),
   222 => (x"7a",x"70",x"88",x"c1"),
   223 => (x"48",x"72",x"4a",x"6b"),
   224 => (x"7b",x"70",x"80",x"c1"),
   225 => (x"52",x"66",x"cc",x"97"),
   226 => (x"c0",x"48",x"66",x"cc"),
   227 => (x"48",x"c0",x"87",x"c2"),
   228 => (x"4a",x"26",x"4b",x"26"),
   229 => (x"5e",x"0e",x"4f",x"26"),
   230 => (x"c8",x"0e",x"5b",x"5a"),
   231 => (x"d4",x"49",x"76",x"8e"),
   232 => (x"a6",x"c4",x"79",x"66"),
   233 => (x"dc",x"79",x"ff",x"49"),
   234 => (x"4b",x"76",x"4a",x"a6"),
   235 => (x"60",x"27",x"1e",x"73"),
   236 => (x"1e",x"00",x"00",x"03"),
   237 => (x"e4",x"c0",x"1e",x"72"),
   238 => (x"8b",x"27",x"1e",x"66"),
   239 => (x"0f",x"00",x"00",x"01"),
   240 => (x"4a",x"70",x"86",x"d0"),
   241 => (x"86",x"c8",x"48",x"72"),
   242 => (x"4a",x"26",x"4b",x"26"),
   243 => (x"5e",x"0e",x"4f",x"26"),
   244 => (x"c8",x"0e",x"5b",x"5a"),
   245 => (x"d4",x"49",x"76",x"8e"),
   246 => (x"a6",x"c4",x"79",x"66"),
   247 => (x"79",x"66",x"d8",x"49"),
   248 => (x"4a",x"a6",x"e0",x"c0"),
   249 => (x"1e",x"73",x"4b",x"76"),
   250 => (x"00",x"03",x"60",x"27"),
   251 => (x"1e",x"72",x"1e",x"00"),
   252 => (x"1e",x"66",x"e8",x"c0"),
   253 => (x"00",x"01",x"8b",x"27"),
   254 => (x"86",x"d0",x"0f",x"00"),
   255 => (x"48",x"72",x"4a",x"70"),
   256 => (x"4b",x"26",x"86",x"c8"),
   257 => (x"4f",x"26",x"4a",x"26"),
   258 => (x"c8",x"1e",x"72",x"1e"),
   259 => (x"d0",x"49",x"76",x"8e"),
   260 => (x"a6",x"c4",x"79",x"66"),
   261 => (x"76",x"79",x"ff",x"49"),
   262 => (x"27",x"1e",x"72",x"4a"),
   263 => (x"00",x"00",x"03",x"60"),
   264 => (x"66",x"e0",x"c0",x"1e"),
   265 => (x"66",x"e0",x"c0",x"1e"),
   266 => (x"01",x"8b",x"27",x"1e"),
   267 => (x"d0",x"0f",x"00",x"00"),
   268 => (x"72",x"4a",x"70",x"86"),
   269 => (x"26",x"86",x"c8",x"48"),
   270 => (x"0e",x"4f",x"26",x"4a"),
   271 => (x"0e",x"5b",x"5a",x"5e"),
   272 => (x"cc",x"4b",x"66",x"d0"),
   273 => (x"66",x"cc",x"7b",x"66"),
   274 => (x"06",x"6a",x"27",x"1e"),
   275 => (x"c4",x"0f",x"00",x"00"),
   276 => (x"72",x"4a",x"70",x"86"),
   277 => (x"c2",x"c0",x"05",x"9a"),
   278 => (x"cc",x"7b",x"c3",x"87"),
   279 => (x"66",x"cc",x"4a",x"66"),
   280 => (x"02",x"a9",x"c0",x"49"),
   281 => (x"c1",x"87",x"db",x"c0"),
   282 => (x"da",x"c0",x"02",x"aa"),
   283 => (x"02",x"aa",x"c2",x"87"),
   284 => (x"c3",x"87",x"ed",x"c0"),
   285 => (x"ee",x"c0",x"02",x"aa"),
   286 => (x"02",x"aa",x"c4",x"87"),
   287 => (x"c0",x"87",x"e6",x"c0"),
   288 => (x"7b",x"c0",x"87",x"e5"),
   289 => (x"27",x"87",x"e0",x"c0"),
   290 => (x"00",x"00",x"18",x"18"),
   291 => (x"e4",x"c1",x"49",x"bf"),
   292 => (x"c0",x"06",x"a9",x"b7"),
   293 => (x"7b",x"c0",x"87",x"c5"),
   294 => (x"c3",x"87",x"cc",x"c0"),
   295 => (x"87",x"c7",x"c0",x"7b"),
   296 => (x"c2",x"c0",x"7b",x"c1"),
   297 => (x"26",x"7b",x"c2",x"87"),
   298 => (x"26",x"4a",x"26",x"4b"),
   299 => (x"1e",x"72",x"1e",x"4f"),
   300 => (x"c2",x"4a",x"66",x"c8"),
   301 => (x"48",x"66",x"cc",x"82"),
   302 => (x"66",x"d0",x"80",x"72"),
   303 => (x"26",x"79",x"70",x"49"),
   304 => (x"0e",x"4f",x"26",x"4a"),
   305 => (x"5c",x"5b",x"5a",x"5e"),
   306 => (x"c0",x"1e",x"0e",x"5d"),
   307 => (x"c5",x"4d",x"66",x"e0"),
   308 => (x"c4",x"4c",x"75",x"85"),
   309 => (x"84",x"66",x"d8",x"94"),
   310 => (x"7c",x"66",x"e4",x"c0"),
   311 => (x"82",x"c1",x"4a",x"75"),
   312 => (x"93",x"c4",x"4b",x"72"),
   313 => (x"6c",x"83",x"66",x"d8"),
   314 => (x"de",x"4b",x"75",x"7b"),
   315 => (x"d8",x"93",x"c4",x"83"),
   316 => (x"7b",x"75",x"83",x"66"),
   317 => (x"79",x"75",x"49",x"76"),
   318 => (x"01",x"ad",x"b7",x"72"),
   319 => (x"6e",x"87",x"df",x"c0"),
   320 => (x"c3",x"4b",x"75",x"4c"),
   321 => (x"66",x"dc",x"93",x"c8"),
   322 => (x"c4",x"4a",x"74",x"83"),
   323 => (x"75",x"82",x"73",x"92"),
   324 => (x"75",x"84",x"c1",x"7a"),
   325 => (x"72",x"82",x"c1",x"4a"),
   326 => (x"ff",x"06",x"ac",x"b7"),
   327 => (x"4b",x"75",x"87",x"e3"),
   328 => (x"dc",x"93",x"c8",x"c3"),
   329 => (x"4a",x"75",x"83",x"66"),
   330 => (x"92",x"c4",x"8a",x"c1"),
   331 => (x"48",x"6a",x"82",x"73"),
   332 => (x"7a",x"70",x"80",x"c1"),
   333 => (x"92",x"c4",x"4a",x"75"),
   334 => (x"72",x"4b",x"66",x"d8"),
   335 => (x"d4",x"4c",x"75",x"83"),
   336 => (x"94",x"c8",x"c3",x"84"),
   337 => (x"74",x"84",x"66",x"dc"),
   338 => (x"27",x"7a",x"6b",x"82"),
   339 => (x"00",x"00",x"18",x"18"),
   340 => (x"26",x"79",x"c5",x"49"),
   341 => (x"4c",x"26",x"4d",x"26"),
   342 => (x"4a",x"26",x"4b",x"26"),
   343 => (x"5e",x"0e",x"4f",x"26"),
   344 => (x"0e",x"5c",x"5b",x"5a"),
   345 => (x"4c",x"66",x"d0",x"97"),
   346 => (x"c0",x"c1",x"4b",x"74"),
   347 => (x"93",x"c0",x"c0",x"c0"),
   348 => (x"93",x"b7",x"c0",x"c4"),
   349 => (x"66",x"d4",x"97",x"4b"),
   350 => (x"c0",x"c0",x"c1",x"4a"),
   351 => (x"c4",x"92",x"c0",x"c0"),
   352 => (x"4a",x"92",x"b7",x"c0"),
   353 => (x"02",x"ab",x"b7",x"72"),
   354 => (x"c0",x"87",x"c5",x"c0"),
   355 => (x"87",x"ca",x"c0",x"48"),
   356 => (x"00",x"18",x"20",x"27"),
   357 => (x"51",x"74",x"49",x"00"),
   358 => (x"4c",x"26",x"48",x"c1"),
   359 => (x"4a",x"26",x"4b",x"26"),
   360 => (x"5e",x"0e",x"4f",x"26"),
   361 => (x"0e",x"5c",x"5b",x"5a"),
   362 => (x"4c",x"6e",x"97",x"1e"),
   363 => (x"66",x"d8",x"4b",x"c2"),
   364 => (x"73",x"82",x"c1",x"4a"),
   365 => (x"4a",x"6a",x"97",x"82"),
   366 => (x"c0",x"c0",x"c0",x"c1"),
   367 => (x"c0",x"c4",x"92",x"c0"),
   368 => (x"72",x"4a",x"92",x"b7"),
   369 => (x"4a",x"66",x"d8",x"1e"),
   370 => (x"6a",x"97",x"82",x"73"),
   371 => (x"c0",x"c0",x"c1",x"4a"),
   372 => (x"c4",x"92",x"c0",x"c0"),
   373 => (x"4a",x"92",x"b7",x"c0"),
   374 => (x"5e",x"27",x"1e",x"72"),
   375 => (x"0f",x"00",x"00",x"05"),
   376 => (x"4a",x"70",x"86",x"c8"),
   377 => (x"c0",x"05",x"9a",x"72"),
   378 => (x"c1",x"c1",x"87",x"c5"),
   379 => (x"c2",x"83",x"c1",x"4c"),
   380 => (x"fe",x"06",x"ab",x"b7"),
   381 => (x"4a",x"74",x"87",x"f8"),
   382 => (x"c0",x"c0",x"c0",x"c1"),
   383 => (x"c0",x"c4",x"92",x"c0"),
   384 => (x"c1",x"4a",x"92",x"b7"),
   385 => (x"04",x"aa",x"b7",x"d7"),
   386 => (x"74",x"87",x"d7",x"c0"),
   387 => (x"c0",x"c0",x"c1",x"4a"),
   388 => (x"c4",x"92",x"c0",x"c0"),
   389 => (x"4a",x"92",x"b7",x"c0"),
   390 => (x"aa",x"b7",x"da",x"c1"),
   391 => (x"87",x"c2",x"c0",x"03"),
   392 => (x"4a",x"74",x"4b",x"c7"),
   393 => (x"c0",x"c0",x"c0",x"c1"),
   394 => (x"c0",x"c4",x"92",x"c0"),
   395 => (x"c1",x"4a",x"92",x"b7"),
   396 => (x"c0",x"05",x"aa",x"d2"),
   397 => (x"48",x"c1",x"87",x"c5"),
   398 => (x"d4",x"87",x"e6",x"c0"),
   399 => (x"66",x"d8",x"4a",x"66"),
   400 => (x"06",x"e1",x"27",x"49"),
   401 => (x"70",x"0f",x"00",x"00"),
   402 => (x"aa",x"b7",x"c0",x"4a"),
   403 => (x"87",x"cf",x"c0",x"06"),
   404 => (x"80",x"c7",x"48",x"73"),
   405 => (x"00",x"18",x"1c",x"27"),
   406 => (x"48",x"c1",x"58",x"00"),
   407 => (x"c0",x"87",x"c2",x"c0"),
   408 => (x"4c",x"26",x"26",x"48"),
   409 => (x"4a",x"26",x"4b",x"26"),
   410 => (x"c4",x"1e",x"4f",x"26"),
   411 => (x"a9",x"c2",x"49",x"66"),
   412 => (x"87",x"c5",x"c0",x"05"),
   413 => (x"c2",x"c0",x"48",x"c1"),
   414 => (x"26",x"48",x"c0",x"87"),
   415 => (x"1e",x"73",x"1e",x"4f"),
   416 => (x"e7",x"02",x"9a",x"72"),
   417 => (x"c1",x"48",x"c0",x"87"),
   418 => (x"06",x"a9",x"72",x"4b"),
   419 => (x"82",x"72",x"87",x"d1"),
   420 => (x"73",x"87",x"c9",x"06"),
   421 => (x"01",x"a9",x"72",x"83"),
   422 => (x"87",x"c3",x"87",x"f4"),
   423 => (x"72",x"3a",x"b2",x"c1"),
   424 => (x"73",x"89",x"03",x"a9"),
   425 => (x"2a",x"c1",x"07",x"80"),
   426 => (x"87",x"f3",x"05",x"2b"),
   427 => (x"4f",x"26",x"4b",x"26"),
   428 => (x"c4",x"1e",x"75",x"1e"),
   429 => (x"a1",x"b7",x"71",x"4d"),
   430 => (x"c1",x"b9",x"ff",x"04"),
   431 => (x"07",x"bd",x"c3",x"81"),
   432 => (x"04",x"a2",x"b7",x"72"),
   433 => (x"82",x"c1",x"ba",x"ff"),
   434 => (x"fe",x"07",x"bd",x"c1"),
   435 => (x"2d",x"c1",x"87",x"ef"),
   436 => (x"c1",x"b8",x"ff",x"04"),
   437 => (x"04",x"2d",x"07",x"80"),
   438 => (x"81",x"c1",x"b9",x"ff"),
   439 => (x"26",x"4d",x"26",x"07"),
   440 => (x"1e",x"72",x"1e",x"4f"),
   441 => (x"02",x"11",x"48",x"12"),
   442 => (x"02",x"88",x"87",x"c4"),
   443 => (x"4a",x"26",x"87",x"f6"),
   444 => (x"ff",x"1e",x"4f",x"26"),
   445 => (x"26",x"48",x"bf",x"c8"),
   446 => (x"5a",x"5e",x"0e",x"4f"),
   447 => (x"0e",x"5d",x"5c",x"5b"),
   448 => (x"66",x"c4",x"8e",x"d0"),
   449 => (x"18",x"14",x"27",x"4c"),
   450 => (x"27",x"49",x"00",x"00"),
   451 => (x"00",x"00",x"40",x"18"),
   452 => (x"18",x"10",x"27",x"79"),
   453 => (x"27",x"49",x"00",x"00"),
   454 => (x"00",x"00",x"40",x"48"),
   455 => (x"40",x"48",x"27",x"79"),
   456 => (x"27",x"49",x"00",x"00"),
   457 => (x"00",x"00",x"40",x"18"),
   458 => (x"40",x"4c",x"27",x"79"),
   459 => (x"c0",x"49",x"00",x"00"),
   460 => (x"40",x"50",x"27",x"79"),
   461 => (x"c2",x"49",x"00",x"00"),
   462 => (x"40",x"54",x"27",x"79"),
   463 => (x"c0",x"49",x"00",x"00"),
   464 => (x"58",x"27",x"79",x"e8"),
   465 => (x"49",x"00",x"00",x"40"),
   466 => (x"00",x"11",x"d2",x"27"),
   467 => (x"1e",x"72",x"48",x"00"),
   468 => (x"41",x"20",x"41",x"20"),
   469 => (x"41",x"20",x"41",x"20"),
   470 => (x"41",x"20",x"41",x"20"),
   471 => (x"51",x"10",x"41",x"20"),
   472 => (x"51",x"10",x"51",x"10"),
   473 => (x"78",x"27",x"4a",x"26"),
   474 => (x"49",x"00",x"00",x"40"),
   475 => (x"00",x"11",x"f1",x"27"),
   476 => (x"1e",x"72",x"48",x"00"),
   477 => (x"41",x"20",x"41",x"20"),
   478 => (x"41",x"20",x"41",x"20"),
   479 => (x"41",x"20",x"41",x"20"),
   480 => (x"51",x"10",x"41",x"20"),
   481 => (x"51",x"10",x"51",x"10"),
   482 => (x"4c",x"27",x"4a",x"26"),
   483 => (x"49",x"00",x"00",x"1f"),
   484 => (x"10",x"27",x"79",x"ca"),
   485 => (x"1e",x"00",x"00",x"12"),
   486 => (x"00",x"03",x"3d",x"27"),
   487 => (x"86",x"c4",x"0f",x"00"),
   488 => (x"00",x"12",x"12",x"27"),
   489 => (x"3d",x"27",x"1e",x"00"),
   490 => (x"0f",x"00",x"00",x"03"),
   491 => (x"42",x"27",x"86",x"c4"),
   492 => (x"1e",x"00",x"00",x"12"),
   493 => (x"00",x"03",x"3d",x"27"),
   494 => (x"86",x"c4",x"0f",x"00"),
   495 => (x"00",x"17",x"f8",x"27"),
   496 => (x"c0",x"02",x"bf",x"00"),
   497 => (x"59",x"27",x"87",x"df"),
   498 => (x"1e",x"00",x"00",x"10"),
   499 => (x"00",x"03",x"3d",x"27"),
   500 => (x"86",x"c4",x"0f",x"00"),
   501 => (x"00",x"10",x"85",x"27"),
   502 => (x"3d",x"27",x"1e",x"00"),
   503 => (x"0f",x"00",x"00",x"03"),
   504 => (x"dc",x"c0",x"86",x"c4"),
   505 => (x"10",x"87",x"27",x"87"),
   506 => (x"27",x"1e",x"00",x"00"),
   507 => (x"00",x"00",x"03",x"3d"),
   508 => (x"27",x"86",x"c4",x"0f"),
   509 => (x"00",x"00",x"10",x"b6"),
   510 => (x"03",x"3d",x"27",x"1e"),
   511 => (x"c4",x"0f",x"00",x"00"),
   512 => (x"17",x"fc",x"27",x"86"),
   513 => (x"1e",x"bf",x"00",x"00"),
   514 => (x"00",x"12",x"44",x"27"),
   515 => (x"3d",x"27",x"1e",x"00"),
   516 => (x"0f",x"00",x"00",x"03"),
   517 => (x"f2",x"27",x"86",x"c8"),
   518 => (x"0f",x"00",x"00",x"06"),
   519 => (x"00",x"40",x"04",x"27"),
   520 => (x"4d",x"c1",x"58",x"00"),
   521 => (x"00",x"17",x"fc",x"27"),
   522 => (x"c0",x"49",x"bf",x"00"),
   523 => (x"c6",x"06",x"a9",x"b7"),
   524 => (x"33",x"27",x"87",x"f2"),
   525 => (x"0f",x"00",x"00",x"10"),
   526 => (x"00",x"0f",x"f3",x"27"),
   527 => (x"49",x"76",x"0f",x"00"),
   528 => (x"4c",x"c3",x"79",x"c2"),
   529 => (x"00",x"40",x"98",x"27"),
   530 => (x"d7",x"27",x"49",x"00"),
   531 => (x"48",x"00",x"00",x"10"),
   532 => (x"41",x"20",x"1e",x"72"),
   533 => (x"41",x"20",x"41",x"20"),
   534 => (x"41",x"20",x"41",x"20"),
   535 => (x"41",x"20",x"41",x"20"),
   536 => (x"51",x"10",x"51",x"10"),
   537 => (x"4a",x"26",x"51",x"10"),
   538 => (x"c1",x"49",x"a6",x"c8"),
   539 => (x"40",x"98",x"27",x"79"),
   540 => (x"27",x"1e",x"00",x"00"),
   541 => (x"00",x"00",x"40",x"78"),
   542 => (x"05",x"a2",x"27",x"1e"),
   543 => (x"c8",x"0f",x"00",x"00"),
   544 => (x"72",x"4a",x"70",x"86"),
   545 => (x"c5",x"c0",x"05",x"9a"),
   546 => (x"c0",x"4a",x"c1",x"87"),
   547 => (x"4a",x"c0",x"87",x"c2"),
   548 => (x"00",x"18",x"1c",x"27"),
   549 => (x"79",x"72",x"49",x"00"),
   550 => (x"06",x"ac",x"b7",x"6e"),
   551 => (x"6e",x"87",x"eb",x"c0"),
   552 => (x"72",x"92",x"c5",x"4a"),
   553 => (x"d0",x"88",x"74",x"48"),
   554 => (x"a6",x"cc",x"58",x"a6"),
   555 => (x"74",x"1e",x"72",x"4a"),
   556 => (x"1e",x"66",x"c8",x"1e"),
   557 => (x"00",x"04",x"ad",x"27"),
   558 => (x"86",x"cc",x"0f",x"00"),
   559 => (x"80",x"c1",x"48",x"6e"),
   560 => (x"6e",x"58",x"a6",x"c4"),
   561 => (x"ff",x"01",x"ac",x"b7"),
   562 => (x"66",x"cc",x"87",x"d5"),
   563 => (x"1e",x"66",x"c4",x"1e"),
   564 => (x"00",x"18",x"f0",x"27"),
   565 => (x"28",x"27",x"1e",x"00"),
   566 => (x"1e",x"00",x"00",x"18"),
   567 => (x"00",x"04",x"c3",x"27"),
   568 => (x"86",x"d0",x"0f",x"00"),
   569 => (x"00",x"18",x"10",x"27"),
   570 => (x"27",x"1e",x"bf",x"00"),
   571 => (x"00",x"00",x"0e",x"d6"),
   572 => (x"c4",x"86",x"c4",x"0f"),
   573 => (x"c1",x"c1",x"49",x"a6"),
   574 => (x"18",x"21",x"27",x"51"),
   575 => (x"bf",x"97",x"00",x"00"),
   576 => (x"c0",x"c0",x"c1",x"4a"),
   577 => (x"c4",x"92",x"c0",x"c0"),
   578 => (x"4a",x"92",x"b7",x"c0"),
   579 => (x"aa",x"b7",x"c1",x"c1"),
   580 => (x"87",x"d5",x"c2",x"04"),
   581 => (x"97",x"1e",x"c3",x"c1"),
   582 => (x"c1",x"4a",x"66",x"c8"),
   583 => (x"c0",x"c0",x"c0",x"c0"),
   584 => (x"b7",x"c0",x"c4",x"92"),
   585 => (x"1e",x"72",x"4a",x"92"),
   586 => (x"00",x"05",x"5e",x"27"),
   587 => (x"86",x"c8",x"0f",x"00"),
   588 => (x"66",x"c8",x"4a",x"70"),
   589 => (x"fd",x"c0",x"05",x"aa"),
   590 => (x"4a",x"a6",x"c8",x"87"),
   591 => (x"1e",x"c0",x"1e",x"72"),
   592 => (x"00",x"04",x"3b",x"27"),
   593 => (x"86",x"c8",x"0f",x"00"),
   594 => (x"00",x"40",x"98",x"27"),
   595 => (x"b8",x"27",x"49",x"00"),
   596 => (x"48",x"00",x"00",x"10"),
   597 => (x"41",x"20",x"1e",x"72"),
   598 => (x"41",x"20",x"41",x"20"),
   599 => (x"41",x"20",x"41",x"20"),
   600 => (x"41",x"20",x"41",x"20"),
   601 => (x"51",x"10",x"51",x"10"),
   602 => (x"4a",x"26",x"51",x"10"),
   603 => (x"18",x"27",x"4c",x"75"),
   604 => (x"49",x"00",x"00",x"18"),
   605 => (x"c4",x"97",x"79",x"75"),
   606 => (x"80",x"c1",x"48",x"66"),
   607 => (x"50",x"08",x"a6",x"c4"),
   608 => (x"4b",x"66",x"c4",x"97"),
   609 => (x"c0",x"c0",x"c0",x"c1"),
   610 => (x"c0",x"c4",x"93",x"c0"),
   611 => (x"27",x"4b",x"93",x"b7"),
   612 => (x"00",x"00",x"18",x"21"),
   613 => (x"c1",x"4a",x"bf",x"97"),
   614 => (x"c0",x"c0",x"c0",x"c0"),
   615 => (x"b7",x"c0",x"c4",x"92"),
   616 => (x"b7",x"72",x"4a",x"92"),
   617 => (x"eb",x"fd",x"06",x"ab"),
   618 => (x"74",x"94",x"6e",x"87"),
   619 => (x"d0",x"1e",x"72",x"49"),
   620 => (x"b0",x"27",x"4a",x"66"),
   621 => (x"0f",x"00",x"00",x"06"),
   622 => (x"48",x"70",x"4a",x"26"),
   623 => (x"74",x"58",x"a6",x"c4"),
   624 => (x"8a",x"66",x"cc",x"4a"),
   625 => (x"4c",x"72",x"92",x"c7"),
   626 => (x"4a",x"76",x"8c",x"6e"),
   627 => (x"70",x"27",x"1e",x"72"),
   628 => (x"0f",x"00",x"00",x"0f"),
   629 => (x"85",x"c1",x"86",x"c4"),
   630 => (x"00",x"17",x"fc",x"27"),
   631 => (x"ad",x"b7",x"bf",x"00"),
   632 => (x"87",x"ce",x"f9",x"06"),
   633 => (x"00",x"06",x"f2",x"27"),
   634 => (x"08",x"27",x"0f",x"00"),
   635 => (x"58",x"00",x"00",x"40"),
   636 => (x"00",x"12",x"71",x"27"),
   637 => (x"3d",x"27",x"1e",x"00"),
   638 => (x"0f",x"00",x"00",x"03"),
   639 => (x"81",x"27",x"86",x"c4"),
   640 => (x"1e",x"00",x"00",x"12"),
   641 => (x"00",x"03",x"3d",x"27"),
   642 => (x"86",x"c4",x"0f",x"00"),
   643 => (x"00",x"12",x"83",x"27"),
   644 => (x"3d",x"27",x"1e",x"00"),
   645 => (x"0f",x"00",x"00",x"03"),
   646 => (x"b9",x"27",x"86",x"c4"),
   647 => (x"1e",x"00",x"00",x"12"),
   648 => (x"00",x"03",x"3d",x"27"),
   649 => (x"86",x"c4",x"0f",x"00"),
   650 => (x"00",x"18",x"18",x"27"),
   651 => (x"27",x"1e",x"bf",x"00"),
   652 => (x"00",x"00",x"12",x"bb"),
   653 => (x"03",x"3d",x"27",x"1e"),
   654 => (x"c8",x"0f",x"00",x"00"),
   655 => (x"27",x"1e",x"c5",x"86"),
   656 => (x"00",x"00",x"12",x"d4"),
   657 => (x"03",x"3d",x"27",x"1e"),
   658 => (x"c8",x"0f",x"00",x"00"),
   659 => (x"18",x"1c",x"27",x"86"),
   660 => (x"1e",x"bf",x"00",x"00"),
   661 => (x"00",x"12",x"ed",x"27"),
   662 => (x"3d",x"27",x"1e",x"00"),
   663 => (x"0f",x"00",x"00",x"03"),
   664 => (x"1e",x"c1",x"86",x"c8"),
   665 => (x"00",x"13",x"06",x"27"),
   666 => (x"3d",x"27",x"1e",x"00"),
   667 => (x"0f",x"00",x"00",x"03"),
   668 => (x"20",x"27",x"86",x"c8"),
   669 => (x"97",x"00",x"00",x"18"),
   670 => (x"c0",x"c1",x"4a",x"bf"),
   671 => (x"92",x"c0",x"c0",x"c0"),
   672 => (x"92",x"b7",x"c0",x"c4"),
   673 => (x"27",x"1e",x"72",x"4a"),
   674 => (x"00",x"00",x"13",x"1f"),
   675 => (x"03",x"3d",x"27",x"1e"),
   676 => (x"c8",x"0f",x"00",x"00"),
   677 => (x"1e",x"c1",x"c1",x"86"),
   678 => (x"00",x"13",x"38",x"27"),
   679 => (x"3d",x"27",x"1e",x"00"),
   680 => (x"0f",x"00",x"00",x"03"),
   681 => (x"21",x"27",x"86",x"c8"),
   682 => (x"97",x"00",x"00",x"18"),
   683 => (x"c0",x"c1",x"4a",x"bf"),
   684 => (x"92",x"c0",x"c0",x"c0"),
   685 => (x"92",x"b7",x"c0",x"c4"),
   686 => (x"27",x"1e",x"72",x"4a"),
   687 => (x"00",x"00",x"13",x"51"),
   688 => (x"03",x"3d",x"27",x"1e"),
   689 => (x"c8",x"0f",x"00",x"00"),
   690 => (x"1e",x"c2",x"c1",x"86"),
   691 => (x"00",x"13",x"6a",x"27"),
   692 => (x"3d",x"27",x"1e",x"00"),
   693 => (x"0f",x"00",x"00",x"03"),
   694 => (x"48",x"27",x"86",x"c8"),
   695 => (x"bf",x"00",x"00",x"18"),
   696 => (x"13",x"83",x"27",x"1e"),
   697 => (x"27",x"1e",x"00",x"00"),
   698 => (x"00",x"00",x"03",x"3d"),
   699 => (x"c7",x"86",x"c8",x"0f"),
   700 => (x"13",x"9c",x"27",x"1e"),
   701 => (x"27",x"1e",x"00",x"00"),
   702 => (x"00",x"00",x"03",x"3d"),
   703 => (x"27",x"86",x"c8",x"0f"),
   704 => (x"00",x"00",x"1f",x"4c"),
   705 => (x"b5",x"27",x"1e",x"bf"),
   706 => (x"1e",x"00",x"00",x"13"),
   707 => (x"00",x"03",x"3d",x"27"),
   708 => (x"86",x"c8",x"0f",x"00"),
   709 => (x"00",x"13",x"ce",x"27"),
   710 => (x"3d",x"27",x"1e",x"00"),
   711 => (x"0f",x"00",x"00",x"03"),
   712 => (x"f8",x"27",x"86",x"c4"),
   713 => (x"1e",x"00",x"00",x"13"),
   714 => (x"00",x"03",x"3d",x"27"),
   715 => (x"86",x"c4",x"0f",x"00"),
   716 => (x"00",x"18",x"10",x"27"),
   717 => (x"1e",x"bf",x"bf",x"00"),
   718 => (x"00",x"14",x"04",x"27"),
   719 => (x"3d",x"27",x"1e",x"00"),
   720 => (x"0f",x"00",x"00",x"03"),
   721 => (x"1d",x"27",x"86",x"c8"),
   722 => (x"1e",x"00",x"00",x"14"),
   723 => (x"00",x"03",x"3d",x"27"),
   724 => (x"86",x"c4",x"0f",x"00"),
   725 => (x"00",x"18",x"10",x"27"),
   726 => (x"c4",x"4a",x"bf",x"00"),
   727 => (x"27",x"1e",x"6a",x"82"),
   728 => (x"00",x"00",x"14",x"4e"),
   729 => (x"03",x"3d",x"27",x"1e"),
   730 => (x"c8",x"0f",x"00",x"00"),
   731 => (x"27",x"1e",x"c0",x"86"),
   732 => (x"00",x"00",x"14",x"67"),
   733 => (x"03",x"3d",x"27",x"1e"),
   734 => (x"c8",x"0f",x"00",x"00"),
   735 => (x"18",x"10",x"27",x"86"),
   736 => (x"4a",x"bf",x"00",x"00"),
   737 => (x"1e",x"6a",x"82",x"c8"),
   738 => (x"00",x"14",x"80",x"27"),
   739 => (x"3d",x"27",x"1e",x"00"),
   740 => (x"0f",x"00",x"00",x"03"),
   741 => (x"1e",x"c2",x"86",x"c8"),
   742 => (x"00",x"14",x"99",x"27"),
   743 => (x"3d",x"27",x"1e",x"00"),
   744 => (x"0f",x"00",x"00",x"03"),
   745 => (x"10",x"27",x"86",x"c8"),
   746 => (x"bf",x"00",x"00",x"18"),
   747 => (x"6a",x"82",x"cc",x"4a"),
   748 => (x"14",x"b2",x"27",x"1e"),
   749 => (x"27",x"1e",x"00",x"00"),
   750 => (x"00",x"00",x"03",x"3d"),
   751 => (x"d1",x"86",x"c8",x"0f"),
   752 => (x"14",x"cb",x"27",x"1e"),
   753 => (x"27",x"1e",x"00",x"00"),
   754 => (x"00",x"00",x"03",x"3d"),
   755 => (x"27",x"86",x"c8",x"0f"),
   756 => (x"00",x"00",x"18",x"10"),
   757 => (x"82",x"d0",x"4a",x"bf"),
   758 => (x"e4",x"27",x"1e",x"72"),
   759 => (x"1e",x"00",x"00",x"14"),
   760 => (x"00",x"03",x"3d",x"27"),
   761 => (x"86",x"c8",x"0f",x"00"),
   762 => (x"00",x"14",x"fd",x"27"),
   763 => (x"3d",x"27",x"1e",x"00"),
   764 => (x"0f",x"00",x"00",x"03"),
   765 => (x"32",x"27",x"86",x"c4"),
   766 => (x"1e",x"00",x"00",x"15"),
   767 => (x"00",x"03",x"3d",x"27"),
   768 => (x"86",x"c4",x"0f",x"00"),
   769 => (x"00",x"18",x"14",x"27"),
   770 => (x"1e",x"bf",x"bf",x"00"),
   771 => (x"00",x"15",x"43",x"27"),
   772 => (x"3d",x"27",x"1e",x"00"),
   773 => (x"0f",x"00",x"00",x"03"),
   774 => (x"5c",x"27",x"86",x"c8"),
   775 => (x"1e",x"00",x"00",x"15"),
   776 => (x"00",x"03",x"3d",x"27"),
   777 => (x"86",x"c4",x"0f",x"00"),
   778 => (x"00",x"18",x"14",x"27"),
   779 => (x"c4",x"4a",x"bf",x"00"),
   780 => (x"27",x"1e",x"6a",x"82"),
   781 => (x"00",x"00",x"15",x"9c"),
   782 => (x"03",x"3d",x"27",x"1e"),
   783 => (x"c8",x"0f",x"00",x"00"),
   784 => (x"27",x"1e",x"c0",x"86"),
   785 => (x"00",x"00",x"15",x"b5"),
   786 => (x"03",x"3d",x"27",x"1e"),
   787 => (x"c8",x"0f",x"00",x"00"),
   788 => (x"18",x"14",x"27",x"86"),
   789 => (x"4a",x"bf",x"00",x"00"),
   790 => (x"1e",x"6a",x"82",x"c8"),
   791 => (x"00",x"15",x"ce",x"27"),
   792 => (x"3d",x"27",x"1e",x"00"),
   793 => (x"0f",x"00",x"00",x"03"),
   794 => (x"1e",x"c1",x"86",x"c8"),
   795 => (x"00",x"15",x"e7",x"27"),
   796 => (x"3d",x"27",x"1e",x"00"),
   797 => (x"0f",x"00",x"00",x"03"),
   798 => (x"14",x"27",x"86",x"c8"),
   799 => (x"bf",x"00",x"00",x"18"),
   800 => (x"6a",x"82",x"cc",x"4a"),
   801 => (x"16",x"00",x"27",x"1e"),
   802 => (x"27",x"1e",x"00",x"00"),
   803 => (x"00",x"00",x"03",x"3d"),
   804 => (x"d2",x"86",x"c8",x"0f"),
   805 => (x"16",x"19",x"27",x"1e"),
   806 => (x"27",x"1e",x"00",x"00"),
   807 => (x"00",x"00",x"03",x"3d"),
   808 => (x"27",x"86",x"c8",x"0f"),
   809 => (x"00",x"00",x"18",x"14"),
   810 => (x"82",x"d0",x"4a",x"bf"),
   811 => (x"32",x"27",x"1e",x"72"),
   812 => (x"1e",x"00",x"00",x"16"),
   813 => (x"00",x"03",x"3d",x"27"),
   814 => (x"86",x"c8",x"0f",x"00"),
   815 => (x"00",x"16",x"4b",x"27"),
   816 => (x"3d",x"27",x"1e",x"00"),
   817 => (x"0f",x"00",x"00",x"03"),
   818 => (x"1e",x"6e",x"86",x"c4"),
   819 => (x"00",x"16",x"80",x"27"),
   820 => (x"3d",x"27",x"1e",x"00"),
   821 => (x"0f",x"00",x"00",x"03"),
   822 => (x"1e",x"c5",x"86",x"c8"),
   823 => (x"00",x"16",x"99",x"27"),
   824 => (x"3d",x"27",x"1e",x"00"),
   825 => (x"0f",x"00",x"00",x"03"),
   826 => (x"1e",x"74",x"86",x"c8"),
   827 => (x"00",x"16",x"b2",x"27"),
   828 => (x"3d",x"27",x"1e",x"00"),
   829 => (x"0f",x"00",x"00",x"03"),
   830 => (x"1e",x"cd",x"86",x"c8"),
   831 => (x"00",x"16",x"cb",x"27"),
   832 => (x"3d",x"27",x"1e",x"00"),
   833 => (x"0f",x"00",x"00",x"03"),
   834 => (x"66",x"cc",x"86",x"c8"),
   835 => (x"16",x"e4",x"27",x"1e"),
   836 => (x"27",x"1e",x"00",x"00"),
   837 => (x"00",x"00",x"03",x"3d"),
   838 => (x"c7",x"86",x"c8",x"0f"),
   839 => (x"16",x"fd",x"27",x"1e"),
   840 => (x"27",x"1e",x"00",x"00"),
   841 => (x"00",x"00",x"03",x"3d"),
   842 => (x"c8",x"86",x"c8",x"0f"),
   843 => (x"16",x"27",x"1e",x"66"),
   844 => (x"1e",x"00",x"00",x"17"),
   845 => (x"00",x"03",x"3d",x"27"),
   846 => (x"86",x"c8",x"0f",x"00"),
   847 => (x"2f",x"27",x"1e",x"c1"),
   848 => (x"1e",x"00",x"00",x"17"),
   849 => (x"00",x"03",x"3d",x"27"),
   850 => (x"86",x"c8",x"0f",x"00"),
   851 => (x"00",x"40",x"78",x"27"),
   852 => (x"48",x"27",x"1e",x"00"),
   853 => (x"1e",x"00",x"00",x"17"),
   854 => (x"00",x"03",x"3d",x"27"),
   855 => (x"86",x"c8",x"0f",x"00"),
   856 => (x"00",x"17",x"61",x"27"),
   857 => (x"3d",x"27",x"1e",x"00"),
   858 => (x"0f",x"00",x"00",x"03"),
   859 => (x"98",x"27",x"86",x"c4"),
   860 => (x"1e",x"00",x"00",x"40"),
   861 => (x"00",x"17",x"96",x"27"),
   862 => (x"3d",x"27",x"1e",x"00"),
   863 => (x"0f",x"00",x"00",x"03"),
   864 => (x"af",x"27",x"86",x"c8"),
   865 => (x"1e",x"00",x"00",x"17"),
   866 => (x"00",x"03",x"3d",x"27"),
   867 => (x"86",x"c4",x"0f",x"00"),
   868 => (x"00",x"17",x"e4",x"27"),
   869 => (x"3d",x"27",x"1e",x"00"),
   870 => (x"0f",x"00",x"00",x"03"),
   871 => (x"04",x"27",x"86",x"c4"),
   872 => (x"bf",x"00",x"00",x"40"),
   873 => (x"40",x"00",x"27",x"4a"),
   874 => (x"8a",x"bf",x"00",x"00"),
   875 => (x"00",x"40",x"08",x"27"),
   876 => (x"79",x"72",x"49",x"00"),
   877 => (x"e6",x"27",x"1e",x"72"),
   878 => (x"1e",x"00",x"00",x"17"),
   879 => (x"00",x"03",x"3d",x"27"),
   880 => (x"86",x"c8",x"0f",x"00"),
   881 => (x"00",x"40",x"08",x"27"),
   882 => (x"c1",x"49",x"bf",x"00"),
   883 => (x"03",x"a9",x"b7",x"f8"),
   884 => (x"27",x"87",x"ea",x"c0"),
   885 => (x"00",x"00",x"10",x"f6"),
   886 => (x"03",x"3d",x"27",x"1e"),
   887 => (x"c4",x"0f",x"00",x"00"),
   888 => (x"11",x"2c",x"27",x"86"),
   889 => (x"27",x"1e",x"00",x"00"),
   890 => (x"00",x"00",x"03",x"3d"),
   891 => (x"27",x"86",x"c4",x"0f"),
   892 => (x"00",x"00",x"11",x"4c"),
   893 => (x"03",x"3d",x"27",x"1e"),
   894 => (x"c4",x"0f",x"00",x"00"),
   895 => (x"40",x"08",x"27",x"86"),
   896 => (x"4a",x"bf",x"00",x"00"),
   897 => (x"e8",x"cf",x"4b",x"72"),
   898 => (x"72",x"49",x"73",x"93"),
   899 => (x"17",x"fc",x"27",x"1e"),
   900 => (x"4a",x"bf",x"00",x"00"),
   901 => (x"00",x"06",x"b0",x"27"),
   902 => (x"4a",x"26",x"0f",x"00"),
   903 => (x"10",x"27",x"48",x"70"),
   904 => (x"58",x"00",x"00",x"40"),
   905 => (x"00",x"17",x"fc",x"27"),
   906 => (x"73",x"4b",x"bf",x"00"),
   907 => (x"94",x"e8",x"cf",x"4c"),
   908 => (x"1e",x"72",x"49",x"74"),
   909 => (x"b0",x"27",x"4a",x"72"),
   910 => (x"0f",x"00",x"00",x"06"),
   911 => (x"48",x"70",x"4a",x"26"),
   912 => (x"00",x"40",x"14",x"27"),
   913 => (x"f9",x"c8",x"58",x"00"),
   914 => (x"72",x"49",x"73",x"93"),
   915 => (x"27",x"4a",x"72",x"1e"),
   916 => (x"00",x"00",x"06",x"b0"),
   917 => (x"70",x"4a",x"26",x"0f"),
   918 => (x"40",x"18",x"27",x"48"),
   919 => (x"27",x"58",x"00",x"00"),
   920 => (x"00",x"00",x"11",x"4e"),
   921 => (x"03",x"3d",x"27",x"1e"),
   922 => (x"c4",x"0f",x"00",x"00"),
   923 => (x"40",x"0c",x"27",x"86"),
   924 => (x"1e",x"bf",x"00",x"00"),
   925 => (x"00",x"11",x"7b",x"27"),
   926 => (x"3d",x"27",x"1e",x"00"),
   927 => (x"0f",x"00",x"00",x"03"),
   928 => (x"80",x"27",x"86",x"c8"),
   929 => (x"1e",x"00",x"00",x"11"),
   930 => (x"00",x"03",x"3d",x"27"),
   931 => (x"86",x"c4",x"0f",x"00"),
   932 => (x"00",x"40",x"10",x"27"),
   933 => (x"27",x"1e",x"bf",x"00"),
   934 => (x"00",x"00",x"11",x"ad"),
   935 => (x"03",x"3d",x"27",x"1e"),
   936 => (x"c8",x"0f",x"00",x"00"),
   937 => (x"40",x"14",x"27",x"86"),
   938 => (x"1e",x"bf",x"00",x"00"),
   939 => (x"00",x"11",x"b2",x"27"),
   940 => (x"3d",x"27",x"1e",x"00"),
   941 => (x"0f",x"00",x"00",x"03"),
   942 => (x"d0",x"27",x"86",x"c8"),
   943 => (x"1e",x"00",x"00",x"11"),
   944 => (x"00",x"03",x"3d",x"27"),
   945 => (x"86",x"c4",x"0f",x"00"),
   946 => (x"86",x"d0",x"48",x"c0"),
   947 => (x"4c",x"26",x"4d",x"26"),
   948 => (x"4a",x"26",x"4b",x"26"),
   949 => (x"5e",x"0e",x"4f",x"26"),
   950 => (x"5d",x"5c",x"5b",x"5a"),
   951 => (x"bf",x"66",x"d4",x"0e"),
   952 => (x"27",x"4d",x"72",x"4a"),
   953 => (x"00",x"00",x"18",x"10"),
   954 => (x"1e",x"72",x"48",x"bf"),
   955 => (x"49",x"a2",x"f0",x"c0"),
   956 => (x"a9",x"72",x"42",x"20"),
   957 => (x"26",x"87",x"f9",x"05"),
   958 => (x"4c",x"66",x"d4",x"4a"),
   959 => (x"7c",x"c5",x"84",x"cc"),
   960 => (x"83",x"cc",x"4b",x"72"),
   961 => (x"66",x"d4",x"7b",x"6c"),
   962 => (x"1e",x"72",x"7a",x"bf"),
   963 => (x"00",x"0f",x"bb",x"27"),
   964 => (x"86",x"c4",x"0f",x"00"),
   965 => (x"05",x"6a",x"82",x"c4"),
   966 => (x"75",x"87",x"f4",x"c0"),
   967 => (x"75",x"83",x"c8",x"4b"),
   968 => (x"c6",x"82",x"cc",x"4a"),
   969 => (x"d8",x"1e",x"73",x"7a"),
   970 => (x"83",x"c8",x"4b",x"66"),
   971 => (x"3b",x"27",x"1e",x"6b"),
   972 => (x"0f",x"00",x"00",x"04"),
   973 => (x"10",x"27",x"86",x"c8"),
   974 => (x"bf",x"00",x"00",x"18"),
   975 => (x"1e",x"72",x"7d",x"bf"),
   976 => (x"1e",x"6a",x"1e",x"ca"),
   977 => (x"00",x"04",x"ad",x"27"),
   978 => (x"86",x"cc",x"0f",x"00"),
   979 => (x"d4",x"87",x"d7",x"c0"),
   980 => (x"d4",x"4a",x"bf",x"66"),
   981 => (x"72",x"48",x"49",x"66"),
   982 => (x"a1",x"f0",x"c0",x"1e"),
   983 => (x"71",x"41",x"20",x"4a"),
   984 => (x"87",x"f9",x"05",x"aa"),
   985 => (x"4d",x"26",x"4a",x"26"),
   986 => (x"4b",x"26",x"4c",x"26"),
   987 => (x"4f",x"26",x"4a",x"26"),
   988 => (x"5b",x"5a",x"5e",x"0e"),
   989 => (x"1e",x"0e",x"5d",x"5c"),
   990 => (x"66",x"d8",x"4d",x"6e"),
   991 => (x"ca",x"4b",x"6c",x"4c"),
   992 => (x"18",x"20",x"27",x"83"),
   993 => (x"bf",x"97",x"00",x"00"),
   994 => (x"c0",x"c0",x"c1",x"4a"),
   995 => (x"c4",x"92",x"c0",x"c0"),
   996 => (x"4a",x"92",x"b7",x"c0"),
   997 => (x"05",x"aa",x"c1",x"c1"),
   998 => (x"c1",x"87",x"cf",x"c0"),
   999 => (x"27",x"48",x"73",x"8b"),
  1000 => (x"00",x"00",x"18",x"18"),
  1001 => (x"7c",x"70",x"88",x"bf"),
  1002 => (x"9d",x"75",x"4d",x"c0"),
  1003 => (x"87",x"d1",x"ff",x"05"),
  1004 => (x"26",x"4d",x"26",x"26"),
  1005 => (x"26",x"4b",x"26",x"4c"),
  1006 => (x"1e",x"4f",x"26",x"4a"),
  1007 => (x"10",x"27",x"1e",x"72"),
  1008 => (x"bf",x"00",x"00",x"18"),
  1009 => (x"87",x"cb",x"c0",x"02"),
  1010 => (x"27",x"49",x"66",x"c8"),
  1011 => (x"00",x"00",x"18",x"10"),
  1012 => (x"27",x"79",x"bf",x"bf"),
  1013 => (x"00",x"00",x"18",x"10"),
  1014 => (x"82",x"cc",x"4a",x"bf"),
  1015 => (x"18",x"27",x"1e",x"72"),
  1016 => (x"bf",x"00",x"00",x"18"),
  1017 => (x"27",x"1e",x"ca",x"1e"),
  1018 => (x"00",x"00",x"04",x"ad"),
  1019 => (x"26",x"86",x"cc",x"0f"),
  1020 => (x"1e",x"4f",x"26",x"4a"),
  1021 => (x"20",x"27",x"1e",x"72"),
  1022 => (x"97",x"00",x"00",x"18"),
  1023 => (x"c0",x"c1",x"4a",x"bf"),
  1024 => (x"92",x"c0",x"c0",x"c0"),
  1025 => (x"92",x"b7",x"c0",x"c4"),
  1026 => (x"aa",x"c1",x"c1",x"4a"),
  1027 => (x"87",x"c5",x"c0",x"02"),
  1028 => (x"c2",x"c0",x"4a",x"c0"),
  1029 => (x"27",x"4a",x"c1",x"87"),
  1030 => (x"00",x"00",x"18",x"1c"),
  1031 => (x"b0",x"72",x"48",x"bf"),
  1032 => (x"00",x"18",x"20",x"27"),
  1033 => (x"21",x"27",x"58",x"00"),
  1034 => (x"49",x"00",x"00",x"18"),
  1035 => (x"26",x"51",x"c2",x"c1"),
  1036 => (x"1e",x"4f",x"26",x"4a"),
  1037 => (x"00",x"18",x"20",x"27"),
  1038 => (x"c1",x"c1",x"49",x"00"),
  1039 => (x"18",x"1c",x"27",x"51"),
  1040 => (x"c0",x"49",x"00",x"00"),
  1041 => (x"00",x"4f",x"26",x"79"),
  1042 => (x"33",x"32",x"31",x"30"),
  1043 => (x"37",x"36",x"35",x"34"),
  1044 => (x"42",x"41",x"39",x"38"),
  1045 => (x"46",x"45",x"44",x"43"),
  1046 => (x"6f",x"72",x"50",x"00"),
  1047 => (x"6d",x"61",x"72",x"67"),
  1048 => (x"6d",x"6f",x"63",x"20"),
  1049 => (x"65",x"6c",x"69",x"70"),
  1050 => (x"69",x"77",x"20",x"64"),
  1051 => (x"27",x"20",x"68",x"74"),
  1052 => (x"69",x"67",x"65",x"72"),
  1053 => (x"72",x"65",x"74",x"73"),
  1054 => (x"74",x"61",x"20",x"27"),
  1055 => (x"62",x"69",x"72",x"74"),
  1056 => (x"0a",x"65",x"74",x"75"),
  1057 => (x"50",x"00",x"0a",x"00"),
  1058 => (x"72",x"67",x"6f",x"72"),
  1059 => (x"63",x"20",x"6d",x"61"),
  1060 => (x"69",x"70",x"6d",x"6f"),
  1061 => (x"20",x"64",x"65",x"6c"),
  1062 => (x"68",x"74",x"69",x"77"),
  1063 => (x"20",x"74",x"75",x"6f"),
  1064 => (x"67",x"65",x"72",x"27"),
  1065 => (x"65",x"74",x"73",x"69"),
  1066 => (x"61",x"20",x"27",x"72"),
  1067 => (x"69",x"72",x"74",x"74"),
  1068 => (x"65",x"74",x"75",x"62"),
  1069 => (x"00",x"0a",x"00",x"0a"),
  1070 => (x"59",x"52",x"48",x"44"),
  1071 => (x"4e",x"4f",x"54",x"53"),
  1072 => (x"52",x"50",x"20",x"45"),
  1073 => (x"41",x"52",x"47",x"4f"),
  1074 => (x"33",x"20",x"2c",x"4d"),
  1075 => (x"20",x"44",x"52",x"27"),
  1076 => (x"49",x"52",x"54",x"53"),
  1077 => (x"44",x"00",x"47",x"4e"),
  1078 => (x"53",x"59",x"52",x"48"),
  1079 => (x"45",x"4e",x"4f",x"54"),
  1080 => (x"4f",x"52",x"50",x"20"),
  1081 => (x"4d",x"41",x"52",x"47"),
  1082 => (x"27",x"32",x"20",x"2c"),
  1083 => (x"53",x"20",x"44",x"4e"),
  1084 => (x"4e",x"49",x"52",x"54"),
  1085 => (x"65",x"4d",x"00",x"47"),
  1086 => (x"72",x"75",x"73",x"61"),
  1087 => (x"74",x"20",x"64",x"65"),
  1088 => (x"20",x"65",x"6d",x"69"),
  1089 => (x"20",x"6f",x"6f",x"74"),
  1090 => (x"6c",x"61",x"6d",x"73"),
  1091 => (x"6f",x"74",x"20",x"6c"),
  1092 => (x"74",x"62",x"6f",x"20"),
  1093 => (x"20",x"6e",x"69",x"61"),
  1094 => (x"6e",x"61",x"65",x"6d"),
  1095 => (x"66",x"67",x"6e",x"69"),
  1096 => (x"72",x"20",x"6c",x"75"),
  1097 => (x"6c",x"75",x"73",x"65"),
  1098 => (x"00",x"0a",x"73",x"74"),
  1099 => (x"61",x"65",x"6c",x"50"),
  1100 => (x"69",x"20",x"65",x"73"),
  1101 => (x"65",x"72",x"63",x"6e"),
  1102 => (x"20",x"65",x"73",x"61"),
  1103 => (x"62",x"6d",x"75",x"6e"),
  1104 => (x"6f",x"20",x"72",x"65"),
  1105 => (x"75",x"72",x"20",x"66"),
  1106 => (x"00",x"0a",x"73",x"6e"),
  1107 => (x"69",x"4d",x"00",x"0a"),
  1108 => (x"73",x"6f",x"72",x"63"),
  1109 => (x"6e",x"6f",x"63",x"65"),
  1110 => (x"66",x"20",x"73",x"64"),
  1111 => (x"6f",x"20",x"72",x"6f"),
  1112 => (x"72",x"20",x"65",x"6e"),
  1113 => (x"74",x"20",x"6e",x"75"),
  1114 => (x"75",x"6f",x"72",x"68"),
  1115 => (x"44",x"20",x"68",x"67"),
  1116 => (x"73",x"79",x"72",x"68"),
  1117 => (x"65",x"6e",x"6f",x"74"),
  1118 => (x"25",x"00",x"20",x"3a"),
  1119 => (x"00",x"0a",x"20",x"64"),
  1120 => (x"79",x"72",x"68",x"44"),
  1121 => (x"6e",x"6f",x"74",x"73"),
  1122 => (x"70",x"20",x"73",x"65"),
  1123 => (x"53",x"20",x"72",x"65"),
  1124 => (x"6e",x"6f",x"63",x"65"),
  1125 => (x"20",x"20",x"3a",x"64"),
  1126 => (x"20",x"20",x"20",x"20"),
  1127 => (x"20",x"20",x"20",x"20"),
  1128 => (x"20",x"20",x"20",x"20"),
  1129 => (x"20",x"20",x"20",x"20"),
  1130 => (x"20",x"20",x"20",x"20"),
  1131 => (x"20",x"64",x"25",x"00"),
  1132 => (x"41",x"56",x"00",x"0a"),
  1133 => (x"49",x"4d",x"20",x"58"),
  1134 => (x"72",x"20",x"53",x"50"),
  1135 => (x"6e",x"69",x"74",x"61"),
  1136 => (x"20",x"2a",x"20",x"67"),
  1137 => (x"30",x"30",x"30",x"31"),
  1138 => (x"25",x"20",x"3d",x"20"),
  1139 => (x"00",x"0a",x"20",x"64"),
  1140 => (x"48",x"44",x"00",x"0a"),
  1141 => (x"54",x"53",x"59",x"52"),
  1142 => (x"20",x"45",x"4e",x"4f"),
  1143 => (x"47",x"4f",x"52",x"50"),
  1144 => (x"2c",x"4d",x"41",x"52"),
  1145 => (x"4d",x"4f",x"53",x"20"),
  1146 => (x"54",x"53",x"20",x"45"),
  1147 => (x"47",x"4e",x"49",x"52"),
  1148 => (x"52",x"48",x"44",x"00"),
  1149 => (x"4f",x"54",x"53",x"59"),
  1150 => (x"50",x"20",x"45",x"4e"),
  1151 => (x"52",x"47",x"4f",x"52"),
  1152 => (x"20",x"2c",x"4d",x"41"),
  1153 => (x"54",x"53",x"27",x"31"),
  1154 => (x"52",x"54",x"53",x"20"),
  1155 => (x"00",x"47",x"4e",x"49"),
  1156 => (x"68",x"44",x"00",x"0a"),
  1157 => (x"74",x"73",x"79",x"72"),
  1158 => (x"20",x"65",x"6e",x"6f"),
  1159 => (x"63",x"6e",x"65",x"42"),
  1160 => (x"72",x"61",x"6d",x"68"),
  1161 => (x"56",x"20",x"2c",x"6b"),
  1162 => (x"69",x"73",x"72",x"65"),
  1163 => (x"32",x"20",x"6e",x"6f"),
  1164 => (x"28",x"20",x"31",x"2e"),
  1165 => (x"67",x"6e",x"61",x"4c"),
  1166 => (x"65",x"67",x"61",x"75"),
  1167 => (x"29",x"43",x"20",x"3a"),
  1168 => (x"00",x"0a",x"00",x"0a"),
  1169 => (x"63",x"65",x"78",x"45"),
  1170 => (x"6f",x"69",x"74",x"75"),
  1171 => (x"74",x"73",x"20",x"6e"),
  1172 => (x"73",x"74",x"72",x"61"),
  1173 => (x"64",x"25",x"20",x"2c"),
  1174 => (x"6e",x"75",x"72",x"20"),
  1175 => (x"68",x"74",x"20",x"73"),
  1176 => (x"67",x"75",x"6f",x"72"),
  1177 => (x"68",x"44",x"20",x"68"),
  1178 => (x"74",x"73",x"79",x"72"),
  1179 => (x"0a",x"65",x"6e",x"6f"),
  1180 => (x"65",x"78",x"45",x"00"),
  1181 => (x"69",x"74",x"75",x"63"),
  1182 => (x"65",x"20",x"6e",x"6f"),
  1183 => (x"0a",x"73",x"64",x"6e"),
  1184 => (x"46",x"00",x"0a",x"00"),
  1185 => (x"6c",x"61",x"6e",x"69"),
  1186 => (x"6c",x"61",x"76",x"20"),
  1187 => (x"20",x"73",x"65",x"75"),
  1188 => (x"74",x"20",x"66",x"6f"),
  1189 => (x"76",x"20",x"65",x"68"),
  1190 => (x"61",x"69",x"72",x"61"),
  1191 => (x"73",x"65",x"6c",x"62"),
  1192 => (x"65",x"73",x"75",x"20"),
  1193 => (x"6e",x"69",x"20",x"64"),
  1194 => (x"65",x"68",x"74",x"20"),
  1195 => (x"6e",x"65",x"62",x"20"),
  1196 => (x"61",x"6d",x"68",x"63"),
  1197 => (x"0a",x"3a",x"6b",x"72"),
  1198 => (x"49",x"00",x"0a",x"00"),
  1199 => (x"47",x"5f",x"74",x"6e"),
  1200 => (x"3a",x"62",x"6f",x"6c"),
  1201 => (x"20",x"20",x"20",x"20"),
  1202 => (x"20",x"20",x"20",x"20"),
  1203 => (x"20",x"20",x"20",x"20"),
  1204 => (x"00",x"0a",x"64",x"25"),
  1205 => (x"20",x"20",x"20",x"20"),
  1206 => (x"20",x"20",x"20",x"20"),
  1207 => (x"75",x"6f",x"68",x"73"),
  1208 => (x"62",x"20",x"64",x"6c"),
  1209 => (x"20",x"20",x"3a",x"65"),
  1210 => (x"0a",x"64",x"25",x"20"),
  1211 => (x"6f",x"6f",x"42",x"00"),
  1212 => (x"6c",x"47",x"5f",x"6c"),
  1213 => (x"20",x"3a",x"62",x"6f"),
  1214 => (x"20",x"20",x"20",x"20"),
  1215 => (x"20",x"20",x"20",x"20"),
  1216 => (x"64",x"25",x"20",x"20"),
  1217 => (x"20",x"20",x"00",x"0a"),
  1218 => (x"20",x"20",x"20",x"20"),
  1219 => (x"68",x"73",x"20",x"20"),
  1220 => (x"64",x"6c",x"75",x"6f"),
  1221 => (x"3a",x"65",x"62",x"20"),
  1222 => (x"25",x"20",x"20",x"20"),
  1223 => (x"43",x"00",x"0a",x"64"),
  1224 => (x"5f",x"31",x"5f",x"68"),
  1225 => (x"62",x"6f",x"6c",x"47"),
  1226 => (x"20",x"20",x"20",x"3a"),
  1227 => (x"20",x"20",x"20",x"20"),
  1228 => (x"20",x"20",x"20",x"20"),
  1229 => (x"00",x"0a",x"63",x"25"),
  1230 => (x"20",x"20",x"20",x"20"),
  1231 => (x"20",x"20",x"20",x"20"),
  1232 => (x"75",x"6f",x"68",x"73"),
  1233 => (x"62",x"20",x"64",x"6c"),
  1234 => (x"20",x"20",x"3a",x"65"),
  1235 => (x"0a",x"63",x"25",x"20"),
  1236 => (x"5f",x"68",x"43",x"00"),
  1237 => (x"6c",x"47",x"5f",x"32"),
  1238 => (x"20",x"3a",x"62",x"6f"),
  1239 => (x"20",x"20",x"20",x"20"),
  1240 => (x"20",x"20",x"20",x"20"),
  1241 => (x"63",x"25",x"20",x"20"),
  1242 => (x"20",x"20",x"00",x"0a"),
  1243 => (x"20",x"20",x"20",x"20"),
  1244 => (x"68",x"73",x"20",x"20"),
  1245 => (x"64",x"6c",x"75",x"6f"),
  1246 => (x"3a",x"65",x"62",x"20"),
  1247 => (x"25",x"20",x"20",x"20"),
  1248 => (x"41",x"00",x"0a",x"63"),
  1249 => (x"31",x"5f",x"72",x"72"),
  1250 => (x"6f",x"6c",x"47",x"5f"),
  1251 => (x"5d",x"38",x"5b",x"62"),
  1252 => (x"20",x"20",x"20",x"3a"),
  1253 => (x"20",x"20",x"20",x"20"),
  1254 => (x"00",x"0a",x"64",x"25"),
  1255 => (x"20",x"20",x"20",x"20"),
  1256 => (x"20",x"20",x"20",x"20"),
  1257 => (x"75",x"6f",x"68",x"73"),
  1258 => (x"62",x"20",x"64",x"6c"),
  1259 => (x"20",x"20",x"3a",x"65"),
  1260 => (x"0a",x"64",x"25",x"20"),
  1261 => (x"72",x"72",x"41",x"00"),
  1262 => (x"47",x"5f",x"32",x"5f"),
  1263 => (x"5b",x"62",x"6f",x"6c"),
  1264 => (x"37",x"5b",x"5d",x"38"),
  1265 => (x"20",x"20",x"3a",x"5d"),
  1266 => (x"64",x"25",x"20",x"20"),
  1267 => (x"20",x"20",x"00",x"0a"),
  1268 => (x"20",x"20",x"20",x"20"),
  1269 => (x"68",x"73",x"20",x"20"),
  1270 => (x"64",x"6c",x"75",x"6f"),
  1271 => (x"3a",x"65",x"62",x"20"),
  1272 => (x"4e",x"20",x"20",x"20"),
  1273 => (x"65",x"62",x"6d",x"75"),
  1274 => (x"66",x"4f",x"5f",x"72"),
  1275 => (x"6e",x"75",x"52",x"5f"),
  1276 => (x"20",x"2b",x"20",x"73"),
  1277 => (x"00",x"0a",x"30",x"31"),
  1278 => (x"5f",x"72",x"74",x"50"),
  1279 => (x"62",x"6f",x"6c",x"47"),
  1280 => (x"00",x"0a",x"3e",x"2d"),
  1281 => (x"74",x"50",x"20",x"20"),
  1282 => (x"6f",x"43",x"5f",x"72"),
  1283 => (x"20",x"3a",x"70",x"6d"),
  1284 => (x"20",x"20",x"20",x"20"),
  1285 => (x"20",x"20",x"20",x"20"),
  1286 => (x"0a",x"64",x"25",x"20"),
  1287 => (x"20",x"20",x"20",x"00"),
  1288 => (x"20",x"20",x"20",x"20"),
  1289 => (x"6f",x"68",x"73",x"20"),
  1290 => (x"20",x"64",x"6c",x"75"),
  1291 => (x"20",x"3a",x"65",x"62"),
  1292 => (x"69",x"28",x"20",x"20"),
  1293 => (x"65",x"6c",x"70",x"6d"),
  1294 => (x"74",x"6e",x"65",x"6d"),
  1295 => (x"6f",x"69",x"74",x"61"),
  1296 => (x"65",x"64",x"2d",x"6e"),
  1297 => (x"64",x"6e",x"65",x"70"),
  1298 => (x"29",x"74",x"6e",x"65"),
  1299 => (x"20",x"20",x"00",x"0a"),
  1300 => (x"63",x"73",x"69",x"44"),
  1301 => (x"20",x"20",x"3a",x"72"),
  1302 => (x"20",x"20",x"20",x"20"),
  1303 => (x"20",x"20",x"20",x"20"),
  1304 => (x"25",x"20",x"20",x"20"),
  1305 => (x"20",x"00",x"0a",x"64"),
  1306 => (x"20",x"20",x"20",x"20"),
  1307 => (x"73",x"20",x"20",x"20"),
  1308 => (x"6c",x"75",x"6f",x"68"),
  1309 => (x"65",x"62",x"20",x"64"),
  1310 => (x"20",x"20",x"20",x"3a"),
  1311 => (x"00",x"0a",x"64",x"25"),
  1312 => (x"6e",x"45",x"20",x"20"),
  1313 => (x"43",x"5f",x"6d",x"75"),
  1314 => (x"3a",x"70",x"6d",x"6f"),
  1315 => (x"20",x"20",x"20",x"20"),
  1316 => (x"20",x"20",x"20",x"20"),
  1317 => (x"0a",x"64",x"25",x"20"),
  1318 => (x"20",x"20",x"20",x"00"),
  1319 => (x"20",x"20",x"20",x"20"),
  1320 => (x"6f",x"68",x"73",x"20"),
  1321 => (x"20",x"64",x"6c",x"75"),
  1322 => (x"20",x"3a",x"65",x"62"),
  1323 => (x"64",x"25",x"20",x"20"),
  1324 => (x"20",x"20",x"00",x"0a"),
  1325 => (x"5f",x"74",x"6e",x"49"),
  1326 => (x"70",x"6d",x"6f",x"43"),
  1327 => (x"20",x"20",x"20",x"3a"),
  1328 => (x"20",x"20",x"20",x"20"),
  1329 => (x"25",x"20",x"20",x"20"),
  1330 => (x"20",x"00",x"0a",x"64"),
  1331 => (x"20",x"20",x"20",x"20"),
  1332 => (x"73",x"20",x"20",x"20"),
  1333 => (x"6c",x"75",x"6f",x"68"),
  1334 => (x"65",x"62",x"20",x"64"),
  1335 => (x"20",x"20",x"20",x"3a"),
  1336 => (x"00",x"0a",x"64",x"25"),
  1337 => (x"74",x"53",x"20",x"20"),
  1338 => (x"6f",x"43",x"5f",x"72"),
  1339 => (x"20",x"3a",x"70",x"6d"),
  1340 => (x"20",x"20",x"20",x"20"),
  1341 => (x"20",x"20",x"20",x"20"),
  1342 => (x"0a",x"73",x"25",x"20"),
  1343 => (x"20",x"20",x"20",x"00"),
  1344 => (x"20",x"20",x"20",x"20"),
  1345 => (x"6f",x"68",x"73",x"20"),
  1346 => (x"20",x"64",x"6c",x"75"),
  1347 => (x"20",x"3a",x"65",x"62"),
  1348 => (x"48",x"44",x"20",x"20"),
  1349 => (x"54",x"53",x"59",x"52"),
  1350 => (x"20",x"45",x"4e",x"4f"),
  1351 => (x"47",x"4f",x"52",x"50"),
  1352 => (x"2c",x"4d",x"41",x"52"),
  1353 => (x"4d",x"4f",x"53",x"20"),
  1354 => (x"54",x"53",x"20",x"45"),
  1355 => (x"47",x"4e",x"49",x"52"),
  1356 => (x"65",x"4e",x"00",x"0a"),
  1357 => (x"50",x"5f",x"74",x"78"),
  1358 => (x"47",x"5f",x"72",x"74"),
  1359 => (x"2d",x"62",x"6f",x"6c"),
  1360 => (x"20",x"00",x"0a",x"3e"),
  1361 => (x"72",x"74",x"50",x"20"),
  1362 => (x"6d",x"6f",x"43",x"5f"),
  1363 => (x"20",x"20",x"3a",x"70"),
  1364 => (x"20",x"20",x"20",x"20"),
  1365 => (x"20",x"20",x"20",x"20"),
  1366 => (x"00",x"0a",x"64",x"25"),
  1367 => (x"20",x"20",x"20",x"20"),
  1368 => (x"20",x"20",x"20",x"20"),
  1369 => (x"75",x"6f",x"68",x"73"),
  1370 => (x"62",x"20",x"64",x"6c"),
  1371 => (x"20",x"20",x"3a",x"65"),
  1372 => (x"6d",x"69",x"28",x"20"),
  1373 => (x"6d",x"65",x"6c",x"70"),
  1374 => (x"61",x"74",x"6e",x"65"),
  1375 => (x"6e",x"6f",x"69",x"74"),
  1376 => (x"70",x"65",x"64",x"2d"),
  1377 => (x"65",x"64",x"6e",x"65"),
  1378 => (x"2c",x"29",x"74",x"6e"),
  1379 => (x"6d",x"61",x"73",x"20"),
  1380 => (x"73",x"61",x"20",x"65"),
  1381 => (x"6f",x"62",x"61",x"20"),
  1382 => (x"00",x"0a",x"65",x"76"),
  1383 => (x"69",x"44",x"20",x"20"),
  1384 => (x"3a",x"72",x"63",x"73"),
  1385 => (x"20",x"20",x"20",x"20"),
  1386 => (x"20",x"20",x"20",x"20"),
  1387 => (x"20",x"20",x"20",x"20"),
  1388 => (x"0a",x"64",x"25",x"20"),
  1389 => (x"20",x"20",x"20",x"00"),
  1390 => (x"20",x"20",x"20",x"20"),
  1391 => (x"6f",x"68",x"73",x"20"),
  1392 => (x"20",x"64",x"6c",x"75"),
  1393 => (x"20",x"3a",x"65",x"62"),
  1394 => (x"64",x"25",x"20",x"20"),
  1395 => (x"20",x"20",x"00",x"0a"),
  1396 => (x"6d",x"75",x"6e",x"45"),
  1397 => (x"6d",x"6f",x"43",x"5f"),
  1398 => (x"20",x"20",x"3a",x"70"),
  1399 => (x"20",x"20",x"20",x"20"),
  1400 => (x"25",x"20",x"20",x"20"),
  1401 => (x"20",x"00",x"0a",x"64"),
  1402 => (x"20",x"20",x"20",x"20"),
  1403 => (x"73",x"20",x"20",x"20"),
  1404 => (x"6c",x"75",x"6f",x"68"),
  1405 => (x"65",x"62",x"20",x"64"),
  1406 => (x"20",x"20",x"20",x"3a"),
  1407 => (x"00",x"0a",x"64",x"25"),
  1408 => (x"6e",x"49",x"20",x"20"),
  1409 => (x"6f",x"43",x"5f",x"74"),
  1410 => (x"20",x"3a",x"70",x"6d"),
  1411 => (x"20",x"20",x"20",x"20"),
  1412 => (x"20",x"20",x"20",x"20"),
  1413 => (x"0a",x"64",x"25",x"20"),
  1414 => (x"20",x"20",x"20",x"00"),
  1415 => (x"20",x"20",x"20",x"20"),
  1416 => (x"6f",x"68",x"73",x"20"),
  1417 => (x"20",x"64",x"6c",x"75"),
  1418 => (x"20",x"3a",x"65",x"62"),
  1419 => (x"64",x"25",x"20",x"20"),
  1420 => (x"20",x"20",x"00",x"0a"),
  1421 => (x"5f",x"72",x"74",x"53"),
  1422 => (x"70",x"6d",x"6f",x"43"),
  1423 => (x"20",x"20",x"20",x"3a"),
  1424 => (x"20",x"20",x"20",x"20"),
  1425 => (x"25",x"20",x"20",x"20"),
  1426 => (x"20",x"00",x"0a",x"73"),
  1427 => (x"20",x"20",x"20",x"20"),
  1428 => (x"73",x"20",x"20",x"20"),
  1429 => (x"6c",x"75",x"6f",x"68"),
  1430 => (x"65",x"62",x"20",x"64"),
  1431 => (x"20",x"20",x"20",x"3a"),
  1432 => (x"59",x"52",x"48",x"44"),
  1433 => (x"4e",x"4f",x"54",x"53"),
  1434 => (x"52",x"50",x"20",x"45"),
  1435 => (x"41",x"52",x"47",x"4f"),
  1436 => (x"53",x"20",x"2c",x"4d"),
  1437 => (x"20",x"45",x"4d",x"4f"),
  1438 => (x"49",x"52",x"54",x"53"),
  1439 => (x"00",x"0a",x"47",x"4e"),
  1440 => (x"5f",x"74",x"6e",x"49"),
  1441 => (x"6f",x"4c",x"5f",x"31"),
  1442 => (x"20",x"20",x"3a",x"63"),
  1443 => (x"20",x"20",x"20",x"20"),
  1444 => (x"20",x"20",x"20",x"20"),
  1445 => (x"0a",x"64",x"25",x"20"),
  1446 => (x"20",x"20",x"20",x"00"),
  1447 => (x"20",x"20",x"20",x"20"),
  1448 => (x"6f",x"68",x"73",x"20"),
  1449 => (x"20",x"64",x"6c",x"75"),
  1450 => (x"20",x"3a",x"65",x"62"),
  1451 => (x"64",x"25",x"20",x"20"),
  1452 => (x"6e",x"49",x"00",x"0a"),
  1453 => (x"5f",x"32",x"5f",x"74"),
  1454 => (x"3a",x"63",x"6f",x"4c"),
  1455 => (x"20",x"20",x"20",x"20"),
  1456 => (x"20",x"20",x"20",x"20"),
  1457 => (x"25",x"20",x"20",x"20"),
  1458 => (x"20",x"00",x"0a",x"64"),
  1459 => (x"20",x"20",x"20",x"20"),
  1460 => (x"73",x"20",x"20",x"20"),
  1461 => (x"6c",x"75",x"6f",x"68"),
  1462 => (x"65",x"62",x"20",x"64"),
  1463 => (x"20",x"20",x"20",x"3a"),
  1464 => (x"00",x"0a",x"64",x"25"),
  1465 => (x"5f",x"74",x"6e",x"49"),
  1466 => (x"6f",x"4c",x"5f",x"33"),
  1467 => (x"20",x"20",x"3a",x"63"),
  1468 => (x"20",x"20",x"20",x"20"),
  1469 => (x"20",x"20",x"20",x"20"),
  1470 => (x"0a",x"64",x"25",x"20"),
  1471 => (x"20",x"20",x"20",x"00"),
  1472 => (x"20",x"20",x"20",x"20"),
  1473 => (x"6f",x"68",x"73",x"20"),
  1474 => (x"20",x"64",x"6c",x"75"),
  1475 => (x"20",x"3a",x"65",x"62"),
  1476 => (x"64",x"25",x"20",x"20"),
  1477 => (x"6e",x"45",x"00",x"0a"),
  1478 => (x"4c",x"5f",x"6d",x"75"),
  1479 => (x"20",x"3a",x"63",x"6f"),
  1480 => (x"20",x"20",x"20",x"20"),
  1481 => (x"20",x"20",x"20",x"20"),
  1482 => (x"25",x"20",x"20",x"20"),
  1483 => (x"20",x"00",x"0a",x"64"),
  1484 => (x"20",x"20",x"20",x"20"),
  1485 => (x"73",x"20",x"20",x"20"),
  1486 => (x"6c",x"75",x"6f",x"68"),
  1487 => (x"65",x"62",x"20",x"64"),
  1488 => (x"20",x"20",x"20",x"3a"),
  1489 => (x"00",x"0a",x"64",x"25"),
  1490 => (x"5f",x"72",x"74",x"53"),
  1491 => (x"6f",x"4c",x"5f",x"31"),
  1492 => (x"20",x"20",x"3a",x"63"),
  1493 => (x"20",x"20",x"20",x"20"),
  1494 => (x"20",x"20",x"20",x"20"),
  1495 => (x"0a",x"73",x"25",x"20"),
  1496 => (x"20",x"20",x"20",x"00"),
  1497 => (x"20",x"20",x"20",x"20"),
  1498 => (x"6f",x"68",x"73",x"20"),
  1499 => (x"20",x"64",x"6c",x"75"),
  1500 => (x"20",x"3a",x"65",x"62"),
  1501 => (x"48",x"44",x"20",x"20"),
  1502 => (x"54",x"53",x"59",x"52"),
  1503 => (x"20",x"45",x"4e",x"4f"),
  1504 => (x"47",x"4f",x"52",x"50"),
  1505 => (x"2c",x"4d",x"41",x"52"),
  1506 => (x"53",x"27",x"31",x"20"),
  1507 => (x"54",x"53",x"20",x"54"),
  1508 => (x"47",x"4e",x"49",x"52"),
  1509 => (x"74",x"53",x"00",x"0a"),
  1510 => (x"5f",x"32",x"5f",x"72"),
  1511 => (x"3a",x"63",x"6f",x"4c"),
  1512 => (x"20",x"20",x"20",x"20"),
  1513 => (x"20",x"20",x"20",x"20"),
  1514 => (x"25",x"20",x"20",x"20"),
  1515 => (x"20",x"00",x"0a",x"73"),
  1516 => (x"20",x"20",x"20",x"20"),
  1517 => (x"73",x"20",x"20",x"20"),
  1518 => (x"6c",x"75",x"6f",x"68"),
  1519 => (x"65",x"62",x"20",x"64"),
  1520 => (x"20",x"20",x"20",x"3a"),
  1521 => (x"59",x"52",x"48",x"44"),
  1522 => (x"4e",x"4f",x"54",x"53"),
  1523 => (x"52",x"50",x"20",x"45"),
  1524 => (x"41",x"52",x"47",x"4f"),
  1525 => (x"32",x"20",x"2c",x"4d"),
  1526 => (x"20",x"44",x"4e",x"27"),
  1527 => (x"49",x"52",x"54",x"53"),
  1528 => (x"00",x"0a",x"47",x"4e"),
  1529 => (x"73",x"55",x"00",x"0a"),
  1530 => (x"74",x"20",x"72",x"65"),
  1531 => (x"3a",x"65",x"6d",x"69"),
  1532 => (x"0a",x"64",x"25",x"20"),
  1533 => (x"00",x"00",x"00",x"00"),
  1534 => (x"00",x"00",x"00",x"00"),
  1535 => (x"00",x"00",x"61",x"a8"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
