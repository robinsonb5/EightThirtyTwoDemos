
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"c9",x"01"),
     1 => (x"cf",x"03",x"87",x"cc"),
     2 => (x"87",x"fd",x"00",x"87"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"36",x"27",x"4f",x"00"),
     5 => (x"4f",x"00",x"00",x"00"),
     6 => (x"0e",x"1e",x"18",x"0e"),
     7 => (x"00",x"00",x"44",x"27"),
     8 => (x"48",x"26",x"0f",x"00"),
     9 => (x"08",x"26",x"80",x"ff"),
    10 => (x"c0",x"c0",x"c2",x"4f"),
    11 => (x"13",x"8f",x"27",x"4e"),
    12 => (x"00",x"0f",x"00",x"00"),
    13 => (x"f0",x"c1",x"87",x"fd"),
    14 => (x"43",x"27",x"4e",x"c0"),
    15 => (x"0f",x"00",x"00",x"00"),
    16 => (x"4f",x"87",x"fd",x"00"),
    17 => (x"0e",x"1e",x"18",x"0e"),
    18 => (x"80",x"ff",x"48",x"26"),
    19 => (x"00",x"4f",x"08",x"26"),
    20 => (x"1e",x"1e",x"72",x"1e"),
    21 => (x"6a",x"4a",x"c0",x"ff"),
    22 => (x"98",x"c0",x"c4",x"48"),
    23 => (x"6e",x"58",x"a6",x"c4"),
    24 => (x"87",x"f3",x"ff",x"02"),
    25 => (x"cc",x"7a",x"66",x"cc"),
    26 => (x"26",x"26",x"48",x"66"),
    27 => (x"0e",x"4f",x"26",x"4a"),
    28 => (x"5c",x"5b",x"5a",x"5e"),
    29 => (x"66",x"d4",x"0e",x"5d"),
    30 => (x"15",x"4c",x"c0",x"4d"),
    31 => (x"02",x"9b",x"73",x"4b"),
    32 => (x"73",x"87",x"d6",x"c0"),
    33 => (x"27",x"1e",x"72",x"4a"),
    34 => (x"00",x"00",x"00",x"50"),
    35 => (x"c1",x"86",x"c4",x"0f"),
    36 => (x"73",x"4b",x"15",x"84"),
    37 => (x"ea",x"ff",x"05",x"9b"),
    38 => (x"26",x"48",x"74",x"87"),
    39 => (x"26",x"4c",x"26",x"4d"),
    40 => (x"26",x"4a",x"26",x"4b"),
    41 => (x"5a",x"5e",x"0e",x"4f"),
    42 => (x"0e",x"5d",x"5c",x"5b"),
    43 => (x"4d",x"66",x"d8",x"1e"),
    44 => (x"00",x"15",x"f8",x"27"),
    45 => (x"49",x"76",x"4b",x"00"),
    46 => (x"00",x"15",x"6a",x"27"),
    47 => (x"4c",x"c0",x"79",x"00"),
    48 => (x"03",x"ad",x"b7",x"c0"),
    49 => (x"c0",x"87",x"cd",x"c0"),
    50 => (x"50",x"27",x"1e",x"ed"),
    51 => (x"0f",x"00",x"00",x"00"),
    52 => (x"8d",x"0d",x"86",x"c4"),
    53 => (x"c0",x"05",x"9d",x"75"),
    54 => (x"f0",x"c0",x"87",x"c6"),
    55 => (x"87",x"f6",x"c0",x"53"),
    56 => (x"c0",x"02",x"9d",x"75"),
    57 => (x"49",x"75",x"87",x"f0"),
    58 => (x"e4",x"c0",x"1e",x"72"),
    59 => (x"20",x"27",x"4a",x"66"),
    60 => (x"0f",x"00",x"00",x"15"),
    61 => (x"4a",x"71",x"4a",x"26"),
    62 => (x"82",x"6e",x"4a",x"72"),
    63 => (x"49",x"75",x"53",x"12"),
    64 => (x"e4",x"c0",x"1e",x"72"),
    65 => (x"20",x"27",x"4a",x"66"),
    66 => (x"0f",x"00",x"00",x"15"),
    67 => (x"4d",x"70",x"4a",x"26"),
    68 => (x"ff",x"05",x"9d",x"75"),
    69 => (x"f8",x"27",x"87",x"d0"),
    70 => (x"b7",x"00",x"00",x"15"),
    71 => (x"de",x"c0",x"02",x"ab"),
    72 => (x"dc",x"8b",x"c1",x"87"),
    73 => (x"6b",x"97",x"49",x"66"),
    74 => (x"48",x"66",x"dc",x"51"),
    75 => (x"e0",x"c0",x"80",x"c1"),
    76 => (x"84",x"c1",x"58",x"a6"),
    77 => (x"00",x"15",x"f8",x"27"),
    78 => (x"05",x"ab",x"b7",x"00"),
    79 => (x"dc",x"87",x"e2",x"ff"),
    80 => (x"51",x"c0",x"49",x"66"),
    81 => (x"26",x"26",x"48",x"74"),
    82 => (x"26",x"4c",x"26",x"4d"),
    83 => (x"26",x"4a",x"26",x"4b"),
    84 => (x"5a",x"5e",x"0e",x"4f"),
    85 => (x"0e",x"5d",x"5c",x"5b"),
    86 => (x"76",x"4c",x"c0",x"1e"),
    87 => (x"dc",x"79",x"c0",x"49"),
    88 => (x"66",x"d8",x"4b",x"a6"),
    89 => (x"48",x"66",x"d8",x"4a"),
    90 => (x"a6",x"dc",x"80",x"c1"),
    91 => (x"d8",x"4d",x"12",x"58"),
    92 => (x"75",x"2d",x"b7",x"35"),
    93 => (x"cb",x"c4",x"02",x"9d"),
    94 => (x"c3",x"02",x"6e",x"87"),
    95 => (x"49",x"76",x"87",x"d7"),
    96 => (x"4a",x"75",x"79",x"c0"),
    97 => (x"02",x"ad",x"e3",x"c1"),
    98 => (x"c1",x"87",x"dd",x"c2"),
    99 => (x"c0",x"02",x"aa",x"e4"),
   100 => (x"ec",x"c1",x"87",x"d8"),
   101 => (x"c8",x"c2",x"02",x"aa"),
   102 => (x"aa",x"f3",x"c1",x"87"),
   103 => (x"87",x"e8",x"c1",x"02"),
   104 => (x"02",x"aa",x"f8",x"c1"),
   105 => (x"c2",x"87",x"f2",x"c0"),
   106 => (x"1e",x"ca",x"87",x"d3"),
   107 => (x"00",x"16",x"48",x"27"),
   108 => (x"83",x"c4",x"1e",x"00"),
   109 => (x"8a",x"c4",x"4a",x"73"),
   110 => (x"a5",x"27",x"1e",x"6a"),
   111 => (x"0f",x"00",x"00",x"00"),
   112 => (x"4a",x"70",x"86",x"cc"),
   113 => (x"84",x"72",x"4c",x"74"),
   114 => (x"00",x"16",x"48",x"27"),
   115 => (x"6f",x"27",x"1e",x"00"),
   116 => (x"0f",x"00",x"00",x"00"),
   117 => (x"d4",x"c2",x"86",x"c4"),
   118 => (x"27",x"1e",x"d0",x"87"),
   119 => (x"00",x"00",x"16",x"48"),
   120 => (x"73",x"83",x"c4",x"1e"),
   121 => (x"6a",x"8a",x"c4",x"4a"),
   122 => (x"00",x"a5",x"27",x"1e"),
   123 => (x"cc",x"0f",x"00",x"00"),
   124 => (x"74",x"4a",x"70",x"86"),
   125 => (x"27",x"84",x"72",x"4c"),
   126 => (x"00",x"00",x"16",x"48"),
   127 => (x"00",x"6f",x"27",x"1e"),
   128 => (x"c4",x"0f",x"00",x"00"),
   129 => (x"87",x"e5",x"c1",x"86"),
   130 => (x"4a",x"73",x"83",x"c4"),
   131 => (x"1e",x"6a",x"8a",x"c4"),
   132 => (x"00",x"00",x"6f",x"27"),
   133 => (x"86",x"c4",x"0f",x"00"),
   134 => (x"4c",x"74",x"4a",x"70"),
   135 => (x"cc",x"c1",x"84",x"72"),
   136 => (x"c1",x"49",x"76",x"87"),
   137 => (x"87",x"c5",x"c1",x"79"),
   138 => (x"4a",x"73",x"83",x"c4"),
   139 => (x"1e",x"6a",x"8a",x"c4"),
   140 => (x"00",x"00",x"50",x"27"),
   141 => (x"86",x"c4",x"0f",x"00"),
   142 => (x"f0",x"c0",x"84",x"c1"),
   143 => (x"1e",x"e5",x"c0",x"87"),
   144 => (x"00",x"00",x"50",x"27"),
   145 => (x"86",x"c4",x"0f",x"00"),
   146 => (x"50",x"27",x"1e",x"75"),
   147 => (x"0f",x"00",x"00",x"00"),
   148 => (x"d8",x"c0",x"86",x"c4"),
   149 => (x"ad",x"e5",x"c0",x"87"),
   150 => (x"87",x"c7",x"c0",x"05"),
   151 => (x"79",x"c1",x"49",x"76"),
   152 => (x"75",x"87",x"ca",x"c0"),
   153 => (x"00",x"50",x"27",x"1e"),
   154 => (x"c4",x"0f",x"00",x"00"),
   155 => (x"4a",x"66",x"d8",x"86"),
   156 => (x"c1",x"48",x"66",x"d8"),
   157 => (x"58",x"a6",x"dc",x"80"),
   158 => (x"35",x"d8",x"4d",x"12"),
   159 => (x"9d",x"75",x"2d",x"b7"),
   160 => (x"87",x"f5",x"fb",x"05"),
   161 => (x"26",x"26",x"48",x"74"),
   162 => (x"26",x"4c",x"26",x"4d"),
   163 => (x"26",x"4a",x"26",x"4b"),
   164 => (x"00",x"1f",x"0f",x"4f"),
   165 => (x"c0",x"1e",x"72",x"1e"),
   166 => (x"49",x"66",x"cc",x"4a"),
   167 => (x"06",x"a9",x"b7",x"c0"),
   168 => (x"c8",x"87",x"d2",x"c0"),
   169 => (x"80",x"c4",x"48",x"66"),
   170 => (x"c1",x"58",x"a6",x"cc"),
   171 => (x"b7",x"66",x"cc",x"82"),
   172 => (x"ee",x"ff",x"04",x"aa"),
   173 => (x"26",x"4a",x"26",x"87"),
   174 => (x"5a",x"5e",x"0e",x"4f"),
   175 => (x"0e",x"5d",x"5c",x"5b"),
   176 => (x"c1",x"4c",x"66",x"d4"),
   177 => (x"73",x"4b",x"c0",x"4d"),
   178 => (x"72",x"92",x"c4",x"4a"),
   179 => (x"15",x"10",x"27",x"4a"),
   180 => (x"6a",x"82",x"00",x"00"),
   181 => (x"6a",x"49",x"6c",x"7c"),
   182 => (x"c0",x"02",x"a9",x"b7"),
   183 => (x"1e",x"6c",x"87",x"e0"),
   184 => (x"92",x"c4",x"4a",x"73"),
   185 => (x"10",x"27",x"4a",x"72"),
   186 => (x"82",x"00",x"00",x"15"),
   187 => (x"7b",x"27",x"1e",x"6a"),
   188 => (x"1e",x"00",x"00",x"15"),
   189 => (x"00",x"01",x"51",x"27"),
   190 => (x"86",x"cc",x"0f",x"00"),
   191 => (x"66",x"d8",x"4d",x"c0"),
   192 => (x"27",x"1e",x"74",x"1e"),
   193 => (x"00",x"00",x"02",x"94"),
   194 => (x"73",x"86",x"c8",x"0f"),
   195 => (x"72",x"92",x"c4",x"4a"),
   196 => (x"15",x"10",x"27",x"4a"),
   197 => (x"6c",x"82",x"00",x"00"),
   198 => (x"a9",x"b7",x"6a",x"49"),
   199 => (x"87",x"e0",x"c0",x"02"),
   200 => (x"4a",x"73",x"1e",x"6c"),
   201 => (x"4a",x"72",x"92",x"c4"),
   202 => (x"00",x"15",x"10",x"27"),
   203 => (x"1e",x"6a",x"82",x"00"),
   204 => (x"00",x"15",x"ba",x"27"),
   205 => (x"51",x"27",x"1e",x"00"),
   206 => (x"0f",x"00",x"00",x"01"),
   207 => (x"4d",x"c0",x"86",x"cc"),
   208 => (x"b7",x"c4",x"83",x"c1"),
   209 => (x"fe",x"fd",x"04",x"ab"),
   210 => (x"26",x"48",x"75",x"87"),
   211 => (x"26",x"4c",x"26",x"4d"),
   212 => (x"26",x"4a",x"26",x"4b"),
   213 => (x"5a",x"5e",x"0e",x"4f"),
   214 => (x"0e",x"5d",x"5c",x"5b"),
   215 => (x"66",x"dc",x"8e",x"c8"),
   216 => (x"73",x"4d",x"c1",x"4b"),
   217 => (x"49",x"a6",x"c4",x"4c"),
   218 => (x"49",x"76",x"79",x"73"),
   219 => (x"4a",x"73",x"79",x"6b"),
   220 => (x"d5",x"c1",x"82",x"cc"),
   221 => (x"d5",x"d5",x"d5",x"d5"),
   222 => (x"ea",x"ea",x"c2",x"7b"),
   223 => (x"7a",x"ea",x"ea",x"ea"),
   224 => (x"7b",x"97",x"cc",x"ff"),
   225 => (x"82",x"cf",x"4a",x"73"),
   226 => (x"6b",x"52",x"f3",x"c0"),
   227 => (x"d5",x"d5",x"c1",x"49"),
   228 => (x"b7",x"cc",x"d7",x"d5"),
   229 => (x"d2",x"c0",x"02",x"a9"),
   230 => (x"27",x"1e",x"6b",x"87"),
   231 => (x"00",x"00",x"06",x"47"),
   232 => (x"01",x"51",x"27",x"1e"),
   233 => (x"c8",x"0f",x"00",x"00"),
   234 => (x"73",x"4d",x"c0",x"86"),
   235 => (x"6a",x"82",x"cc",x"4a"),
   236 => (x"ea",x"f3",x"c0",x"49"),
   237 => (x"b7",x"ea",x"ea",x"ea"),
   238 => (x"d6",x"c0",x"02",x"a9"),
   239 => (x"cc",x"4a",x"73",x"87"),
   240 => (x"27",x"1e",x"6a",x"82"),
   241 => (x"00",x"00",x"06",x"81"),
   242 => (x"01",x"51",x"27",x"1e"),
   243 => (x"c8",x"0f",x"00",x"00"),
   244 => (x"74",x"4d",x"c0",x"86"),
   245 => (x"d2",x"82",x"c1",x"4a"),
   246 => (x"4a",x"66",x"c4",x"52"),
   247 => (x"dc",x"fb",x"82",x"ce"),
   248 => (x"49",x"6b",x"7a",x"9f"),
   249 => (x"d1",x"d5",x"d5",x"c1"),
   250 => (x"a9",x"b7",x"cc",x"cb"),
   251 => (x"87",x"d2",x"c0",x"02"),
   252 => (x"bb",x"27",x"1e",x"6b"),
   253 => (x"1e",x"00",x"00",x"06"),
   254 => (x"00",x"01",x"51",x"27"),
   255 => (x"86",x"c8",x"0f",x"00"),
   256 => (x"4a",x"73",x"4d",x"c0"),
   257 => (x"49",x"6a",x"82",x"cc"),
   258 => (x"ea",x"ca",x"f7",x"fe"),
   259 => (x"c0",x"02",x"a9",x"ea"),
   260 => (x"4a",x"73",x"87",x"d6"),
   261 => (x"1e",x"6a",x"82",x"cc"),
   262 => (x"00",x"06",x"f7",x"27"),
   263 => (x"51",x"27",x"1e",x"00"),
   264 => (x"0f",x"00",x"00",x"01"),
   265 => (x"4d",x"c0",x"86",x"c8"),
   266 => (x"1e",x"66",x"e0",x"c0"),
   267 => (x"94",x"27",x"1e",x"73"),
   268 => (x"0f",x"00",x"00",x"02"),
   269 => (x"49",x"6b",x"86",x"c8"),
   270 => (x"d1",x"d5",x"d5",x"c1"),
   271 => (x"a9",x"b7",x"cc",x"cb"),
   272 => (x"87",x"d2",x"c0",x"02"),
   273 => (x"33",x"27",x"1e",x"6b"),
   274 => (x"1e",x"00",x"00",x"07"),
   275 => (x"00",x"01",x"51",x"27"),
   276 => (x"86",x"c8",x"0f",x"00"),
   277 => (x"4a",x"73",x"4d",x"c0"),
   278 => (x"49",x"6a",x"82",x"cc"),
   279 => (x"ea",x"ca",x"f7",x"fe"),
   280 => (x"c0",x"02",x"a9",x"ea"),
   281 => (x"4a",x"73",x"87",x"d6"),
   282 => (x"1e",x"6a",x"82",x"cc"),
   283 => (x"00",x"07",x"6c",x"27"),
   284 => (x"51",x"27",x"1e",x"00"),
   285 => (x"0f",x"00",x"00",x"01"),
   286 => (x"4d",x"c0",x"86",x"c8"),
   287 => (x"82",x"c2",x"4a",x"74"),
   288 => (x"4a",x"74",x"52",x"cf"),
   289 => (x"52",x"f0",x"82",x"cd"),
   290 => (x"c4",x"48",x"6c",x"97"),
   291 => (x"49",x"6e",x"58",x"a6"),
   292 => (x"a9",x"b7",x"cc",x"c3"),
   293 => (x"87",x"d5",x"c0",x"02"),
   294 => (x"72",x"4a",x"6c",x"97"),
   295 => (x"07",x"a5",x"27",x"1e"),
   296 => (x"27",x"1e",x"00",x"00"),
   297 => (x"00",x"00",x"01",x"51"),
   298 => (x"c0",x"86",x"c8",x"0f"),
   299 => (x"c1",x"4a",x"74",x"4d"),
   300 => (x"c4",x"48",x"12",x"82"),
   301 => (x"49",x"6e",x"58",x"a6"),
   302 => (x"02",x"a9",x"b7",x"d2"),
   303 => (x"74",x"87",x"d9",x"c0"),
   304 => (x"97",x"82",x"c1",x"4a"),
   305 => (x"1e",x"72",x"4a",x"6a"),
   306 => (x"00",x"07",x"cd",x"27"),
   307 => (x"51",x"27",x"1e",x"00"),
   308 => (x"0f",x"00",x"00",x"01"),
   309 => (x"4d",x"c0",x"86",x"c8"),
   310 => (x"82",x"c2",x"4a",x"74"),
   311 => (x"a6",x"c4",x"48",x"12"),
   312 => (x"cf",x"49",x"6e",x"58"),
   313 => (x"c0",x"02",x"a9",x"b7"),
   314 => (x"4a",x"74",x"87",x"d9"),
   315 => (x"6a",x"97",x"82",x"c2"),
   316 => (x"27",x"1e",x"72",x"4a"),
   317 => (x"00",x"00",x"07",x"f5"),
   318 => (x"01",x"51",x"27",x"1e"),
   319 => (x"c8",x"0f",x"00",x"00"),
   320 => (x"74",x"4d",x"c0",x"86"),
   321 => (x"12",x"82",x"c3",x"4a"),
   322 => (x"58",x"a6",x"c4",x"48"),
   323 => (x"d5",x"c1",x"49",x"6e"),
   324 => (x"c0",x"02",x"a9",x"b7"),
   325 => (x"4a",x"74",x"87",x"d9"),
   326 => (x"6a",x"97",x"82",x"c3"),
   327 => (x"27",x"1e",x"72",x"4a"),
   328 => (x"00",x"00",x"08",x"1d"),
   329 => (x"01",x"51",x"27",x"1e"),
   330 => (x"c8",x"0f",x"00",x"00"),
   331 => (x"74",x"4d",x"c0",x"86"),
   332 => (x"12",x"82",x"cc",x"4a"),
   333 => (x"58",x"a6",x"c4",x"48"),
   334 => (x"ea",x"c2",x"49",x"6e"),
   335 => (x"c0",x"02",x"a9",x"b7"),
   336 => (x"4a",x"74",x"87",x"d9"),
   337 => (x"6a",x"97",x"82",x"cc"),
   338 => (x"27",x"1e",x"72",x"4a"),
   339 => (x"00",x"00",x"08",x"45"),
   340 => (x"01",x"51",x"27",x"1e"),
   341 => (x"c8",x"0f",x"00",x"00"),
   342 => (x"74",x"4d",x"c0",x"86"),
   343 => (x"12",x"82",x"cd",x"4a"),
   344 => (x"58",x"a6",x"c4",x"48"),
   345 => (x"f0",x"c3",x"49",x"6e"),
   346 => (x"c0",x"02",x"a9",x"b7"),
   347 => (x"4a",x"74",x"87",x"d9"),
   348 => (x"6a",x"97",x"82",x"cd"),
   349 => (x"27",x"1e",x"72",x"4a"),
   350 => (x"00",x"00",x"08",x"6e"),
   351 => (x"01",x"51",x"27",x"1e"),
   352 => (x"c8",x"0f",x"00",x"00"),
   353 => (x"74",x"4d",x"c0",x"86"),
   354 => (x"12",x"82",x"ce",x"4a"),
   355 => (x"58",x"a6",x"c4",x"48"),
   356 => (x"dc",x"c3",x"49",x"6e"),
   357 => (x"c0",x"02",x"a9",x"b7"),
   358 => (x"4a",x"74",x"87",x"d9"),
   359 => (x"6a",x"97",x"82",x"ce"),
   360 => (x"27",x"1e",x"72",x"4a"),
   361 => (x"00",x"00",x"08",x"97"),
   362 => (x"01",x"51",x"27",x"1e"),
   363 => (x"c8",x"0f",x"00",x"00"),
   364 => (x"74",x"4d",x"c0",x"86"),
   365 => (x"12",x"82",x"cf",x"4a"),
   366 => (x"58",x"a6",x"c4",x"48"),
   367 => (x"fe",x"c3",x"49",x"6e"),
   368 => (x"c0",x"02",x"a9",x"b7"),
   369 => (x"4a",x"74",x"87",x"d9"),
   370 => (x"6a",x"97",x"82",x"cf"),
   371 => (x"27",x"1e",x"72",x"4a"),
   372 => (x"00",x"00",x"08",x"c0"),
   373 => (x"01",x"51",x"27",x"1e"),
   374 => (x"c8",x"0f",x"00",x"00"),
   375 => (x"c4",x"4d",x"c0",x"86"),
   376 => (x"48",x"bf",x"9f",x"66"),
   377 => (x"6e",x"58",x"a6",x"c4"),
   378 => (x"cc",x"cb",x"c1",x"49"),
   379 => (x"c0",x"02",x"a9",x"b7"),
   380 => (x"66",x"c4",x"87",x"d7"),
   381 => (x"72",x"4a",x"bf",x"9f"),
   382 => (x"08",x"e9",x"27",x"1e"),
   383 => (x"27",x"1e",x"00",x"00"),
   384 => (x"00",x"00",x"01",x"51"),
   385 => (x"c0",x"86",x"c8",x"0f"),
   386 => (x"4a",x"66",x"c4",x"4d"),
   387 => (x"6a",x"9f",x"82",x"ce"),
   388 => (x"58",x"a6",x"c4",x"48"),
   389 => (x"fb",x"cf",x"49",x"6e"),
   390 => (x"02",x"a9",x"b7",x"dc"),
   391 => (x"c4",x"87",x"da",x"c0"),
   392 => (x"82",x"ce",x"4a",x"66"),
   393 => (x"72",x"4a",x"6a",x"9f"),
   394 => (x"09",x"11",x"27",x"1e"),
   395 => (x"27",x"1e",x"00",x"00"),
   396 => (x"00",x"00",x"01",x"51"),
   397 => (x"c0",x"86",x"c8",x"0f"),
   398 => (x"c8",x"48",x"75",x"4d"),
   399 => (x"26",x"4d",x"26",x"86"),
   400 => (x"26",x"4b",x"26",x"4c"),
   401 => (x"42",x"4f",x"26",x"4a"),
   402 => (x"20",x"65",x"74",x"79"),
   403 => (x"63",x"65",x"68",x"63"),
   404 => (x"61",x"66",x"20",x"6b"),
   405 => (x"64",x"65",x"6c",x"69"),
   406 => (x"65",x"62",x"28",x"20"),
   407 => (x"65",x"72",x"6f",x"66"),
   408 => (x"63",x"61",x"63",x"20"),
   409 => (x"72",x"20",x"65",x"68"),
   410 => (x"65",x"72",x"66",x"65"),
   411 => (x"20",x"29",x"68",x"73"),
   412 => (x"30",x"20",x"74",x"61"),
   413 => (x"6f",x"67",x"28",x"20"),
   414 => (x"78",x"30",x"20",x"74"),
   415 => (x"0a",x"29",x"64",x"25"),
   416 => (x"74",x"79",x"42",x"00"),
   417 => (x"68",x"63",x"20",x"65"),
   418 => (x"20",x"6b",x"63",x"65"),
   419 => (x"6c",x"69",x"61",x"66"),
   420 => (x"28",x"20",x"64",x"65"),
   421 => (x"6f",x"66",x"65",x"62"),
   422 => (x"63",x"20",x"65",x"72"),
   423 => (x"65",x"68",x"63",x"61"),
   424 => (x"66",x"65",x"72",x"20"),
   425 => (x"68",x"73",x"65",x"72"),
   426 => (x"74",x"61",x"20",x"29"),
   427 => (x"28",x"20",x"33",x"20"),
   428 => (x"20",x"74",x"6f",x"67"),
   429 => (x"64",x"25",x"78",x"30"),
   430 => (x"42",x"00",x"0a",x"29"),
   431 => (x"20",x"65",x"74",x"79"),
   432 => (x"63",x"65",x"68",x"63"),
   433 => (x"20",x"32",x"20",x"6b"),
   434 => (x"6c",x"69",x"61",x"66"),
   435 => (x"28",x"20",x"64",x"65"),
   436 => (x"6f",x"66",x"65",x"62"),
   437 => (x"63",x"20",x"65",x"72"),
   438 => (x"65",x"68",x"63",x"61"),
   439 => (x"66",x"65",x"72",x"20"),
   440 => (x"68",x"73",x"65",x"72"),
   441 => (x"74",x"61",x"20",x"29"),
   442 => (x"28",x"20",x"30",x"20"),
   443 => (x"20",x"74",x"6f",x"67"),
   444 => (x"64",x"25",x"78",x"30"),
   445 => (x"42",x"00",x"0a",x"29"),
   446 => (x"20",x"65",x"74",x"79"),
   447 => (x"63",x"65",x"68",x"63"),
   448 => (x"20",x"32",x"20",x"6b"),
   449 => (x"6c",x"69",x"61",x"66"),
   450 => (x"28",x"20",x"64",x"65"),
   451 => (x"6f",x"66",x"65",x"62"),
   452 => (x"63",x"20",x"65",x"72"),
   453 => (x"65",x"68",x"63",x"61"),
   454 => (x"66",x"65",x"72",x"20"),
   455 => (x"68",x"73",x"65",x"72"),
   456 => (x"74",x"61",x"20",x"29"),
   457 => (x"28",x"20",x"33",x"20"),
   458 => (x"20",x"74",x"6f",x"67"),
   459 => (x"64",x"25",x"78",x"30"),
   460 => (x"42",x"00",x"0a",x"29"),
   461 => (x"20",x"65",x"74",x"79"),
   462 => (x"63",x"65",x"68",x"63"),
   463 => (x"61",x"66",x"20",x"6b"),
   464 => (x"64",x"65",x"6c",x"69"),
   465 => (x"66",x"61",x"28",x"20"),
   466 => (x"20",x"72",x"65",x"74"),
   467 => (x"68",x"63",x"61",x"63"),
   468 => (x"65",x"72",x"20",x"65"),
   469 => (x"73",x"65",x"72",x"66"),
   470 => (x"61",x"20",x"29",x"68"),
   471 => (x"20",x"30",x"20",x"74"),
   472 => (x"74",x"6f",x"67",x"28"),
   473 => (x"25",x"78",x"30",x"20"),
   474 => (x"00",x"0a",x"29",x"64"),
   475 => (x"65",x"74",x"79",x"42"),
   476 => (x"65",x"68",x"63",x"20"),
   477 => (x"66",x"20",x"6b",x"63"),
   478 => (x"65",x"6c",x"69",x"61"),
   479 => (x"61",x"28",x"20",x"64"),
   480 => (x"72",x"65",x"74",x"66"),
   481 => (x"63",x"61",x"63",x"20"),
   482 => (x"72",x"20",x"65",x"68"),
   483 => (x"65",x"72",x"66",x"65"),
   484 => (x"20",x"29",x"68",x"73"),
   485 => (x"33",x"20",x"74",x"61"),
   486 => (x"6f",x"67",x"28",x"20"),
   487 => (x"78",x"30",x"20",x"74"),
   488 => (x"0a",x"29",x"64",x"25"),
   489 => (x"74",x"79",x"42",x"00"),
   490 => (x"65",x"72",x"20",x"65"),
   491 => (x"63",x"20",x"64",x"61"),
   492 => (x"6b",x"63",x"65",x"68"),
   493 => (x"69",x"61",x"66",x"20"),
   494 => (x"20",x"64",x"65",x"6c"),
   495 => (x"30",x"20",x"74",x"61"),
   496 => (x"6f",x"67",x"28",x"20"),
   497 => (x"78",x"30",x"20",x"74"),
   498 => (x"0a",x"29",x"64",x"25"),
   499 => (x"74",x"79",x"42",x"00"),
   500 => (x"65",x"72",x"20",x"65"),
   501 => (x"63",x"20",x"64",x"61"),
   502 => (x"6b",x"63",x"65",x"68"),
   503 => (x"69",x"61",x"66",x"20"),
   504 => (x"20",x"64",x"65",x"6c"),
   505 => (x"31",x"20",x"74",x"61"),
   506 => (x"6f",x"67",x"28",x"20"),
   507 => (x"78",x"30",x"20",x"74"),
   508 => (x"0a",x"29",x"64",x"25"),
   509 => (x"74",x"79",x"42",x"00"),
   510 => (x"65",x"72",x"20",x"65"),
   511 => (x"63",x"20",x"64",x"61"),
   512 => (x"6b",x"63",x"65",x"68"),
   513 => (x"69",x"61",x"66",x"20"),
   514 => (x"20",x"64",x"65",x"6c"),
   515 => (x"32",x"20",x"74",x"61"),
   516 => (x"6f",x"67",x"28",x"20"),
   517 => (x"78",x"30",x"20",x"74"),
   518 => (x"0a",x"29",x"64",x"25"),
   519 => (x"74",x"79",x"42",x"00"),
   520 => (x"65",x"72",x"20",x"65"),
   521 => (x"63",x"20",x"64",x"61"),
   522 => (x"6b",x"63",x"65",x"68"),
   523 => (x"69",x"61",x"66",x"20"),
   524 => (x"20",x"64",x"65",x"6c"),
   525 => (x"33",x"20",x"74",x"61"),
   526 => (x"6f",x"67",x"28",x"20"),
   527 => (x"78",x"30",x"20",x"74"),
   528 => (x"0a",x"29",x"64",x"25"),
   529 => (x"74",x"79",x"42",x"00"),
   530 => (x"65",x"72",x"20",x"65"),
   531 => (x"63",x"20",x"64",x"61"),
   532 => (x"6b",x"63",x"65",x"68"),
   533 => (x"69",x"61",x"66",x"20"),
   534 => (x"20",x"64",x"65",x"6c"),
   535 => (x"31",x"20",x"74",x"61"),
   536 => (x"67",x"28",x"20",x"32"),
   537 => (x"30",x"20",x"74",x"6f"),
   538 => (x"29",x"64",x"25",x"78"),
   539 => (x"79",x"42",x"00",x"0a"),
   540 => (x"72",x"20",x"65",x"74"),
   541 => (x"20",x"64",x"61",x"65"),
   542 => (x"63",x"65",x"68",x"63"),
   543 => (x"61",x"66",x"20",x"6b"),
   544 => (x"64",x"65",x"6c",x"69"),
   545 => (x"20",x"74",x"61",x"20"),
   546 => (x"28",x"20",x"33",x"31"),
   547 => (x"20",x"74",x"6f",x"67"),
   548 => (x"64",x"25",x"78",x"30"),
   549 => (x"42",x"00",x"0a",x"29"),
   550 => (x"20",x"65",x"74",x"79"),
   551 => (x"64",x"61",x"65",x"72"),
   552 => (x"65",x"68",x"63",x"20"),
   553 => (x"66",x"20",x"6b",x"63"),
   554 => (x"65",x"6c",x"69",x"61"),
   555 => (x"74",x"61",x"20",x"64"),
   556 => (x"20",x"34",x"31",x"20"),
   557 => (x"74",x"6f",x"67",x"28"),
   558 => (x"25",x"78",x"30",x"20"),
   559 => (x"00",x"0a",x"29",x"64"),
   560 => (x"65",x"74",x"79",x"42"),
   561 => (x"61",x"65",x"72",x"20"),
   562 => (x"68",x"63",x"20",x"64"),
   563 => (x"20",x"6b",x"63",x"65"),
   564 => (x"6c",x"69",x"61",x"66"),
   565 => (x"61",x"20",x"64",x"65"),
   566 => (x"35",x"31",x"20",x"74"),
   567 => (x"6f",x"67",x"28",x"20"),
   568 => (x"78",x"30",x"20",x"74"),
   569 => (x"0a",x"29",x"64",x"25"),
   570 => (x"72",x"6f",x"57",x"00"),
   571 => (x"65",x"72",x"20",x"64"),
   572 => (x"63",x"20",x"64",x"61"),
   573 => (x"6b",x"63",x"65",x"68"),
   574 => (x"69",x"61",x"66",x"20"),
   575 => (x"20",x"64",x"65",x"6c"),
   576 => (x"30",x"20",x"74",x"61"),
   577 => (x"6f",x"67",x"28",x"20"),
   578 => (x"78",x"30",x"20",x"74"),
   579 => (x"0a",x"29",x"64",x"25"),
   580 => (x"72",x"6f",x"57",x"00"),
   581 => (x"65",x"72",x"20",x"64"),
   582 => (x"63",x"20",x"64",x"61"),
   583 => (x"6b",x"63",x"65",x"68"),
   584 => (x"69",x"61",x"66",x"20"),
   585 => (x"20",x"64",x"65",x"6c"),
   586 => (x"37",x"20",x"74",x"61"),
   587 => (x"6f",x"67",x"28",x"20"),
   588 => (x"78",x"30",x"20",x"74"),
   589 => (x"0a",x"29",x"64",x"25"),
   590 => (x"5a",x"5e",x"0e",x"00"),
   591 => (x"0e",x"5d",x"5c",x"5b"),
   592 => (x"fc",x"ee",x"ea",x"c2"),
   593 => (x"d4",x"4d",x"dd",x"f3"),
   594 => (x"66",x"d4",x"4c",x"66"),
   595 => (x"c8",x"d2",x"c4",x"49"),
   596 => (x"66",x"d4",x"79",x"f3"),
   597 => (x"c1",x"82",x"c4",x"4a"),
   598 => (x"d9",x"d6",x"d5",x"c4"),
   599 => (x"66",x"d4",x"7a",x"f7"),
   600 => (x"c2",x"82",x"c8",x"4a"),
   601 => (x"ea",x"da",x"e6",x"c8"),
   602 => (x"66",x"d4",x"7a",x"fb"),
   603 => (x"c3",x"82",x"cc",x"4a"),
   604 => (x"fb",x"de",x"f7",x"cc"),
   605 => (x"66",x"d4",x"7a",x"ff"),
   606 => (x"c1",x"82",x"d0",x"4a"),
   607 => (x"ea",x"da",x"d5",x"d5"),
   608 => (x"66",x"d4",x"7a",x"ea"),
   609 => (x"4a",x"82",x"c2",x"4a"),
   610 => (x"e2",x"c0",x"4b",x"6a"),
   611 => (x"d5",x"d1",x"f4",x"cc"),
   612 => (x"c0",x"02",x"ab",x"b7"),
   613 => (x"1e",x"73",x"87",x"d0"),
   614 => (x"00",x"0a",x"a3",x"27"),
   615 => (x"51",x"27",x"1e",x"00"),
   616 => (x"0f",x"00",x"00",x"01"),
   617 => (x"4a",x"74",x"86",x"c8"),
   618 => (x"6a",x"4a",x"82",x"c6"),
   619 => (x"dd",x"e6",x"c1",x"4b"),
   620 => (x"b7",x"d9",x"e2",x"f8"),
   621 => (x"d0",x"c0",x"02",x"ab"),
   622 => (x"27",x"1e",x"73",x"87"),
   623 => (x"00",x"00",x"0a",x"de"),
   624 => (x"01",x"51",x"27",x"1e"),
   625 => (x"c8",x"0f",x"00",x"00"),
   626 => (x"ca",x"4a",x"74",x"86"),
   627 => (x"4b",x"6a",x"4a",x"82"),
   628 => (x"c0",x"02",x"ab",x"75"),
   629 => (x"1e",x"73",x"87",x"d0"),
   630 => (x"00",x"0b",x"19",x"27"),
   631 => (x"51",x"27",x"1e",x"00"),
   632 => (x"0f",x"00",x"00",x"01"),
   633 => (x"4a",x"74",x"86",x"c8"),
   634 => (x"6a",x"4a",x"82",x"ce"),
   635 => (x"f5",x"ff",x"ee",x"4b"),
   636 => (x"02",x"ab",x"d5",x"d5"),
   637 => (x"73",x"87",x"d0",x"c0"),
   638 => (x"0b",x"55",x"27",x"1e"),
   639 => (x"27",x"1e",x"00",x"00"),
   640 => (x"00",x"00",x"01",x"51"),
   641 => (x"d8",x"86",x"c8",x"0f"),
   642 => (x"66",x"d8",x"1e",x"66"),
   643 => (x"02",x"94",x"27",x"1e"),
   644 => (x"c8",x"0f",x"00",x"00"),
   645 => (x"c2",x"4a",x"74",x"86"),
   646 => (x"4b",x"6a",x"4a",x"82"),
   647 => (x"f4",x"cc",x"e2",x"c0"),
   648 => (x"ab",x"b7",x"d5",x"d1"),
   649 => (x"87",x"d0",x"c0",x"02"),
   650 => (x"91",x"27",x"1e",x"73"),
   651 => (x"1e",x"00",x"00",x"0b"),
   652 => (x"00",x"01",x"51",x"27"),
   653 => (x"86",x"c8",x"0f",x"00"),
   654 => (x"82",x"c6",x"4a",x"74"),
   655 => (x"c1",x"4b",x"6a",x"4a"),
   656 => (x"e2",x"f8",x"dd",x"e6"),
   657 => (x"02",x"ab",x"b7",x"d9"),
   658 => (x"73",x"87",x"d0",x"c0"),
   659 => (x"0b",x"cb",x"27",x"1e"),
   660 => (x"27",x"1e",x"00",x"00"),
   661 => (x"00",x"00",x"01",x"51"),
   662 => (x"74",x"86",x"c8",x"0f"),
   663 => (x"4a",x"82",x"ca",x"4a"),
   664 => (x"ab",x"75",x"4b",x"6a"),
   665 => (x"87",x"d0",x"c0",x"02"),
   666 => (x"05",x"27",x"1e",x"73"),
   667 => (x"1e",x"00",x"00",x"0c"),
   668 => (x"00",x"01",x"51",x"27"),
   669 => (x"86",x"c8",x"0f",x"00"),
   670 => (x"82",x"ce",x"4a",x"74"),
   671 => (x"ee",x"4b",x"6a",x"4a"),
   672 => (x"d5",x"d5",x"f5",x"ff"),
   673 => (x"d0",x"c0",x"02",x"ab"),
   674 => (x"27",x"1e",x"73",x"87"),
   675 => (x"00",x"00",x"0c",x"40"),
   676 => (x"01",x"51",x"27",x"1e"),
   677 => (x"c8",x"0f",x"00",x"00"),
   678 => (x"26",x"4d",x"26",x"86"),
   679 => (x"26",x"4b",x"26",x"4c"),
   680 => (x"41",x"4f",x"26",x"4a"),
   681 => (x"6e",x"67",x"69",x"6c"),
   682 => (x"65",x"68",x"63",x"20"),
   683 => (x"66",x"20",x"6b",x"63"),
   684 => (x"65",x"6c",x"69",x"61"),
   685 => (x"62",x"28",x"20",x"64"),
   686 => (x"72",x"6f",x"66",x"65"),
   687 => (x"61",x"63",x"20",x"65"),
   688 => (x"20",x"65",x"68",x"63"),
   689 => (x"72",x"66",x"65",x"72"),
   690 => (x"29",x"68",x"73",x"65"),
   691 => (x"20",x"74",x"61",x"20"),
   692 => (x"67",x"28",x"20",x"32"),
   693 => (x"30",x"20",x"74",x"6f"),
   694 => (x"29",x"64",x"25",x"78"),
   695 => (x"6c",x"41",x"00",x"0a"),
   696 => (x"20",x"6e",x"67",x"69"),
   697 => (x"63",x"65",x"68",x"63"),
   698 => (x"61",x"66",x"20",x"6b"),
   699 => (x"64",x"65",x"6c",x"69"),
   700 => (x"65",x"62",x"28",x"20"),
   701 => (x"65",x"72",x"6f",x"66"),
   702 => (x"63",x"61",x"63",x"20"),
   703 => (x"72",x"20",x"65",x"68"),
   704 => (x"65",x"72",x"66",x"65"),
   705 => (x"20",x"29",x"68",x"73"),
   706 => (x"36",x"20",x"74",x"61"),
   707 => (x"6f",x"67",x"28",x"20"),
   708 => (x"78",x"30",x"20",x"74"),
   709 => (x"0a",x"29",x"64",x"25"),
   710 => (x"69",x"6c",x"41",x"00"),
   711 => (x"63",x"20",x"6e",x"67"),
   712 => (x"6b",x"63",x"65",x"68"),
   713 => (x"69",x"61",x"66",x"20"),
   714 => (x"20",x"64",x"65",x"6c"),
   715 => (x"66",x"65",x"62",x"28"),
   716 => (x"20",x"65",x"72",x"6f"),
   717 => (x"68",x"63",x"61",x"63"),
   718 => (x"65",x"72",x"20",x"65"),
   719 => (x"73",x"65",x"72",x"66"),
   720 => (x"61",x"20",x"29",x"68"),
   721 => (x"30",x"31",x"20",x"74"),
   722 => (x"6f",x"67",x"28",x"20"),
   723 => (x"78",x"30",x"20",x"74"),
   724 => (x"0a",x"29",x"64",x"25"),
   725 => (x"69",x"6c",x"41",x"00"),
   726 => (x"63",x"20",x"6e",x"67"),
   727 => (x"6b",x"63",x"65",x"68"),
   728 => (x"69",x"61",x"66",x"20"),
   729 => (x"20",x"64",x"65",x"6c"),
   730 => (x"66",x"65",x"62",x"28"),
   731 => (x"20",x"65",x"72",x"6f"),
   732 => (x"68",x"63",x"61",x"63"),
   733 => (x"65",x"72",x"20",x"65"),
   734 => (x"73",x"65",x"72",x"66"),
   735 => (x"61",x"20",x"29",x"68"),
   736 => (x"34",x"31",x"20",x"74"),
   737 => (x"6f",x"67",x"28",x"20"),
   738 => (x"78",x"30",x"20",x"74"),
   739 => (x"0a",x"29",x"64",x"25"),
   740 => (x"69",x"6c",x"41",x"00"),
   741 => (x"63",x"20",x"6e",x"67"),
   742 => (x"6b",x"63",x"65",x"68"),
   743 => (x"69",x"61",x"66",x"20"),
   744 => (x"20",x"64",x"65",x"6c"),
   745 => (x"74",x"66",x"61",x"28"),
   746 => (x"63",x"20",x"72",x"65"),
   747 => (x"65",x"68",x"63",x"61"),
   748 => (x"66",x"65",x"72",x"20"),
   749 => (x"68",x"73",x"65",x"72"),
   750 => (x"74",x"61",x"20",x"29"),
   751 => (x"28",x"20",x"32",x"20"),
   752 => (x"20",x"74",x"6f",x"67"),
   753 => (x"64",x"25",x"78",x"30"),
   754 => (x"41",x"00",x"0a",x"29"),
   755 => (x"6e",x"67",x"69",x"6c"),
   756 => (x"65",x"68",x"63",x"20"),
   757 => (x"66",x"20",x"6b",x"63"),
   758 => (x"65",x"6c",x"69",x"61"),
   759 => (x"61",x"28",x"20",x"64"),
   760 => (x"72",x"65",x"74",x"66"),
   761 => (x"63",x"61",x"63",x"20"),
   762 => (x"72",x"20",x"65",x"68"),
   763 => (x"65",x"72",x"66",x"65"),
   764 => (x"20",x"29",x"68",x"73"),
   765 => (x"36",x"20",x"74",x"61"),
   766 => (x"6f",x"67",x"28",x"20"),
   767 => (x"78",x"30",x"20",x"74"),
   768 => (x"0a",x"29",x"64",x"25"),
   769 => (x"69",x"6c",x"41",x"00"),
   770 => (x"63",x"20",x"6e",x"67"),
   771 => (x"6b",x"63",x"65",x"68"),
   772 => (x"69",x"61",x"66",x"20"),
   773 => (x"20",x"64",x"65",x"6c"),
   774 => (x"74",x"66",x"61",x"28"),
   775 => (x"63",x"20",x"72",x"65"),
   776 => (x"65",x"68",x"63",x"61"),
   777 => (x"66",x"65",x"72",x"20"),
   778 => (x"68",x"73",x"65",x"72"),
   779 => (x"74",x"61",x"20",x"29"),
   780 => (x"20",x"30",x"31",x"20"),
   781 => (x"74",x"6f",x"67",x"28"),
   782 => (x"25",x"78",x"30",x"20"),
   783 => (x"00",x"0a",x"29",x"64"),
   784 => (x"67",x"69",x"6c",x"41"),
   785 => (x"68",x"63",x"20",x"6e"),
   786 => (x"20",x"6b",x"63",x"65"),
   787 => (x"6c",x"69",x"61",x"66"),
   788 => (x"28",x"20",x"64",x"65"),
   789 => (x"65",x"74",x"66",x"61"),
   790 => (x"61",x"63",x"20",x"72"),
   791 => (x"20",x"65",x"68",x"63"),
   792 => (x"72",x"66",x"65",x"72"),
   793 => (x"29",x"68",x"73",x"65"),
   794 => (x"20",x"74",x"61",x"20"),
   795 => (x"28",x"20",x"34",x"31"),
   796 => (x"20",x"74",x"6f",x"67"),
   797 => (x"64",x"25",x"78",x"30"),
   798 => (x"0e",x"00",x"0a",x"29"),
   799 => (x"5c",x"5b",x"5a",x"5e"),
   800 => (x"e0",x"c0",x"0e",x"5d"),
   801 => (x"49",x"a6",x"c4",x"8e"),
   802 => (x"a6",x"cc",x"79",x"c1"),
   803 => (x"c0",x"79",x"c0",x"49"),
   804 => (x"d2",x"4a",x"66",x"f8"),
   805 => (x"c1",x"48",x"72",x"32"),
   806 => (x"58",x"a6",x"d4",x"88"),
   807 => (x"4c",x"f3",x"c2",x"c3"),
   808 => (x"00",x"0e",x"2a",x"27"),
   809 => (x"51",x"27",x"1e",x"00"),
   810 => (x"0f",x"00",x"00",x"01"),
   811 => (x"a6",x"c8",x"86",x"c4"),
   812 => (x"79",x"fe",x"c1",x"49"),
   813 => (x"c0",x"49",x"a6",x"d4"),
   814 => (x"1e",x"ee",x"c0",x"79"),
   815 => (x"00",x"00",x"50",x"27"),
   816 => (x"86",x"c4",x"0f",x"00"),
   817 => (x"79",x"74",x"49",x"76"),
   818 => (x"4b",x"74",x"4d",x"c0"),
   819 => (x"ff",x"ff",x"ff",x"c3"),
   820 => (x"4a",x"66",x"d4",x"9b"),
   821 => (x"92",x"c4",x"ba",x"73"),
   822 => (x"f4",x"c0",x"4a",x"72"),
   823 => (x"7a",x"73",x"82",x"66"),
   824 => (x"4a",x"74",x"34",x"c1"),
   825 => (x"c0",x"c0",x"c0",x"d0"),
   826 => (x"02",x"9a",x"72",x"9a"),
   827 => (x"c1",x"87",x"c2",x"c0"),
   828 => (x"c8",x"4a",x"74",x"b4"),
   829 => (x"9a",x"c0",x"c0",x"c0"),
   830 => (x"c0",x"02",x"9a",x"72"),
   831 => (x"bc",x"c1",x"87",x"c2"),
   832 => (x"c0",x"c1",x"85",x"c1"),
   833 => (x"ad",x"b7",x"c0",x"c0"),
   834 => (x"87",x"fe",x"fe",x"04"),
   835 => (x"4d",x"c0",x"4c",x"6e"),
   836 => (x"ff",x"c3",x"4a",x"74"),
   837 => (x"d8",x"9a",x"ff",x"ff"),
   838 => (x"79",x"72",x"49",x"a6"),
   839 => (x"72",x"49",x"a6",x"dc"),
   840 => (x"d4",x"4b",x"72",x"79"),
   841 => (x"93",x"c4",x"bb",x"66"),
   842 => (x"f4",x"c0",x"4b",x"73"),
   843 => (x"49",x"76",x"83",x"66"),
   844 => (x"49",x"6e",x"79",x"6b"),
   845 => (x"c0",x"02",x"a9",x"72"),
   846 => (x"a6",x"c4",x"87",x"fa"),
   847 => (x"cc",x"79",x"c0",x"49"),
   848 => (x"f0",x"27",x"1e",x"66"),
   849 => (x"1e",x"00",x"00",x"0d"),
   850 => (x"00",x"01",x"51",x"27"),
   851 => (x"86",x"c8",x"0f",x"00"),
   852 => (x"66",x"dc",x"1e",x"6e"),
   853 => (x"66",x"e4",x"c0",x"1e"),
   854 => (x"ba",x"66",x"dc",x"4a"),
   855 => (x"02",x"27",x"1e",x"72"),
   856 => (x"1e",x"00",x"00",x"0e"),
   857 => (x"00",x"01",x"51",x"27"),
   858 => (x"86",x"d0",x"0f",x"00"),
   859 => (x"c0",x"49",x"a6",x"cc"),
   860 => (x"87",x"c8",x"c0",x"79"),
   861 => (x"c1",x"48",x"66",x"cc"),
   862 => (x"58",x"a6",x"d0",x"80"),
   863 => (x"4a",x"74",x"34",x"c1"),
   864 => (x"c0",x"c0",x"c0",x"d0"),
   865 => (x"02",x"9a",x"72",x"9a"),
   866 => (x"c1",x"87",x"c2",x"c0"),
   867 => (x"c8",x"4a",x"74",x"b4"),
   868 => (x"9a",x"c0",x"c0",x"c0"),
   869 => (x"c0",x"02",x"9a",x"72"),
   870 => (x"bc",x"c1",x"87",x"c2"),
   871 => (x"c0",x"c1",x"85",x"c1"),
   872 => (x"ad",x"b7",x"c0",x"c0"),
   873 => (x"87",x"e8",x"fd",x"04"),
   874 => (x"4a",x"74",x"34",x"c1"),
   875 => (x"c0",x"c0",x"c0",x"d0"),
   876 => (x"02",x"9a",x"72",x"9a"),
   877 => (x"c1",x"87",x"c2",x"c0"),
   878 => (x"c8",x"4a",x"74",x"b4"),
   879 => (x"9a",x"c0",x"c0",x"c0"),
   880 => (x"c0",x"02",x"9a",x"72"),
   881 => (x"bc",x"c1",x"87",x"c2"),
   882 => (x"c1",x"48",x"66",x"c8"),
   883 => (x"58",x"a6",x"cc",x"88"),
   884 => (x"fb",x"05",x"66",x"c8"),
   885 => (x"1e",x"ca",x"87",x"de"),
   886 => (x"00",x"00",x"50",x"27"),
   887 => (x"86",x"c4",x"0f",x"00"),
   888 => (x"c0",x"48",x"66",x"c4"),
   889 => (x"4d",x"26",x"86",x"e0"),
   890 => (x"4b",x"26",x"4c",x"26"),
   891 => (x"4f",x"26",x"4a",x"26"),
   892 => (x"64",x"25",x"78",x"30"),
   893 => (x"6f",x"6f",x"67",x"20"),
   894 => (x"65",x"72",x"20",x"64"),
   895 => (x"2c",x"73",x"64",x"61"),
   896 => (x"72",x"45",x"00",x"20"),
   897 => (x"20",x"72",x"6f",x"72"),
   898 => (x"30",x"20",x"74",x"61"),
   899 => (x"2c",x"64",x"25",x"78"),
   900 => (x"70",x"78",x"65",x"20"),
   901 => (x"65",x"74",x"63",x"65"),
   902 => (x"78",x"30",x"20",x"64"),
   903 => (x"20",x"2c",x"64",x"25"),
   904 => (x"20",x"74",x"6f",x"67"),
   905 => (x"64",x"25",x"78",x"30"),
   906 => (x"68",x"43",x"00",x"0a"),
   907 => (x"69",x"6b",x"63",x"65"),
   908 => (x"6d",x"20",x"67",x"6e"),
   909 => (x"72",x"6f",x"6d",x"65"),
   910 => (x"5e",x"0e",x"00",x"79"),
   911 => (x"5d",x"5c",x"5b",x"5a"),
   912 => (x"c8",x"8e",x"d4",x"0e"),
   913 => (x"79",x"c1",x"49",x"a6"),
   914 => (x"ec",x"c0",x"4d",x"c0"),
   915 => (x"32",x"d2",x"4a",x"66"),
   916 => (x"88",x"c1",x"48",x"72"),
   917 => (x"c3",x"58",x"a6",x"d0"),
   918 => (x"27",x"4b",x"f3",x"c2"),
   919 => (x"00",x"00",x"0f",x"90"),
   920 => (x"01",x"51",x"27",x"1e"),
   921 => (x"c4",x"0f",x"00",x"00"),
   922 => (x"c3",x"49",x"76",x"86"),
   923 => (x"c0",x"79",x"f3",x"c2"),
   924 => (x"ac",x"66",x"cc",x"4c"),
   925 => (x"87",x"f5",x"c0",x"03"),
   926 => (x"92",x"c4",x"4a",x"74"),
   927 => (x"e8",x"c0",x"4a",x"72"),
   928 => (x"7a",x"73",x"82",x"66"),
   929 => (x"4a",x"73",x"33",x"c1"),
   930 => (x"c0",x"c0",x"c0",x"d0"),
   931 => (x"02",x"9a",x"72",x"9a"),
   932 => (x"c1",x"87",x"c2",x"c0"),
   933 => (x"c8",x"4a",x"73",x"b3"),
   934 => (x"9a",x"c0",x"c0",x"c0"),
   935 => (x"c0",x"02",x"9a",x"72"),
   936 => (x"bb",x"c1",x"87",x"c2"),
   937 => (x"66",x"cc",x"84",x"c1"),
   938 => (x"cb",x"ff",x"04",x"ac"),
   939 => (x"c0",x"4b",x"6e",x"87"),
   940 => (x"ac",x"66",x"cc",x"4c"),
   941 => (x"87",x"f9",x"c1",x"03"),
   942 => (x"73",x"49",x"a6",x"c4"),
   943 => (x"c4",x"4a",x"74",x"79"),
   944 => (x"c0",x"4a",x"72",x"92"),
   945 => (x"76",x"82",x"66",x"e8"),
   946 => (x"6e",x"79",x"6a",x"49"),
   947 => (x"02",x"a9",x"73",x"49"),
   948 => (x"c8",x"87",x"f3",x"c0"),
   949 => (x"79",x"c0",x"49",x"a6"),
   950 => (x"4a",x"27",x"1e",x"75"),
   951 => (x"1e",x"00",x"00",x"0f"),
   952 => (x"00",x"01",x"51",x"27"),
   953 => (x"86",x"c8",x"0f",x"00"),
   954 => (x"c4",x"1e",x"66",x"d0"),
   955 => (x"66",x"cc",x"1e",x"66"),
   956 => (x"27",x"1e",x"74",x"1e"),
   957 => (x"00",x"00",x"0f",x"5c"),
   958 => (x"01",x"51",x"27",x"1e"),
   959 => (x"d4",x"0f",x"00",x"00"),
   960 => (x"c0",x"4d",x"c0",x"86"),
   961 => (x"85",x"c1",x"87",x"c2"),
   962 => (x"4a",x"73",x"33",x"c1"),
   963 => (x"c0",x"c0",x"c0",x"d0"),
   964 => (x"02",x"9a",x"72",x"9a"),
   965 => (x"c1",x"87",x"c2",x"c0"),
   966 => (x"c8",x"4a",x"73",x"b3"),
   967 => (x"9a",x"c0",x"c0",x"c0"),
   968 => (x"c0",x"02",x"9a",x"72"),
   969 => (x"bb",x"c1",x"87",x"c2"),
   970 => (x"66",x"cc",x"84",x"c1"),
   971 => (x"c7",x"fe",x"04",x"ac"),
   972 => (x"27",x"1e",x"ca",x"87"),
   973 => (x"00",x"00",x"00",x"50"),
   974 => (x"c8",x"86",x"c4",x"0f"),
   975 => (x"86",x"d4",x"48",x"66"),
   976 => (x"4c",x"26",x"4d",x"26"),
   977 => (x"4a",x"26",x"4b",x"26"),
   978 => (x"78",x"30",x"4f",x"26"),
   979 => (x"67",x"20",x"64",x"25"),
   980 => (x"20",x"64",x"6f",x"6f"),
   981 => (x"64",x"61",x"65",x"72"),
   982 => (x"00",x"20",x"2c",x"73"),
   983 => (x"6f",x"72",x"72",x"45"),
   984 => (x"74",x"61",x"20",x"72"),
   985 => (x"25",x"78",x"30",x"20"),
   986 => (x"65",x"20",x"2c",x"64"),
   987 => (x"63",x"65",x"70",x"78"),
   988 => (x"20",x"64",x"65",x"74"),
   989 => (x"64",x"25",x"78",x"30"),
   990 => (x"6f",x"67",x"20",x"2c"),
   991 => (x"78",x"30",x"20",x"74"),
   992 => (x"6f",x"20",x"64",x"25"),
   993 => (x"6f",x"72",x"20",x"6e"),
   994 => (x"20",x"64",x"6e",x"75"),
   995 => (x"00",x"0a",x"64",x"25"),
   996 => (x"65",x"6e",x"69",x"4c"),
   997 => (x"6d",x"20",x"72",x"61"),
   998 => (x"72",x"6f",x"6d",x"65"),
   999 => (x"68",x"63",x"20",x"79"),
  1000 => (x"00",x"6b",x"63",x"65"),
  1001 => (x"5b",x"5a",x"5e",x"0e"),
  1002 => (x"d4",x"0e",x"5d",x"5c"),
  1003 => (x"ea",x"d5",x"c1",x"8e"),
  1004 => (x"4d",x"fb",x"d2",x"e4"),
  1005 => (x"79",x"c1",x"49",x"76"),
  1006 => (x"a6",x"c4",x"4b",x"c0"),
  1007 => (x"79",x"c0",x"c1",x"49"),
  1008 => (x"e8",x"c0",x"4c",x"c1"),
  1009 => (x"79",x"75",x"49",x"66"),
  1010 => (x"c1",x"49",x"a6",x"c8"),
  1011 => (x"49",x"a6",x"cc",x"79"),
  1012 => (x"a6",x"d0",x"79",x"c1"),
  1013 => (x"cc",x"79",x"c1",x"49"),
  1014 => (x"b2",x"74",x"4a",x"66"),
  1015 => (x"4a",x"72",x"92",x"c4"),
  1016 => (x"82",x"66",x"e8",x"c0"),
  1017 => (x"66",x"cc",x"7a",x"75"),
  1018 => (x"d0",x"30",x"c1",x"48"),
  1019 => (x"66",x"d0",x"58",x"a6"),
  1020 => (x"d4",x"80",x"c1",x"48"),
  1021 => (x"66",x"d0",x"58",x"a6"),
  1022 => (x"a9",x"b7",x"d9",x"49"),
  1023 => (x"87",x"d7",x"ff",x"04"),
  1024 => (x"66",x"c8",x"34",x"c1"),
  1025 => (x"cc",x"80",x"c1",x"48"),
  1026 => (x"66",x"c8",x"58",x"a6"),
  1027 => (x"a9",x"b7",x"d9",x"49"),
  1028 => (x"87",x"f9",x"fe",x"04"),
  1029 => (x"1e",x"66",x"ec",x"c0"),
  1030 => (x"1e",x"66",x"ec",x"c0"),
  1031 => (x"00",x"02",x"94",x"27"),
  1032 => (x"86",x"c8",x"0f",x"00"),
  1033 => (x"e8",x"c0",x"4c",x"c1"),
  1034 => (x"f8",x"f0",x"49",x"66"),
  1035 => (x"79",x"c3",x"cb",x"dd"),
  1036 => (x"c1",x"49",x"a6",x"c8"),
  1037 => (x"c4",x"4a",x"74",x"79"),
  1038 => (x"c0",x"4a",x"72",x"92"),
  1039 => (x"6a",x"82",x"66",x"e8"),
  1040 => (x"dd",x"f8",x"f0",x"49"),
  1041 => (x"05",x"a9",x"c3",x"cb"),
  1042 => (x"73",x"87",x"c7",x"c0"),
  1043 => (x"c0",x"b3",x"74",x"4b"),
  1044 => (x"4a",x"74",x"87",x"f7"),
  1045 => (x"4a",x"72",x"92",x"c4"),
  1046 => (x"82",x"66",x"e8",x"c0"),
  1047 => (x"b7",x"75",x"49",x"6a"),
  1048 => (x"e4",x"c0",x"02",x"a9"),
  1049 => (x"c0",x"49",x"76",x"87"),
  1050 => (x"c4",x"4a",x"74",x"79"),
  1051 => (x"c0",x"4a",x"72",x"92"),
  1052 => (x"6a",x"82",x"66",x"e8"),
  1053 => (x"c2",x"4a",x"74",x"1e"),
  1054 => (x"27",x"1e",x"72",x"32"),
  1055 => (x"00",x"00",x"11",x"2c"),
  1056 => (x"01",x"51",x"27",x"1e"),
  1057 => (x"cc",x"0f",x"00",x"00"),
  1058 => (x"c8",x"34",x"c1",x"86"),
  1059 => (x"80",x"c1",x"48",x"66"),
  1060 => (x"c8",x"58",x"a6",x"cc"),
  1061 => (x"b7",x"d9",x"49",x"66"),
  1062 => (x"d8",x"fe",x"04",x"a9"),
  1063 => (x"73",x"33",x"c2",x"87"),
  1064 => (x"e7",x"c1",x"02",x"9b"),
  1065 => (x"27",x"1e",x"73",x"87"),
  1066 => (x"00",x"00",x"11",x"4b"),
  1067 => (x"01",x"51",x"27",x"1e"),
  1068 => (x"c8",x"0f",x"00",x"00"),
  1069 => (x"02",x"9b",x"73",x"86"),
  1070 => (x"73",x"87",x"ec",x"c0"),
  1071 => (x"c0",x"c0",x"c2",x"4a"),
  1072 => (x"72",x"9a",x"c0",x"c0"),
  1073 => (x"c4",x"c0",x"05",x"9a"),
  1074 => (x"c0",x"49",x"76",x"87"),
  1075 => (x"c1",x"4a",x"73",x"79"),
  1076 => (x"c3",x"4b",x"72",x"32"),
  1077 => (x"ff",x"ff",x"ff",x"ff"),
  1078 => (x"48",x"66",x"c4",x"9b"),
  1079 => (x"a6",x"c8",x"28",x"c1"),
  1080 => (x"05",x"9b",x"73",x"58"),
  1081 => (x"6e",x"87",x"d4",x"ff"),
  1082 => (x"87",x"db",x"c0",x"02"),
  1083 => (x"c1",x"49",x"66",x"c4"),
  1084 => (x"c0",x"03",x"a9",x"c0"),
  1085 => (x"62",x"27",x"87",x"d1"),
  1086 => (x"1e",x"00",x"00",x"11"),
  1087 => (x"00",x"01",x"51",x"27"),
  1088 => (x"86",x"c4",x"0f",x"00"),
  1089 => (x"c4",x"87",x"c5",x"c0"),
  1090 => (x"79",x"c1",x"49",x"a6"),
  1091 => (x"27",x"1e",x"66",x"c4"),
  1092 => (x"00",x"00",x"11",x"ac"),
  1093 => (x"01",x"51",x"27",x"1e"),
  1094 => (x"c8",x"0f",x"00",x"00"),
  1095 => (x"48",x"66",x"c4",x"86"),
  1096 => (x"4d",x"26",x"86",x"d4"),
  1097 => (x"4b",x"26",x"4c",x"26"),
  1098 => (x"4f",x"26",x"4a",x"26"),
  1099 => (x"20",x"64",x"61",x"42"),
  1100 => (x"61",x"74",x"61",x"64"),
  1101 => (x"75",x"6f",x"66",x"20"),
  1102 => (x"61",x"20",x"64",x"6e"),
  1103 => (x"78",x"30",x"20",x"74"),
  1104 => (x"28",x"20",x"64",x"25"),
  1105 => (x"64",x"25",x"78",x"30"),
  1106 => (x"41",x"00",x"0a",x"29"),
  1107 => (x"73",x"61",x"69",x"6c"),
  1108 => (x"66",x"20",x"73",x"65"),
  1109 => (x"64",x"6e",x"75",x"6f"),
  1110 => (x"20",x"74",x"61",x"20"),
  1111 => (x"64",x"25",x"78",x"30"),
  1112 => (x"41",x"28",x"00",x"0a"),
  1113 => (x"73",x"61",x"69",x"6c"),
  1114 => (x"70",x"20",x"73",x"65"),
  1115 => (x"61",x"62",x"6f",x"72"),
  1116 => (x"20",x"79",x"6c",x"62"),
  1117 => (x"70",x"6d",x"69",x"73"),
  1118 => (x"69",x"20",x"79",x"6c"),
  1119 => (x"63",x"69",x"64",x"6e"),
  1120 => (x"20",x"65",x"74",x"61"),
  1121 => (x"74",x"61",x"68",x"74"),
  1122 => (x"4d",x"41",x"52",x"20"),
  1123 => (x"20",x"73",x"69",x"0a"),
  1124 => (x"6c",x"61",x"6d",x"73"),
  1125 => (x"20",x"72",x"65",x"6c"),
  1126 => (x"6e",x"61",x"68",x"74"),
  1127 => (x"20",x"34",x"36",x"20"),
  1128 => (x"61",x"67",x"65",x"6d"),
  1129 => (x"65",x"74",x"79",x"62"),
  1130 => (x"00",x"0a",x"29",x"73"),
  1131 => (x"41",x"52",x"44",x"53"),
  1132 => (x"69",x"73",x"20",x"4d"),
  1133 => (x"28",x"20",x"65",x"7a"),
  1134 => (x"75",x"73",x"73",x"61"),
  1135 => (x"67",x"6e",x"69",x"6d"),
  1136 => (x"20",x"6f",x"6e",x"20"),
  1137 => (x"72",x"64",x"64",x"61"),
  1138 => (x"20",x"73",x"73",x"65"),
  1139 => (x"6c",x"75",x"61",x"66"),
  1140 => (x"20",x"29",x"73",x"74"),
  1141 => (x"30",x"20",x"73",x"69"),
  1142 => (x"20",x"64",x"25",x"78"),
  1143 => (x"61",x"67",x"65",x"6d"),
  1144 => (x"65",x"74",x"79",x"62"),
  1145 => (x"0e",x"00",x"0a",x"73"),
  1146 => (x"5c",x"5b",x"5a",x"5e"),
  1147 => (x"dd",x"c3",x"0e",x"5d"),
  1148 => (x"c0",x"fc",x"ef",x"fb"),
  1149 => (x"ea",x"d9",x"c2",x"4d"),
  1150 => (x"4c",x"cc",x"ef",x"eb"),
  1151 => (x"d1",x"4b",x"66",x"d4"),
  1152 => (x"c4",x"cd",x"e3",x"c8"),
  1153 => (x"c4",x"4a",x"73",x"7b"),
  1154 => (x"d9",x"d5",x"c1",x"82"),
  1155 => (x"7a",x"c8",x"de",x"e7"),
  1156 => (x"82",x"c8",x"4a",x"73"),
  1157 => (x"4a",x"73",x"7a",x"74"),
  1158 => (x"7a",x"75",x"82",x"cc"),
  1159 => (x"c8",x"d1",x"49",x"6b"),
  1160 => (x"b7",x"c4",x"cd",x"e3"),
  1161 => (x"d0",x"c0",x"02",x"a9"),
  1162 => (x"27",x"1e",x"6b",x"87"),
  1163 => (x"00",x"00",x"12",x"ab"),
  1164 => (x"01",x"51",x"27",x"1e"),
  1165 => (x"c8",x"0f",x"00",x"00"),
  1166 => (x"c4",x"4a",x"73",x"86"),
  1167 => (x"c1",x"49",x"6a",x"82"),
  1168 => (x"de",x"e7",x"d9",x"d5"),
  1169 => (x"02",x"a9",x"b7",x"c8"),
  1170 => (x"73",x"87",x"d4",x"c0"),
  1171 => (x"6a",x"82",x"c4",x"4a"),
  1172 => (x"12",x"e4",x"27",x"1e"),
  1173 => (x"27",x"1e",x"00",x"00"),
  1174 => (x"00",x"00",x"01",x"51"),
  1175 => (x"73",x"86",x"c8",x"0f"),
  1176 => (x"6a",x"82",x"c8",x"4a"),
  1177 => (x"02",x"a9",x"74",x"49"),
  1178 => (x"73",x"87",x"d4",x"c0"),
  1179 => (x"6a",x"82",x"c8",x"4a"),
  1180 => (x"13",x"1d",x"27",x"1e"),
  1181 => (x"27",x"1e",x"00",x"00"),
  1182 => (x"00",x"00",x"01",x"51"),
  1183 => (x"73",x"86",x"c8",x"0f"),
  1184 => (x"6a",x"82",x"cc",x"4a"),
  1185 => (x"02",x"a9",x"75",x"49"),
  1186 => (x"73",x"87",x"d4",x"c0"),
  1187 => (x"6a",x"82",x"cc",x"4a"),
  1188 => (x"13",x"56",x"27",x"1e"),
  1189 => (x"27",x"1e",x"00",x"00"),
  1190 => (x"00",x"00",x"01",x"51"),
  1191 => (x"c1",x"86",x"c8",x"0f"),
  1192 => (x"26",x"4d",x"26",x"48"),
  1193 => (x"26",x"4b",x"26",x"4c"),
  1194 => (x"53",x"4f",x"26",x"4a"),
  1195 => (x"6c",x"70",x"6d",x"69"),
  1196 => (x"68",x"63",x"20",x"65"),
  1197 => (x"20",x"6b",x"63",x"65"),
  1198 => (x"6c",x"69",x"61",x"66"),
  1199 => (x"61",x"20",x"64",x"65"),
  1200 => (x"20",x"30",x"20",x"74"),
  1201 => (x"74",x"6f",x"67",x"28"),
  1202 => (x"2c",x"64",x"25",x"20"),
  1203 => (x"70",x"78",x"65",x"20"),
  1204 => (x"65",x"74",x"63",x"65"),
  1205 => (x"78",x"30",x"20",x"64"),
  1206 => (x"32",x"32",x"31",x"31"),
  1207 => (x"34",x"34",x"33",x"33"),
  1208 => (x"00",x"0a",x"29",x"29"),
  1209 => (x"70",x"6d",x"69",x"53"),
  1210 => (x"63",x"20",x"65",x"6c"),
  1211 => (x"6b",x"63",x"65",x"68"),
  1212 => (x"69",x"61",x"66",x"20"),
  1213 => (x"20",x"64",x"65",x"6c"),
  1214 => (x"31",x"20",x"74",x"61"),
  1215 => (x"6f",x"67",x"28",x"20"),
  1216 => (x"64",x"25",x"20",x"74"),
  1217 => (x"78",x"65",x"20",x"2c"),
  1218 => (x"74",x"63",x"65",x"70"),
  1219 => (x"30",x"20",x"64",x"65"),
  1220 => (x"36",x"35",x"35",x"78"),
  1221 => (x"38",x"37",x"37",x"36"),
  1222 => (x"0a",x"29",x"29",x"38"),
  1223 => (x"6d",x"69",x"53",x"00"),
  1224 => (x"20",x"65",x"6c",x"70"),
  1225 => (x"63",x"65",x"68",x"63"),
  1226 => (x"61",x"66",x"20",x"6b"),
  1227 => (x"64",x"65",x"6c",x"69"),
  1228 => (x"20",x"74",x"61",x"20"),
  1229 => (x"67",x"28",x"20",x"32"),
  1230 => (x"25",x"20",x"74",x"6f"),
  1231 => (x"65",x"20",x"2c",x"64"),
  1232 => (x"63",x"65",x"70",x"78"),
  1233 => (x"20",x"64",x"65",x"74"),
  1234 => (x"39",x"39",x"78",x"30"),
  1235 => (x"62",x"62",x"61",x"61"),
  1236 => (x"29",x"29",x"63",x"63"),
  1237 => (x"69",x"53",x"00",x"0a"),
  1238 => (x"65",x"6c",x"70",x"6d"),
  1239 => (x"65",x"68",x"63",x"20"),
  1240 => (x"66",x"20",x"6b",x"63"),
  1241 => (x"65",x"6c",x"69",x"61"),
  1242 => (x"74",x"61",x"20",x"64"),
  1243 => (x"28",x"20",x"33",x"20"),
  1244 => (x"20",x"74",x"6f",x"67"),
  1245 => (x"20",x"2c",x"64",x"25"),
  1246 => (x"65",x"70",x"78",x"65"),
  1247 => (x"64",x"65",x"74",x"63"),
  1248 => (x"64",x"78",x"30",x"20"),
  1249 => (x"66",x"65",x"65",x"64"),
  1250 => (x"29",x"30",x"30",x"66"),
  1251 => (x"0e",x"00",x"0a",x"29"),
  1252 => (x"5c",x"5b",x"5a",x"5e"),
  1253 => (x"c0",x"c1",x"0e",x"5d"),
  1254 => (x"e0",x"c0",x"4d",x"c0"),
  1255 => (x"c0",x"c0",x"c0",x"c0"),
  1256 => (x"73",x"1e",x"75",x"4b"),
  1257 => (x"11",x"e7",x"27",x"1e"),
  1258 => (x"c8",x"0f",x"00",x"00"),
  1259 => (x"72",x"4a",x"70",x"86"),
  1260 => (x"ce",x"c0",x"02",x"9a"),
  1261 => (x"14",x"7a",x"27",x"87"),
  1262 => (x"27",x"1e",x"00",x"00"),
  1263 => (x"00",x"00",x"01",x"51"),
  1264 => (x"75",x"86",x"c4",x"0f"),
  1265 => (x"27",x"1e",x"73",x"1e"),
  1266 => (x"00",x"00",x"02",x"b9"),
  1267 => (x"70",x"86",x"c8",x"0f"),
  1268 => (x"02",x"9a",x"72",x"4a"),
  1269 => (x"27",x"87",x"ce",x"c0"),
  1270 => (x"00",x"00",x"14",x"90"),
  1271 => (x"01",x"51",x"27",x"1e"),
  1272 => (x"c4",x"0f",x"00",x"00"),
  1273 => (x"73",x"1e",x"75",x"86"),
  1274 => (x"03",x"55",x"27",x"1e"),
  1275 => (x"c8",x"0f",x"00",x"00"),
  1276 => (x"72",x"4a",x"70",x"86"),
  1277 => (x"ce",x"c0",x"02",x"9a"),
  1278 => (x"14",x"b2",x"27",x"87"),
  1279 => (x"27",x"1e",x"00",x"00"),
  1280 => (x"00",x"00",x"01",x"51"),
  1281 => (x"75",x"86",x"c4",x"0f"),
  1282 => (x"27",x"1e",x"73",x"1e"),
  1283 => (x"00",x"00",x"0f",x"a4"),
  1284 => (x"70",x"86",x"c8",x"0f"),
  1285 => (x"02",x"9c",x"74",x"4c"),
  1286 => (x"27",x"87",x"ce",x"c0"),
  1287 => (x"00",x"00",x"14",x"cb"),
  1288 => (x"01",x"51",x"27",x"1e"),
  1289 => (x"c4",x"0f",x"00",x"00"),
  1290 => (x"73",x"1e",x"74",x"86"),
  1291 => (x"0e",x"3a",x"27",x"1e"),
  1292 => (x"c8",x"0f",x"00",x"00"),
  1293 => (x"72",x"4a",x"70",x"86"),
  1294 => (x"ce",x"c0",x"02",x"9a"),
  1295 => (x"14",x"e2",x"27",x"87"),
  1296 => (x"27",x"1e",x"00",x"00"),
  1297 => (x"00",x"00",x"01",x"51"),
  1298 => (x"74",x"86",x"c4",x"0f"),
  1299 => (x"27",x"1e",x"73",x"1e"),
  1300 => (x"00",x"00",x"0c",x"7b"),
  1301 => (x"70",x"86",x"c8",x"0f"),
  1302 => (x"02",x"9a",x"72",x"4a"),
  1303 => (x"27",x"87",x"c2",x"fd"),
  1304 => (x"00",x"00",x"14",x"f9"),
  1305 => (x"01",x"51",x"27",x"1e"),
  1306 => (x"c4",x"0f",x"00",x"00"),
  1307 => (x"87",x"f1",x"fc",x"86"),
  1308 => (x"4c",x"26",x"4d",x"26"),
  1309 => (x"4a",x"26",x"4b",x"26"),
  1310 => (x"69",x"53",x"4f",x"26"),
  1311 => (x"65",x"6c",x"70",x"6d"),
  1312 => (x"65",x"68",x"63",x"20"),
  1313 => (x"70",x"20",x"6b",x"63"),
  1314 => (x"65",x"73",x"73",x"61"),
  1315 => (x"00",x"0a",x"2e",x"64"),
  1316 => (x"73",x"72",x"69",x"46"),
  1317 => (x"74",x"73",x"20",x"74"),
  1318 => (x"20",x"65",x"67",x"61"),
  1319 => (x"69",x"6e",x"61",x"73"),
  1320 => (x"63",x"20",x"79",x"74"),
  1321 => (x"6b",x"63",x"65",x"68"),
  1322 => (x"73",x"61",x"70",x"20"),
  1323 => (x"2e",x"64",x"65",x"73"),
  1324 => (x"79",x"42",x"00",x"0a"),
  1325 => (x"28",x"20",x"65",x"74"),
  1326 => (x"29",x"6d",x"71",x"64"),
  1327 => (x"65",x"68",x"63",x"20"),
  1328 => (x"70",x"20",x"6b",x"63"),
  1329 => (x"65",x"73",x"73",x"61"),
  1330 => (x"41",x"00",x"0a",x"64"),
  1331 => (x"65",x"72",x"64",x"64"),
  1332 => (x"63",x"20",x"73",x"73"),
  1333 => (x"6b",x"63",x"65",x"68"),
  1334 => (x"73",x"61",x"70",x"20"),
  1335 => (x"2e",x"64",x"65",x"73"),
  1336 => (x"69",x"4c",x"00",x"0a"),
  1337 => (x"72",x"61",x"65",x"6e"),
  1338 => (x"65",x"68",x"63",x"20"),
  1339 => (x"70",x"20",x"6b",x"63"),
  1340 => (x"65",x"73",x"73",x"61"),
  1341 => (x"0a",x"0a",x"2e",x"64"),
  1342 => (x"53",x"46",x"4c",x"00"),
  1343 => (x"68",x"63",x"20",x"52"),
  1344 => (x"20",x"6b",x"63",x"65"),
  1345 => (x"73",x"73",x"61",x"70"),
  1346 => (x"0a",x"2e",x"64",x"65"),
  1347 => (x"90",x"66",x"00",x"0a"),
  1348 => (x"00",x"00",x"00",x"00"),
  1349 => (x"55",x"55",x"55",x"55"),
  1350 => (x"aa",x"aa",x"aa",x"aa"),
  1351 => (x"ff",x"ff",x"ff",x"ff"),
  1352 => (x"72",x"1e",x"73",x"1e"),
  1353 => (x"87",x"d9",x"02",x"9a"),
  1354 => (x"4b",x"c1",x"48",x"c0"),
  1355 => (x"82",x"01",x"a9",x"72"),
  1356 => (x"87",x"f8",x"83",x"73"),
  1357 => (x"89",x"03",x"a9",x"72"),
  1358 => (x"c1",x"07",x"80",x"73"),
  1359 => (x"f3",x"05",x"2b",x"2a"),
  1360 => (x"26",x"4b",x"26",x"87"),
  1361 => (x"1e",x"75",x"1e",x"4f"),
  1362 => (x"a1",x"71",x"4d",x"c0"),
  1363 => (x"c1",x"b9",x"ff",x"04"),
  1364 => (x"72",x"07",x"bd",x"81"),
  1365 => (x"ba",x"ff",x"04",x"a2"),
  1366 => (x"07",x"bd",x"82",x"c1"),
  1367 => (x"9d",x"75",x"87",x"c2"),
  1368 => (x"c1",x"b8",x"ff",x"05"),
  1369 => (x"4d",x"25",x"07",x"80"),
  1370 => (x"31",x"30",x"4f",x"26"),
  1371 => (x"35",x"34",x"33",x"32"),
  1372 => (x"39",x"38",x"37",x"36"),
  1373 => (x"44",x"43",x"42",x"41"),
  1374 => (x"53",x"00",x"46",x"45"),
  1375 => (x"74",x"69",x"6e",x"61"),
  1376 => (x"68",x"63",x"20",x"79"),
  1377 => (x"20",x"6b",x"63",x"65"),
  1378 => (x"6c",x"69",x"61",x"66"),
  1379 => (x"28",x"20",x"64",x"65"),
  1380 => (x"6f",x"66",x"65",x"62"),
  1381 => (x"63",x"20",x"65",x"72"),
  1382 => (x"65",x"68",x"63",x"61"),
  1383 => (x"66",x"65",x"72",x"20"),
  1384 => (x"68",x"73",x"65",x"72"),
  1385 => (x"6e",x"6f",x"20",x"29"),
  1386 => (x"25",x"78",x"30",x"20"),
  1387 => (x"67",x"28",x"20",x"64"),
  1388 => (x"30",x"20",x"74",x"6f"),
  1389 => (x"29",x"64",x"25",x"78"),
  1390 => (x"61",x"53",x"00",x"0a"),
  1391 => (x"79",x"74",x"69",x"6e"),
  1392 => (x"65",x"68",x"63",x"20"),
  1393 => (x"66",x"20",x"6b",x"63"),
  1394 => (x"65",x"6c",x"69",x"61"),
  1395 => (x"61",x"28",x"20",x"64"),
  1396 => (x"72",x"65",x"74",x"66"),
  1397 => (x"63",x"61",x"63",x"20"),
  1398 => (x"72",x"20",x"65",x"68"),
  1399 => (x"65",x"72",x"66",x"65"),
  1400 => (x"20",x"29",x"68",x"73"),
  1401 => (x"30",x"20",x"6e",x"6f"),
  1402 => (x"20",x"64",x"25",x"78"),
  1403 => (x"74",x"6f",x"67",x"28"),
  1404 => (x"25",x"78",x"30",x"20"),
  1405 => (x"00",x"0a",x"29",x"64"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
