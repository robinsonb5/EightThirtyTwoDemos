
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"d4",x"01"),
     1 => (x"18",x"0e",x"87",x"d7"),
     2 => (x"3e",x"27",x"0e",x"1e"),
     3 => (x"0f",x"00",x"00",x"00"),
     4 => (x"80",x"ff",x"48",x"26"),
     5 => (x"27",x"4f",x"08",x"26"),
     6 => (x"00",x"00",x"00",x"23"),
     7 => (x"00",x"30",x"27",x"4f"),
     8 => (x"c2",x"4f",x"00",x"00"),
     9 => (x"27",x"4e",x"c0",x"c0"),
    10 => (x"00",x"00",x"16",x"04"),
    11 => (x"87",x"fd",x"00",x"0f"),
    12 => (x"4e",x"c0",x"f0",x"c1"),
    13 => (x"00",x"00",x"3d",x"27"),
    14 => (x"fd",x"00",x"0f",x"00"),
    15 => (x"1e",x"4f",x"4f",x"87"),
    16 => (x"ff",x"1e",x"1e",x"72"),
    17 => (x"48",x"6a",x"4a",x"c0"),
    18 => (x"c4",x"98",x"c0",x"c4"),
    19 => (x"02",x"6e",x"58",x"a6"),
    20 => (x"cc",x"87",x"f3",x"ff"),
    21 => (x"66",x"cc",x"7a",x"66"),
    22 => (x"4a",x"26",x"26",x"48"),
    23 => (x"5e",x"0e",x"4f",x"26"),
    24 => (x"5d",x"5c",x"5b",x"5a"),
    25 => (x"4b",x"66",x"d4",x"0e"),
    26 => (x"4c",x"13",x"4d",x"c0"),
    27 => (x"c0",x"02",x"9c",x"74"),
    28 => (x"4a",x"74",x"87",x"d6"),
    29 => (x"3f",x"27",x"1e",x"72"),
    30 => (x"0f",x"00",x"00",x"00"),
    31 => (x"85",x"c1",x"86",x"c4"),
    32 => (x"9c",x"74",x"4c",x"13"),
    33 => (x"87",x"ea",x"ff",x"05"),
    34 => (x"4d",x"26",x"48",x"75"),
    35 => (x"4b",x"26",x"4c",x"26"),
    36 => (x"4f",x"26",x"4a",x"26"),
    37 => (x"5b",x"5a",x"5e",x"0e"),
    38 => (x"d0",x"0e",x"5d",x"5c"),
    39 => (x"c4",x"4c",x"c0",x"8e"),
    40 => (x"79",x"c0",x"49",x"a6"),
    41 => (x"4b",x"a6",x"e8",x"c0"),
    42 => (x"4a",x"66",x"e4",x"c0"),
    43 => (x"48",x"66",x"e4",x"c0"),
    44 => (x"e8",x"c0",x"80",x"c1"),
    45 => (x"48",x"12",x"58",x"a6"),
    46 => (x"c0",x"c0",x"c0",x"c1"),
    47 => (x"c0",x"c4",x"90",x"c0"),
    48 => (x"c4",x"48",x"90",x"b7"),
    49 => (x"02",x"6e",x"58",x"a6"),
    50 => (x"c4",x"87",x"c3",x"c5"),
    51 => (x"ff",x"c3",x"02",x"66"),
    52 => (x"49",x"a6",x"c4",x"87"),
    53 => (x"4a",x"6e",x"79",x"c0"),
    54 => (x"f0",x"c0",x"49",x"6e"),
    55 => (x"c5",x"c3",x"02",x"a9"),
    56 => (x"aa",x"e3",x"c1",x"87"),
    57 => (x"87",x"c6",x"c3",x"02"),
    58 => (x"02",x"aa",x"e4",x"c1"),
    59 => (x"c1",x"87",x"e3",x"c0"),
    60 => (x"c2",x"02",x"aa",x"ec"),
    61 => (x"f0",x"c1",x"87",x"f0"),
    62 => (x"d5",x"c0",x"02",x"aa"),
    63 => (x"aa",x"f3",x"c1",x"87"),
    64 => (x"87",x"c9",x"c2",x"02"),
    65 => (x"02",x"aa",x"f5",x"c1"),
    66 => (x"c1",x"87",x"c7",x"c0"),
    67 => (x"c2",x"05",x"aa",x"f8"),
    68 => (x"83",x"c4",x"87",x"f1"),
    69 => (x"8a",x"c4",x"4a",x"73"),
    70 => (x"79",x"6a",x"49",x"76"),
    71 => (x"dc",x"c1",x"02",x"6e"),
    72 => (x"49",x"a6",x"c8",x"87"),
    73 => (x"a6",x"cc",x"79",x"c0"),
    74 => (x"6e",x"79",x"c0",x"49"),
    75 => (x"2a",x"b7",x"dc",x"4a"),
    76 => (x"9d",x"cf",x"4d",x"72"),
    77 => (x"30",x"c4",x"48",x"6e"),
    78 => (x"75",x"58",x"a6",x"c4"),
    79 => (x"c5",x"c0",x"02",x"9d"),
    80 => (x"49",x"a6",x"c8",x"87"),
    81 => (x"b7",x"c9",x"79",x"c1"),
    82 => (x"c6",x"c0",x"06",x"ad"),
    83 => (x"85",x"f7",x"c0",x"87"),
    84 => (x"c0",x"87",x"c3",x"c0"),
    85 => (x"66",x"c8",x"85",x"f0"),
    86 => (x"87",x"cc",x"c0",x"02"),
    87 => (x"3f",x"27",x"1e",x"75"),
    88 => (x"0f",x"00",x"00",x"00"),
    89 => (x"84",x"c1",x"86",x"c4"),
    90 => (x"c1",x"48",x"66",x"cc"),
    91 => (x"58",x"a6",x"d0",x"80"),
    92 => (x"c8",x"49",x"66",x"cc"),
    93 => (x"fe",x"04",x"a9",x"b7"),
    94 => (x"ee",x"c1",x"87",x"f1"),
    95 => (x"1e",x"f0",x"c0",x"87"),
    96 => (x"00",x"00",x"3f",x"27"),
    97 => (x"86",x"c4",x"0f",x"00"),
    98 => (x"de",x"c1",x"84",x"c1"),
    99 => (x"73",x"83",x"c4",x"87"),
   100 => (x"6a",x"8a",x"c4",x"4a"),
   101 => (x"00",x"5e",x"27",x"1e"),
   102 => (x"c4",x"0f",x"00",x"00"),
   103 => (x"74",x"4a",x"70",x"86"),
   104 => (x"c1",x"84",x"72",x"4c"),
   105 => (x"a6",x"c4",x"87",x"c5"),
   106 => (x"c0",x"79",x"c1",x"49"),
   107 => (x"83",x"c4",x"87",x"fd"),
   108 => (x"8a",x"c4",x"4a",x"73"),
   109 => (x"3f",x"27",x"1e",x"6a"),
   110 => (x"0f",x"00",x"00",x"00"),
   111 => (x"84",x"c1",x"86",x"c4"),
   112 => (x"6e",x"87",x"e8",x"c0"),
   113 => (x"00",x"3f",x"27",x"1e"),
   114 => (x"c4",x"0f",x"00",x"00"),
   115 => (x"87",x"db",x"c0",x"86"),
   116 => (x"e5",x"c0",x"49",x"6e"),
   117 => (x"c8",x"c0",x"05",x"a9"),
   118 => (x"49",x"a6",x"c4",x"87"),
   119 => (x"ca",x"c0",x"79",x"c1"),
   120 => (x"27",x"1e",x"6e",x"87"),
   121 => (x"00",x"00",x"00",x"3f"),
   122 => (x"c0",x"86",x"c4",x"0f"),
   123 => (x"c0",x"4a",x"66",x"e4"),
   124 => (x"c1",x"48",x"66",x"e4"),
   125 => (x"a6",x"e8",x"c0",x"80"),
   126 => (x"c1",x"48",x"12",x"58"),
   127 => (x"c0",x"c0",x"c0",x"c0"),
   128 => (x"b7",x"c0",x"c4",x"90"),
   129 => (x"a6",x"c4",x"48",x"90"),
   130 => (x"fa",x"05",x"6e",x"58"),
   131 => (x"48",x"74",x"87",x"fd"),
   132 => (x"4d",x"26",x"86",x"d0"),
   133 => (x"4b",x"26",x"4c",x"26"),
   134 => (x"4f",x"26",x"4a",x"26"),
   135 => (x"00",x"00",x"00",x"00"),
   136 => (x"ff",x"1e",x"75",x"1e"),
   137 => (x"ff",x"c3",x"4d",x"d4"),
   138 => (x"48",x"6d",x"7d",x"49"),
   139 => (x"7d",x"71",x"38",x"c8"),
   140 => (x"38",x"c8",x"b0",x"6d"),
   141 => (x"b0",x"6d",x"7d",x"71"),
   142 => (x"7d",x"71",x"38",x"c8"),
   143 => (x"38",x"c8",x"b0",x"6d"),
   144 => (x"4f",x"26",x"4d",x"26"),
   145 => (x"ff",x"1e",x"75",x"1e"),
   146 => (x"ff",x"c3",x"4d",x"d4"),
   147 => (x"48",x"6d",x"7d",x"49"),
   148 => (x"7d",x"71",x"30",x"c8"),
   149 => (x"30",x"c8",x"b0",x"6d"),
   150 => (x"b0",x"6d",x"7d",x"71"),
   151 => (x"7d",x"71",x"30",x"c8"),
   152 => (x"4d",x"26",x"b0",x"6d"),
   153 => (x"75",x"1e",x"4f",x"26"),
   154 => (x"4d",x"d4",x"ff",x"1e"),
   155 => (x"c8",x"49",x"66",x"cc"),
   156 => (x"fe",x"7d",x"48",x"66"),
   157 => (x"c9",x"02",x"67",x"e6"),
   158 => (x"39",x"d8",x"07",x"31"),
   159 => (x"39",x"09",x"7d",x"09"),
   160 => (x"39",x"09",x"7d",x"09"),
   161 => (x"39",x"09",x"7d",x"09"),
   162 => (x"38",x"d0",x"7d",x"09"),
   163 => (x"f1",x"c9",x"7d",x"70"),
   164 => (x"ff",x"c3",x"49",x"c0"),
   165 => (x"a8",x"08",x"6d",x"48"),
   166 => (x"08",x"87",x"c7",x"05"),
   167 => (x"05",x"89",x"c1",x"7d"),
   168 => (x"4d",x"26",x"87",x"f3"),
   169 => (x"ff",x"1e",x"4f",x"26"),
   170 => (x"c8",x"c3",x"49",x"d4"),
   171 => (x"80",x"79",x"ff",x"48"),
   172 => (x"26",x"87",x"fa",x"05"),
   173 => (x"5a",x"5e",x"0e",x"4f"),
   174 => (x"0e",x"5d",x"5c",x"5b"),
   175 => (x"c1",x"f0",x"ff",x"c0"),
   176 => (x"c0",x"c1",x"4d",x"f7"),
   177 => (x"c0",x"c0",x"c0",x"c0"),
   178 => (x"02",x"a6",x"27",x"4b"),
   179 => (x"c4",x"0f",x"00",x"00"),
   180 => (x"c0",x"4c",x"df",x"f8"),
   181 => (x"27",x"1e",x"75",x"1e"),
   182 => (x"00",x"00",x"02",x"66"),
   183 => (x"70",x"86",x"c8",x"0f"),
   184 => (x"aa",x"b7",x"c1",x"4a"),
   185 => (x"87",x"ef",x"c0",x"05"),
   186 => (x"c3",x"49",x"d4",x"ff"),
   187 => (x"1e",x"73",x"79",x"ff"),
   188 => (x"c1",x"f0",x"e1",x"c0"),
   189 => (x"66",x"27",x"1e",x"e9"),
   190 => (x"0f",x"00",x"00",x"02"),
   191 => (x"4a",x"70",x"86",x"c8"),
   192 => (x"c0",x"05",x"9a",x"72"),
   193 => (x"d4",x"ff",x"87",x"cb"),
   194 => (x"79",x"ff",x"c3",x"49"),
   195 => (x"d0",x"c0",x"48",x"c1"),
   196 => (x"02",x"a6",x"27",x"87"),
   197 => (x"c1",x"0f",x"00",x"00"),
   198 => (x"05",x"9c",x"74",x"8c"),
   199 => (x"c0",x"87",x"f4",x"fe"),
   200 => (x"26",x"4d",x"26",x"48"),
   201 => (x"26",x"4b",x"26",x"4c"),
   202 => (x"0e",x"4f",x"26",x"4a"),
   203 => (x"5c",x"5b",x"5a",x"5e"),
   204 => (x"f0",x"ff",x"c0",x"0e"),
   205 => (x"ff",x"4c",x"c1",x"c1"),
   206 => (x"ff",x"c3",x"49",x"d4"),
   207 => (x"18",x"16",x"27",x"79"),
   208 => (x"27",x"1e",x"00",x"00"),
   209 => (x"00",x"00",x"00",x"5e"),
   210 => (x"d3",x"86",x"c4",x"0f"),
   211 => (x"74",x"1e",x"c0",x"4b"),
   212 => (x"02",x"66",x"27",x"1e"),
   213 => (x"c8",x"0f",x"00",x"00"),
   214 => (x"72",x"4a",x"70",x"86"),
   215 => (x"cb",x"c0",x"05",x"9a"),
   216 => (x"49",x"d4",x"ff",x"87"),
   217 => (x"c1",x"79",x"ff",x"c3"),
   218 => (x"87",x"d0",x"c0",x"48"),
   219 => (x"00",x"02",x"a6",x"27"),
   220 => (x"8b",x"c1",x"0f",x"00"),
   221 => (x"ff",x"05",x"9b",x"73"),
   222 => (x"48",x"c0",x"87",x"d3"),
   223 => (x"4b",x"26",x"4c",x"26"),
   224 => (x"4f",x"26",x"4a",x"26"),
   225 => (x"5b",x"5a",x"5e",x"0e"),
   226 => (x"1e",x"0e",x"5d",x"5c"),
   227 => (x"ff",x"4d",x"ff",x"c3"),
   228 => (x"a6",x"27",x"4c",x"d4"),
   229 => (x"0f",x"00",x"00",x"02"),
   230 => (x"c0",x"1e",x"ea",x"c6"),
   231 => (x"c8",x"c1",x"f0",x"e1"),
   232 => (x"02",x"66",x"27",x"1e"),
   233 => (x"c8",x"0f",x"00",x"00"),
   234 => (x"72",x"4a",x"70",x"86"),
   235 => (x"04",x"e3",x"27",x"1e"),
   236 => (x"27",x"1e",x"00",x"00"),
   237 => (x"00",x"00",x"00",x"94"),
   238 => (x"c1",x"86",x"c8",x"0f"),
   239 => (x"c0",x"02",x"aa",x"b7"),
   240 => (x"2b",x"27",x"87",x"cb"),
   241 => (x"0f",x"00",x"00",x"03"),
   242 => (x"c9",x"c3",x"48",x"c0"),
   243 => (x"02",x"44",x"27",x"87"),
   244 => (x"70",x"0f",x"00",x"00"),
   245 => (x"ff",x"ff",x"cf",x"4a"),
   246 => (x"b7",x"ea",x"c6",x"9a"),
   247 => (x"cb",x"c0",x"02",x"aa"),
   248 => (x"03",x"2b",x"27",x"87"),
   249 => (x"c0",x"0f",x"00",x"00"),
   250 => (x"87",x"ea",x"c2",x"48"),
   251 => (x"49",x"76",x"7c",x"75"),
   252 => (x"27",x"79",x"f1",x"c0"),
   253 => (x"00",x"00",x"02",x"b5"),
   254 => (x"72",x"4a",x"70",x"0f"),
   255 => (x"eb",x"c1",x"02",x"9a"),
   256 => (x"c0",x"1e",x"c0",x"87"),
   257 => (x"fa",x"c1",x"f0",x"ff"),
   258 => (x"02",x"66",x"27",x"1e"),
   259 => (x"c8",x"0f",x"00",x"00"),
   260 => (x"73",x"4b",x"70",x"86"),
   261 => (x"c3",x"c1",x"05",x"9b"),
   262 => (x"27",x"1e",x"73",x"87"),
   263 => (x"00",x"00",x"04",x"a1"),
   264 => (x"00",x"94",x"27",x"1e"),
   265 => (x"c8",x"0f",x"00",x"00"),
   266 => (x"6c",x"7c",x"75",x"86"),
   267 => (x"73",x"9b",x"75",x"4b"),
   268 => (x"04",x"ad",x"27",x"1e"),
   269 => (x"27",x"1e",x"00",x"00"),
   270 => (x"00",x"00",x"00",x"94"),
   271 => (x"75",x"86",x"c8",x"0f"),
   272 => (x"75",x"7c",x"75",x"7c"),
   273 => (x"73",x"7c",x"75",x"7c"),
   274 => (x"9a",x"c0",x"c1",x"4a"),
   275 => (x"c0",x"02",x"9a",x"72"),
   276 => (x"48",x"c1",x"87",x"c5"),
   277 => (x"c0",x"87",x"ff",x"c0"),
   278 => (x"87",x"fa",x"c0",x"48"),
   279 => (x"bb",x"27",x"1e",x"73"),
   280 => (x"1e",x"00",x"00",x"04"),
   281 => (x"00",x"00",x"94",x"27"),
   282 => (x"86",x"c8",x"0f",x"00"),
   283 => (x"b7",x"c2",x"49",x"6e"),
   284 => (x"d3",x"c0",x"05",x"a9"),
   285 => (x"04",x"c7",x"27",x"87"),
   286 => (x"27",x"1e",x"00",x"00"),
   287 => (x"00",x"00",x"00",x"94"),
   288 => (x"c0",x"86",x"c4",x"0f"),
   289 => (x"87",x"ce",x"c0",x"48"),
   290 => (x"88",x"c1",x"48",x"6e"),
   291 => (x"6e",x"58",x"a6",x"c4"),
   292 => (x"87",x"df",x"fd",x"05"),
   293 => (x"26",x"26",x"48",x"c0"),
   294 => (x"26",x"4c",x"26",x"4d"),
   295 => (x"26",x"4a",x"26",x"4b"),
   296 => (x"44",x"4d",x"43",x"4f"),
   297 => (x"25",x"20",x"38",x"35"),
   298 => (x"20",x"20",x"0a",x"64"),
   299 => (x"44",x"4d",x"43",x"00"),
   300 => (x"32",x"5f",x"38",x"35"),
   301 => (x"0a",x"64",x"25",x"20"),
   302 => (x"43",x"00",x"20",x"20"),
   303 => (x"38",x"35",x"44",x"4d"),
   304 => (x"0a",x"64",x"25",x"20"),
   305 => (x"53",x"00",x"20",x"20"),
   306 => (x"20",x"43",x"48",x"44"),
   307 => (x"74",x"69",x"6e",x"49"),
   308 => (x"69",x"6c",x"61",x"69"),
   309 => (x"69",x"74",x"61",x"7a"),
   310 => (x"65",x"20",x"6e",x"6f"),
   311 => (x"72",x"6f",x"72",x"72"),
   312 => (x"63",x"00",x"0a",x"21"),
   313 => (x"43",x"5f",x"64",x"6d"),
   314 => (x"20",x"38",x"44",x"4d"),
   315 => (x"70",x"73",x"65",x"72"),
   316 => (x"65",x"73",x"6e",x"6f"),
   317 => (x"64",x"25",x"20",x"3a"),
   318 => (x"5e",x"0e",x"00",x"0a"),
   319 => (x"5d",x"5c",x"5b",x"5a"),
   320 => (x"d0",x"ff",x"1e",x"0e"),
   321 => (x"c0",x"c0",x"c8",x"4c"),
   322 => (x"02",x"1c",x"27",x"4b"),
   323 => (x"c1",x"49",x"00",x"00"),
   324 => (x"06",x"17",x"27",x"79"),
   325 => (x"27",x"1e",x"00",x"00"),
   326 => (x"00",x"00",x"00",x"5e"),
   327 => (x"c7",x"86",x"c4",x"0f"),
   328 => (x"73",x"48",x"6c",x"4d"),
   329 => (x"58",x"a6",x"c4",x"98"),
   330 => (x"cc",x"c0",x"02",x"6e"),
   331 => (x"73",x"48",x"6c",x"87"),
   332 => (x"58",x"a6",x"c4",x"98"),
   333 => (x"f4",x"ff",x"05",x"6e"),
   334 => (x"27",x"7c",x"c0",x"87"),
   335 => (x"00",x"00",x"02",x"a6"),
   336 => (x"73",x"48",x"6c",x"0f"),
   337 => (x"58",x"a6",x"c4",x"98"),
   338 => (x"cc",x"c0",x"02",x"6e"),
   339 => (x"73",x"48",x"6c",x"87"),
   340 => (x"58",x"a6",x"c4",x"98"),
   341 => (x"f4",x"ff",x"05",x"6e"),
   342 => (x"c0",x"7c",x"c1",x"87"),
   343 => (x"d0",x"e5",x"c0",x"1e"),
   344 => (x"27",x"1e",x"c0",x"c1"),
   345 => (x"00",x"00",x"02",x"66"),
   346 => (x"70",x"86",x"c8",x"0f"),
   347 => (x"aa",x"b7",x"c1",x"4a"),
   348 => (x"87",x"c2",x"c0",x"05"),
   349 => (x"b7",x"c2",x"4d",x"c1"),
   350 => (x"d3",x"c0",x"05",x"ad"),
   351 => (x"06",x"12",x"27",x"87"),
   352 => (x"27",x"1e",x"00",x"00"),
   353 => (x"00",x"00",x"00",x"5e"),
   354 => (x"c0",x"86",x"c4",x"0f"),
   355 => (x"87",x"f7",x"c1",x"48"),
   356 => (x"9d",x"75",x"8d",x"c1"),
   357 => (x"87",x"c9",x"fe",x"05"),
   358 => (x"00",x"03",x"84",x"27"),
   359 => (x"20",x"27",x"0f",x"00"),
   360 => (x"58",x"00",x"00",x"02"),
   361 => (x"00",x"02",x"1c",x"27"),
   362 => (x"c0",x"05",x"bf",x"00"),
   363 => (x"1e",x"c1",x"87",x"d0"),
   364 => (x"c1",x"f0",x"ff",x"c0"),
   365 => (x"66",x"27",x"1e",x"d0"),
   366 => (x"0f",x"00",x"00",x"02"),
   367 => (x"d4",x"ff",x"86",x"c8"),
   368 => (x"79",x"ff",x"c3",x"49"),
   369 => (x"00",x"08",x"ad",x"27"),
   370 => (x"b0",x"27",x"0f",x"00"),
   371 => (x"58",x"00",x"00",x"19"),
   372 => (x"00",x"19",x"ac",x"27"),
   373 => (x"27",x"1e",x"bf",x"00"),
   374 => (x"00",x"00",x"06",x"1b"),
   375 => (x"00",x"94",x"27",x"1e"),
   376 => (x"c8",x"0f",x"00",x"00"),
   377 => (x"73",x"48",x"6c",x"86"),
   378 => (x"58",x"a6",x"c4",x"98"),
   379 => (x"cc",x"c0",x"02",x"6e"),
   380 => (x"73",x"48",x"6c",x"87"),
   381 => (x"58",x"a6",x"c4",x"98"),
   382 => (x"f4",x"ff",x"05",x"6e"),
   383 => (x"ff",x"7c",x"c0",x"87"),
   384 => (x"ff",x"c3",x"49",x"d4"),
   385 => (x"26",x"48",x"c1",x"79"),
   386 => (x"4c",x"26",x"4d",x"26"),
   387 => (x"4a",x"26",x"4b",x"26"),
   388 => (x"45",x"49",x"4f",x"26"),
   389 => (x"53",x"00",x"52",x"52"),
   390 => (x"53",x"00",x"49",x"50"),
   391 => (x"61",x"63",x"20",x"44"),
   392 => (x"73",x"20",x"64",x"72"),
   393 => (x"20",x"65",x"7a",x"69"),
   394 => (x"25",x"20",x"73",x"69"),
   395 => (x"0e",x"00",x"0a",x"64"),
   396 => (x"5c",x"5b",x"5a",x"5e"),
   397 => (x"c3",x"1e",x"0e",x"5d"),
   398 => (x"d4",x"ff",x"4d",x"ff"),
   399 => (x"ff",x"7c",x"75",x"4c"),
   400 => (x"c8",x"48",x"bf",x"d0"),
   401 => (x"c4",x"98",x"c0",x"c0"),
   402 => (x"02",x"6e",x"58",x"a6"),
   403 => (x"c8",x"87",x"d2",x"c0"),
   404 => (x"ff",x"4a",x"c0",x"c0"),
   405 => (x"72",x"48",x"bf",x"d0"),
   406 => (x"58",x"a6",x"c4",x"98"),
   407 => (x"f2",x"ff",x"05",x"6e"),
   408 => (x"49",x"d0",x"ff",x"87"),
   409 => (x"75",x"79",x"c1",x"c4"),
   410 => (x"1e",x"66",x"d8",x"7c"),
   411 => (x"c1",x"f0",x"ff",x"c0"),
   412 => (x"66",x"27",x"1e",x"d8"),
   413 => (x"0f",x"00",x"00",x"02"),
   414 => (x"4a",x"70",x"86",x"c8"),
   415 => (x"c0",x"02",x"9a",x"72"),
   416 => (x"37",x"27",x"87",x"d3"),
   417 => (x"1e",x"00",x"00",x"07"),
   418 => (x"00",x"00",x"5e",x"27"),
   419 => (x"86",x"c4",x"0f",x"00"),
   420 => (x"d7",x"c2",x"48",x"c1"),
   421 => (x"c3",x"7c",x"75",x"87"),
   422 => (x"49",x"76",x"7c",x"fe"),
   423 => (x"66",x"dc",x"79",x"c0"),
   424 => (x"4b",x"72",x"4a",x"bf"),
   425 => (x"73",x"2b",x"b7",x"d8"),
   426 => (x"70",x"98",x"75",x"48"),
   427 => (x"d0",x"4b",x"72",x"7c"),
   428 => (x"48",x"73",x"2b",x"b7"),
   429 => (x"7c",x"70",x"98",x"75"),
   430 => (x"b7",x"c8",x"4b",x"72"),
   431 => (x"75",x"48",x"73",x"2b"),
   432 => (x"72",x"7c",x"70",x"98"),
   433 => (x"70",x"98",x"75",x"48"),
   434 => (x"48",x"66",x"dc",x"7c"),
   435 => (x"e0",x"c0",x"80",x"c4"),
   436 => (x"48",x"6e",x"58",x"a6"),
   437 => (x"a6",x"c4",x"80",x"c1"),
   438 => (x"c2",x"49",x"6e",x"58"),
   439 => (x"04",x"a9",x"b7",x"c0"),
   440 => (x"75",x"87",x"fb",x"fe"),
   441 => (x"75",x"7c",x"75",x"7c"),
   442 => (x"e0",x"da",x"d8",x"7c"),
   443 => (x"6c",x"7c",x"75",x"4b"),
   444 => (x"72",x"9a",x"75",x"4a"),
   445 => (x"c8",x"c0",x"05",x"9a"),
   446 => (x"73",x"8b",x"c1",x"87"),
   447 => (x"ec",x"ff",x"05",x"9b"),
   448 => (x"ff",x"7c",x"75",x"87"),
   449 => (x"c8",x"48",x"bf",x"d0"),
   450 => (x"c4",x"98",x"c0",x"c0"),
   451 => (x"02",x"6e",x"58",x"a6"),
   452 => (x"c8",x"87",x"d2",x"c0"),
   453 => (x"ff",x"4a",x"c0",x"c0"),
   454 => (x"72",x"48",x"bf",x"d0"),
   455 => (x"58",x"a6",x"c4",x"98"),
   456 => (x"f2",x"ff",x"05",x"6e"),
   457 => (x"49",x"d0",x"ff",x"87"),
   458 => (x"48",x"c0",x"79",x"c0"),
   459 => (x"26",x"4d",x"26",x"26"),
   460 => (x"26",x"4b",x"26",x"4c"),
   461 => (x"57",x"4f",x"26",x"4a"),
   462 => (x"65",x"74",x"69",x"72"),
   463 => (x"69",x"61",x"66",x"20"),
   464 => (x"0a",x"64",x"65",x"6c"),
   465 => (x"5a",x"5e",x"0e",x"00"),
   466 => (x"0e",x"5d",x"5c",x"5b"),
   467 => (x"4c",x"66",x"d8",x"1e"),
   468 => (x"76",x"4b",x"66",x"dc"),
   469 => (x"c5",x"79",x"c0",x"49"),
   470 => (x"4d",x"df",x"cd",x"ee"),
   471 => (x"c3",x"49",x"d4",x"ff"),
   472 => (x"d4",x"ff",x"79",x"ff"),
   473 => (x"ff",x"c3",x"4a",x"bf"),
   474 => (x"b7",x"fe",x"c3",x"9a"),
   475 => (x"e5",x"c1",x"05",x"aa"),
   476 => (x"19",x"a8",x"27",x"87"),
   477 => (x"c0",x"49",x"00",x"00"),
   478 => (x"ab",x"b7",x"c4",x"79"),
   479 => (x"87",x"e4",x"c0",x"04"),
   480 => (x"00",x"02",x"20",x"27"),
   481 => (x"4a",x"70",x"0f",x"00"),
   482 => (x"84",x"c4",x"7c",x"72"),
   483 => (x"00",x"19",x"a8",x"27"),
   484 => (x"72",x"48",x"bf",x"00"),
   485 => (x"19",x"ac",x"27",x"80"),
   486 => (x"c4",x"58",x"00",x"00"),
   487 => (x"ab",x"b7",x"c4",x"8b"),
   488 => (x"87",x"dc",x"ff",x"03"),
   489 => (x"06",x"ab",x"b7",x"c0"),
   490 => (x"ff",x"87",x"e5",x"c0"),
   491 => (x"ff",x"c3",x"4d",x"d4"),
   492 => (x"72",x"4a",x"6d",x"7d"),
   493 => (x"84",x"c1",x"7c",x"97"),
   494 => (x"00",x"19",x"a8",x"27"),
   495 => (x"72",x"48",x"bf",x"00"),
   496 => (x"19",x"ac",x"27",x"80"),
   497 => (x"c1",x"58",x"00",x"00"),
   498 => (x"ab",x"b7",x"c0",x"8b"),
   499 => (x"87",x"de",x"ff",x"01"),
   500 => (x"49",x"76",x"4d",x"c1"),
   501 => (x"8d",x"c1",x"79",x"c1"),
   502 => (x"fd",x"05",x"9d",x"75"),
   503 => (x"d4",x"ff",x"87",x"fe"),
   504 => (x"79",x"ff",x"c3",x"49"),
   505 => (x"26",x"26",x"48",x"6e"),
   506 => (x"26",x"4c",x"26",x"4d"),
   507 => (x"26",x"4a",x"26",x"4b"),
   508 => (x"5a",x"5e",x"0e",x"4f"),
   509 => (x"0e",x"5d",x"5c",x"5b"),
   510 => (x"4b",x"d0",x"ff",x"1e"),
   511 => (x"4a",x"c0",x"c0",x"c8"),
   512 => (x"d4",x"ff",x"4c",x"c0"),
   513 => (x"79",x"ff",x"c3",x"49"),
   514 => (x"98",x"72",x"48",x"6b"),
   515 => (x"6e",x"58",x"a6",x"c4"),
   516 => (x"87",x"cc",x"c0",x"02"),
   517 => (x"98",x"72",x"48",x"6b"),
   518 => (x"6e",x"58",x"a6",x"c4"),
   519 => (x"87",x"f4",x"ff",x"05"),
   520 => (x"ff",x"7b",x"c1",x"c4"),
   521 => (x"ff",x"c3",x"49",x"d4"),
   522 => (x"1e",x"66",x"d8",x"79"),
   523 => (x"c1",x"f0",x"ff",x"c0"),
   524 => (x"66",x"27",x"1e",x"d1"),
   525 => (x"0f",x"00",x"00",x"02"),
   526 => (x"4d",x"70",x"86",x"c8"),
   527 => (x"c0",x"02",x"9d",x"75"),
   528 => (x"1e",x"75",x"87",x"d6"),
   529 => (x"27",x"1e",x"66",x"dc"),
   530 => (x"00",x"00",x"08",x"8d"),
   531 => (x"00",x"94",x"27",x"1e"),
   532 => (x"cc",x"0f",x"00",x"00"),
   533 => (x"87",x"e8",x"c0",x"86"),
   534 => (x"c0",x"1e",x"c0",x"c8"),
   535 => (x"fb",x"1e",x"66",x"e0"),
   536 => (x"86",x"c8",x"87",x"e3"),
   537 => (x"48",x"6b",x"4c",x"70"),
   538 => (x"a6",x"c4",x"98",x"72"),
   539 => (x"c0",x"02",x"6e",x"58"),
   540 => (x"48",x"6b",x"87",x"cc"),
   541 => (x"a6",x"c4",x"98",x"72"),
   542 => (x"ff",x"05",x"6e",x"58"),
   543 => (x"7b",x"c0",x"87",x"f4"),
   544 => (x"26",x"26",x"48",x"74"),
   545 => (x"26",x"4c",x"26",x"4d"),
   546 => (x"26",x"4a",x"26",x"4b"),
   547 => (x"61",x"65",x"52",x"4f"),
   548 => (x"6f",x"63",x"20",x"64"),
   549 => (x"6e",x"61",x"6d",x"6d"),
   550 => (x"61",x"66",x"20",x"64"),
   551 => (x"64",x"65",x"6c",x"69"),
   552 => (x"20",x"74",x"61",x"20"),
   553 => (x"28",x"20",x"64",x"25"),
   554 => (x"0a",x"29",x"64",x"25"),
   555 => (x"5a",x"5e",x"0e",x"00"),
   556 => (x"0e",x"5d",x"5c",x"5b"),
   557 => (x"c0",x"1e",x"c0",x"1e"),
   558 => (x"c9",x"c1",x"f0",x"ff"),
   559 => (x"02",x"66",x"27",x"1e"),
   560 => (x"c8",x"0f",x"00",x"00"),
   561 => (x"27",x"1e",x"d2",x"86"),
   562 => (x"00",x"00",x"19",x"b8"),
   563 => (x"87",x"f5",x"f9",x"1e"),
   564 => (x"4d",x"c0",x"86",x"c8"),
   565 => (x"b7",x"d2",x"85",x"c1"),
   566 => (x"f7",x"ff",x"04",x"ad"),
   567 => (x"19",x"b8",x"27",x"87"),
   568 => (x"bf",x"97",x"00",x"00"),
   569 => (x"9a",x"c0",x"c3",x"4a"),
   570 => (x"aa",x"b7",x"c0",x"c1"),
   571 => (x"87",x"f2",x"c0",x"05"),
   572 => (x"00",x"19",x"bf",x"27"),
   573 => (x"4a",x"bf",x"97",x"00"),
   574 => (x"c0",x"27",x"32",x"d0"),
   575 => (x"97",x"00",x"00",x"19"),
   576 => (x"33",x"c8",x"4b",x"bf"),
   577 => (x"b2",x"73",x"4a",x"72"),
   578 => (x"00",x"19",x"c1",x"27"),
   579 => (x"4b",x"bf",x"97",x"00"),
   580 => (x"b2",x"73",x"4a",x"72"),
   581 => (x"ff",x"ff",x"ff",x"cf"),
   582 => (x"c1",x"4d",x"72",x"9a"),
   583 => (x"c3",x"35",x"ca",x"85"),
   584 => (x"c1",x"27",x"87",x"cb"),
   585 => (x"97",x"00",x"00",x"19"),
   586 => (x"32",x"c1",x"4a",x"bf"),
   587 => (x"c2",x"27",x"9a",x"c6"),
   588 => (x"97",x"00",x"00",x"19"),
   589 => (x"b7",x"c7",x"4b",x"bf"),
   590 => (x"73",x"4a",x"72",x"2b"),
   591 => (x"19",x"bd",x"27",x"b2"),
   592 => (x"bf",x"97",x"00",x"00"),
   593 => (x"cf",x"48",x"73",x"4b"),
   594 => (x"58",x"a6",x"c4",x"98"),
   595 => (x"00",x"19",x"be",x"27"),
   596 => (x"4b",x"bf",x"97",x"00"),
   597 => (x"33",x"ca",x"9b",x"c3"),
   598 => (x"00",x"19",x"bf",x"27"),
   599 => (x"4c",x"bf",x"97",x"00"),
   600 => (x"4b",x"73",x"34",x"c2"),
   601 => (x"c0",x"27",x"b3",x"74"),
   602 => (x"97",x"00",x"00",x"19"),
   603 => (x"c0",x"c3",x"4c",x"bf"),
   604 => (x"2c",x"b7",x"c6",x"9c"),
   605 => (x"b3",x"74",x"4b",x"73"),
   606 => (x"66",x"c4",x"1e",x"73"),
   607 => (x"27",x"1e",x"72",x"1e"),
   608 => (x"00",x"00",x"09",x"fa"),
   609 => (x"00",x"94",x"27",x"1e"),
   610 => (x"d0",x"0f",x"00",x"00"),
   611 => (x"c1",x"82",x"c2",x"86"),
   612 => (x"70",x"30",x"72",x"48"),
   613 => (x"27",x"1e",x"72",x"4a"),
   614 => (x"00",x"00",x"0a",x"27"),
   615 => (x"00",x"94",x"27",x"1e"),
   616 => (x"c8",x"0f",x"00",x"00"),
   617 => (x"6e",x"48",x"c1",x"86"),
   618 => (x"58",x"a6",x"c4",x"30"),
   619 => (x"4d",x"73",x"83",x"c1"),
   620 => (x"1e",x"6e",x"95",x"72"),
   621 => (x"30",x"27",x"1e",x"75"),
   622 => (x"1e",x"00",x"00",x"0a"),
   623 => (x"00",x"00",x"94",x"27"),
   624 => (x"86",x"cc",x"0f",x"00"),
   625 => (x"c0",x"c8",x"49",x"6e"),
   626 => (x"c0",x"06",x"a9",x"b7"),
   627 => (x"4a",x"6e",x"87",x"cf"),
   628 => (x"b7",x"c1",x"35",x"c1"),
   629 => (x"b7",x"c0",x"c8",x"2a"),
   630 => (x"f3",x"ff",x"01",x"aa"),
   631 => (x"27",x"1e",x"75",x"87"),
   632 => (x"00",x"00",x"0a",x"46"),
   633 => (x"00",x"94",x"27",x"1e"),
   634 => (x"c8",x"0f",x"00",x"00"),
   635 => (x"26",x"48",x"75",x"86"),
   636 => (x"4c",x"26",x"4d",x"26"),
   637 => (x"4a",x"26",x"4b",x"26"),
   638 => (x"5f",x"63",x"4f",x"26"),
   639 => (x"65",x"7a",x"69",x"73"),
   640 => (x"6c",x"75",x"6d",x"5f"),
   641 => (x"25",x"20",x"3a",x"74"),
   642 => (x"72",x"20",x"2c",x"64"),
   643 => (x"5f",x"64",x"61",x"65"),
   644 => (x"6c",x"5f",x"6c",x"62"),
   645 => (x"20",x"3a",x"6e",x"65"),
   646 => (x"20",x"2c",x"64",x"25"),
   647 => (x"7a",x"69",x"73",x"63"),
   648 => (x"25",x"20",x"3a",x"65"),
   649 => (x"4d",x"00",x"0a",x"64"),
   650 => (x"20",x"74",x"6c",x"75"),
   651 => (x"00",x"0a",x"64",x"25"),
   652 => (x"62",x"20",x"64",x"25"),
   653 => (x"6b",x"63",x"6f",x"6c"),
   654 => (x"66",x"6f",x"20",x"73"),
   655 => (x"7a",x"69",x"73",x"20"),
   656 => (x"64",x"25",x"20",x"65"),
   657 => (x"64",x"25",x"00",x"0a"),
   658 => (x"6f",x"6c",x"62",x"20"),
   659 => (x"20",x"73",x"6b",x"63"),
   660 => (x"35",x"20",x"66",x"6f"),
   661 => (x"62",x"20",x"32",x"31"),
   662 => (x"73",x"65",x"74",x"79"),
   663 => (x"5e",x"0e",x"00",x"0a"),
   664 => (x"5d",x"5c",x"5b",x"5a"),
   665 => (x"4d",x"66",x"d4",x"0e"),
   666 => (x"66",x"dc",x"4c",x"c0"),
   667 => (x"a9",x"b7",x"c0",x"49"),
   668 => (x"87",x"fb",x"c0",x"06"),
   669 => (x"c0",x"c1",x"4b",x"15"),
   670 => (x"93",x"c0",x"c0",x"c0"),
   671 => (x"93",x"b7",x"c0",x"c4"),
   672 => (x"97",x"66",x"d8",x"4b"),
   673 => (x"c0",x"c1",x"4a",x"bf"),
   674 => (x"92",x"c0",x"c0",x"c0"),
   675 => (x"92",x"b7",x"c0",x"c4"),
   676 => (x"48",x"66",x"d8",x"4a"),
   677 => (x"a6",x"dc",x"80",x"c1"),
   678 => (x"ab",x"b7",x"72",x"58"),
   679 => (x"87",x"c5",x"c0",x"02"),
   680 => (x"cc",x"c0",x"48",x"c1"),
   681 => (x"dc",x"84",x"c1",x"87"),
   682 => (x"04",x"ac",x"b7",x"66"),
   683 => (x"c0",x"87",x"c5",x"ff"),
   684 => (x"26",x"4d",x"26",x"48"),
   685 => (x"26",x"4b",x"26",x"4c"),
   686 => (x"0e",x"4f",x"26",x"4a"),
   687 => (x"5c",x"5b",x"5a",x"5e"),
   688 => (x"e0",x"27",x"0e",x"5d"),
   689 => (x"49",x"00",x"00",x"1b"),
   690 => (x"ee",x"27",x"79",x"c0"),
   691 => (x"1e",x"00",x"00",x"18"),
   692 => (x"00",x"00",x"5e",x"27"),
   693 => (x"86",x"c4",x"0f",x"00"),
   694 => (x"00",x"19",x"d8",x"27"),
   695 => (x"1e",x"c0",x"1e",x"00"),
   696 => (x"00",x"07",x"f1",x"27"),
   697 => (x"86",x"c8",x"0f",x"00"),
   698 => (x"9a",x"72",x"4a",x"70"),
   699 => (x"87",x"d3",x"c0",x"05"),
   700 => (x"00",x"18",x"1a",x"27"),
   701 => (x"5e",x"27",x"1e",x"00"),
   702 => (x"0f",x"00",x"00",x"00"),
   703 => (x"48",x"c0",x"86",x"c4"),
   704 => (x"27",x"87",x"d8",x"cf"),
   705 => (x"00",x"00",x"18",x"fb"),
   706 => (x"00",x"5e",x"27",x"1e"),
   707 => (x"c4",x"0f",x"00",x"00"),
   708 => (x"27",x"4c",x"c0",x"86"),
   709 => (x"00",x"00",x"1c",x"0c"),
   710 => (x"c8",x"79",x"c1",x"49"),
   711 => (x"19",x"12",x"27",x"1e"),
   712 => (x"27",x"1e",x"00",x"00"),
   713 => (x"00",x"00",x"1a",x"0e"),
   714 => (x"0a",x"5e",x"27",x"1e"),
   715 => (x"cc",x"0f",x"00",x"00"),
   716 => (x"72",x"4a",x"70",x"86"),
   717 => (x"c8",x"c0",x"05",x"9a"),
   718 => (x"1c",x"0c",x"27",x"87"),
   719 => (x"c0",x"49",x"00",x"00"),
   720 => (x"27",x"1e",x"c8",x"79"),
   721 => (x"00",x"00",x"19",x"1b"),
   722 => (x"1a",x"2a",x"27",x"1e"),
   723 => (x"27",x"1e",x"00",x"00"),
   724 => (x"00",x"00",x"0a",x"5e"),
   725 => (x"70",x"86",x"cc",x"0f"),
   726 => (x"05",x"9a",x"72",x"4a"),
   727 => (x"27",x"87",x"c8",x"c0"),
   728 => (x"00",x"00",x"1c",x"0c"),
   729 => (x"27",x"79",x"c0",x"49"),
   730 => (x"00",x"00",x"1c",x"0c"),
   731 => (x"24",x"27",x"1e",x"bf"),
   732 => (x"1e",x"00",x"00",x"19"),
   733 => (x"00",x"00",x"94",x"27"),
   734 => (x"86",x"c8",x"0f",x"00"),
   735 => (x"00",x"1c",x"0c",x"27"),
   736 => (x"c3",x"02",x"bf",x"00"),
   737 => (x"d8",x"27",x"87",x"c0"),
   738 => (x"4d",x"00",x"00",x"19"),
   739 => (x"00",x"1b",x"96",x"27"),
   740 => (x"d6",x"27",x"4b",x"00"),
   741 => (x"9f",x"00",x"00",x"1b"),
   742 => (x"1e",x"72",x"4a",x"bf"),
   743 => (x"00",x"1b",x"d6",x"27"),
   744 => (x"d8",x"27",x"4a",x"00"),
   745 => (x"8a",x"00",x"00",x"19"),
   746 => (x"1e",x"d0",x"1e",x"72"),
   747 => (x"27",x"1e",x"c0",x"c8"),
   748 => (x"00",x"00",x"18",x"4c"),
   749 => (x"00",x"94",x"27",x"1e"),
   750 => (x"d4",x"0f",x"00",x"00"),
   751 => (x"c8",x"4a",x"73",x"86"),
   752 => (x"27",x"4c",x"6a",x"82"),
   753 => (x"00",x"00",x"1b",x"d6"),
   754 => (x"c5",x"4a",x"bf",x"9f"),
   755 => (x"aa",x"b7",x"ea",x"d6"),
   756 => (x"87",x"d3",x"c0",x"05"),
   757 => (x"82",x"c8",x"4a",x"73"),
   758 => (x"46",x"27",x"1e",x"6a"),
   759 => (x"0f",x"00",x"00",x"12"),
   760 => (x"4c",x"70",x"86",x"c4"),
   761 => (x"75",x"87",x"e4",x"c0"),
   762 => (x"82",x"fe",x"c7",x"4a"),
   763 => (x"ca",x"4a",x"6a",x"9f"),
   764 => (x"aa",x"b7",x"d5",x"e9"),
   765 => (x"87",x"d3",x"c0",x"02"),
   766 => (x"00",x"18",x"2e",x"27"),
   767 => (x"5e",x"27",x"1e",x"00"),
   768 => (x"0f",x"00",x"00",x"00"),
   769 => (x"48",x"c0",x"86",x"c4"),
   770 => (x"74",x"87",x"d0",x"cb"),
   771 => (x"18",x"89",x"27",x"1e"),
   772 => (x"27",x"1e",x"00",x"00"),
   773 => (x"00",x"00",x"00",x"94"),
   774 => (x"27",x"86",x"c8",x"0f"),
   775 => (x"00",x"00",x"19",x"d8"),
   776 => (x"27",x"1e",x"74",x"1e"),
   777 => (x"00",x"00",x"07",x"f1"),
   778 => (x"70",x"86",x"c8",x"0f"),
   779 => (x"05",x"9a",x"72",x"4a"),
   780 => (x"c0",x"87",x"c5",x"c0"),
   781 => (x"87",x"e3",x"ca",x"48"),
   782 => (x"00",x"18",x"a1",x"27"),
   783 => (x"5e",x"27",x"1e",x"00"),
   784 => (x"0f",x"00",x"00",x"00"),
   785 => (x"37",x"27",x"86",x"c4"),
   786 => (x"1e",x"00",x"00",x"19"),
   787 => (x"00",x"00",x"94",x"27"),
   788 => (x"86",x"c4",x"0f",x"00"),
   789 => (x"4f",x"27",x"1e",x"c8"),
   790 => (x"1e",x"00",x"00",x"19"),
   791 => (x"00",x"1a",x"2a",x"27"),
   792 => (x"5e",x"27",x"1e",x"00"),
   793 => (x"0f",x"00",x"00",x"0a"),
   794 => (x"4a",x"70",x"86",x"cc"),
   795 => (x"c0",x"05",x"9a",x"72"),
   796 => (x"e0",x"27",x"87",x"cb"),
   797 => (x"49",x"00",x"00",x"1b"),
   798 => (x"f1",x"c0",x"79",x"c1"),
   799 => (x"27",x"1e",x"c8",x"87"),
   800 => (x"00",x"00",x"19",x"58"),
   801 => (x"1a",x"0e",x"27",x"1e"),
   802 => (x"27",x"1e",x"00",x"00"),
   803 => (x"00",x"00",x"0a",x"5e"),
   804 => (x"70",x"86",x"cc",x"0f"),
   805 => (x"02",x"9a",x"72",x"4a"),
   806 => (x"27",x"87",x"d3",x"c0"),
   807 => (x"00",x"00",x"18",x"c8"),
   808 => (x"00",x"94",x"27",x"1e"),
   809 => (x"c4",x"0f",x"00",x"00"),
   810 => (x"c8",x"48",x"c0",x"86"),
   811 => (x"d6",x"27",x"87",x"ed"),
   812 => (x"97",x"00",x"00",x"1b"),
   813 => (x"d5",x"c1",x"4a",x"bf"),
   814 => (x"c0",x"05",x"aa",x"b7"),
   815 => (x"d7",x"27",x"87",x"d0"),
   816 => (x"97",x"00",x"00",x"1b"),
   817 => (x"ea",x"c2",x"4a",x"bf"),
   818 => (x"c0",x"02",x"aa",x"b7"),
   819 => (x"48",x"c0",x"87",x"c5"),
   820 => (x"27",x"87",x"c8",x"c8"),
   821 => (x"00",x"00",x"19",x"d8"),
   822 => (x"c3",x"4a",x"bf",x"97"),
   823 => (x"02",x"aa",x"b7",x"e9"),
   824 => (x"27",x"87",x"d5",x"c0"),
   825 => (x"00",x"00",x"19",x"d8"),
   826 => (x"c3",x"4a",x"bf",x"97"),
   827 => (x"02",x"aa",x"b7",x"eb"),
   828 => (x"c0",x"87",x"c5",x"c0"),
   829 => (x"87",x"e3",x"c7",x"48"),
   830 => (x"00",x"19",x"e3",x"27"),
   831 => (x"4a",x"bf",x"97",x"00"),
   832 => (x"c0",x"05",x"9a",x"72"),
   833 => (x"e4",x"27",x"87",x"cf"),
   834 => (x"97",x"00",x"00",x"19"),
   835 => (x"b7",x"c2",x"4a",x"bf"),
   836 => (x"c5",x"c0",x"02",x"aa"),
   837 => (x"c7",x"48",x"c0",x"87"),
   838 => (x"e5",x"27",x"87",x"c1"),
   839 => (x"97",x"00",x"00",x"19"),
   840 => (x"dc",x"27",x"48",x"bf"),
   841 => (x"58",x"00",x"00",x"1b"),
   842 => (x"00",x"1b",x"d8",x"27"),
   843 => (x"72",x"4a",x"bf",x"00"),
   844 => (x"27",x"8b",x"c1",x"4b"),
   845 => (x"00",x"00",x"1b",x"dc"),
   846 => (x"73",x"79",x"73",x"49"),
   847 => (x"27",x"1e",x"72",x"1e"),
   848 => (x"00",x"00",x"19",x"61"),
   849 => (x"00",x"94",x"27",x"1e"),
   850 => (x"cc",x"0f",x"00",x"00"),
   851 => (x"19",x"e6",x"27",x"86"),
   852 => (x"bf",x"97",x"00",x"00"),
   853 => (x"27",x"82",x"74",x"4a"),
   854 => (x"00",x"00",x"19",x"e7"),
   855 => (x"c8",x"4b",x"bf",x"97"),
   856 => (x"72",x"48",x"73",x"33"),
   857 => (x"1b",x"f0",x"27",x"80"),
   858 => (x"27",x"58",x"00",x"00"),
   859 => (x"00",x"00",x"19",x"e8"),
   860 => (x"27",x"48",x"bf",x"97"),
   861 => (x"00",x"00",x"1c",x"04"),
   862 => (x"1b",x"e0",x"27",x"58"),
   863 => (x"02",x"bf",x"00",x"00"),
   864 => (x"c8",x"87",x"df",x"c3"),
   865 => (x"18",x"e5",x"27",x"1e"),
   866 => (x"27",x"1e",x"00",x"00"),
   867 => (x"00",x"00",x"1a",x"2a"),
   868 => (x"0a",x"5e",x"27",x"1e"),
   869 => (x"cc",x"0f",x"00",x"00"),
   870 => (x"72",x"4a",x"70",x"86"),
   871 => (x"c5",x"c0",x"02",x"9a"),
   872 => (x"c4",x"48",x"c0",x"87"),
   873 => (x"d8",x"27",x"87",x"f5"),
   874 => (x"bf",x"00",x"00",x"1b"),
   875 => (x"c4",x"48",x"73",x"4b"),
   876 => (x"1c",x"08",x"27",x"30"),
   877 => (x"27",x"58",x"00",x"00"),
   878 => (x"00",x"00",x"1b",x"fc"),
   879 => (x"27",x"79",x"73",x"49"),
   880 => (x"00",x"00",x"19",x"fd"),
   881 => (x"c8",x"4a",x"bf",x"97"),
   882 => (x"19",x"fc",x"27",x"32"),
   883 => (x"bf",x"97",x"00",x"00"),
   884 => (x"74",x"4a",x"72",x"4c"),
   885 => (x"19",x"fe",x"27",x"82"),
   886 => (x"bf",x"97",x"00",x"00"),
   887 => (x"72",x"34",x"d0",x"4c"),
   888 => (x"27",x"82",x"74",x"4a"),
   889 => (x"00",x"00",x"19",x"ff"),
   890 => (x"d8",x"4c",x"bf",x"97"),
   891 => (x"74",x"4a",x"72",x"34"),
   892 => (x"1c",x"08",x"27",x"82"),
   893 => (x"72",x"49",x"00",x"00"),
   894 => (x"27",x"4a",x"72",x"79"),
   895 => (x"00",x"00",x"1c",x"00"),
   896 => (x"4a",x"72",x"92",x"bf"),
   897 => (x"00",x"1b",x"ec",x"27"),
   898 => (x"27",x"82",x"bf",x"00"),
   899 => (x"00",x"00",x"1b",x"f0"),
   900 => (x"27",x"79",x"72",x"49"),
   901 => (x"00",x"00",x"1a",x"05"),
   902 => (x"c8",x"4c",x"bf",x"97"),
   903 => (x"1a",x"04",x"27",x"34"),
   904 => (x"bf",x"97",x"00",x"00"),
   905 => (x"75",x"4c",x"74",x"4d"),
   906 => (x"1a",x"06",x"27",x"84"),
   907 => (x"bf",x"97",x"00",x"00"),
   908 => (x"74",x"35",x"d0",x"4d"),
   909 => (x"27",x"84",x"75",x"4c"),
   910 => (x"00",x"00",x"1a",x"07"),
   911 => (x"cf",x"4d",x"bf",x"97"),
   912 => (x"74",x"35",x"d8",x"9d"),
   913 => (x"27",x"84",x"75",x"4c"),
   914 => (x"00",x"00",x"1b",x"f4"),
   915 => (x"c2",x"79",x"74",x"49"),
   916 => (x"74",x"4b",x"73",x"8c"),
   917 => (x"72",x"48",x"73",x"93"),
   918 => (x"1b",x"fc",x"27",x"80"),
   919 => (x"c1",x"58",x"00",x"00"),
   920 => (x"ea",x"27",x"87",x"f7"),
   921 => (x"97",x"00",x"00",x"19"),
   922 => (x"32",x"c8",x"4a",x"bf"),
   923 => (x"00",x"19",x"e9",x"27"),
   924 => (x"4b",x"bf",x"97",x"00"),
   925 => (x"82",x"73",x"4a",x"72"),
   926 => (x"00",x"1c",x"04",x"27"),
   927 => (x"79",x"72",x"49",x"00"),
   928 => (x"ff",x"c7",x"32",x"c5"),
   929 => (x"27",x"2a",x"c9",x"82"),
   930 => (x"00",x"00",x"1b",x"fc"),
   931 => (x"27",x"79",x"72",x"49"),
   932 => (x"00",x"00",x"19",x"ef"),
   933 => (x"c8",x"4b",x"bf",x"97"),
   934 => (x"19",x"ee",x"27",x"33"),
   935 => (x"bf",x"97",x"00",x"00"),
   936 => (x"74",x"4b",x"73",x"4c"),
   937 => (x"1c",x"08",x"27",x"83"),
   938 => (x"73",x"49",x"00",x"00"),
   939 => (x"27",x"4b",x"73",x"79"),
   940 => (x"00",x"00",x"1c",x"00"),
   941 => (x"4b",x"73",x"93",x"bf"),
   942 => (x"00",x"1b",x"ec",x"27"),
   943 => (x"27",x"83",x"bf",x"00"),
   944 => (x"00",x"00",x"1b",x"f8"),
   945 => (x"27",x"79",x"73",x"49"),
   946 => (x"00",x"00",x"1b",x"f4"),
   947 => (x"73",x"79",x"c0",x"49"),
   948 => (x"27",x"80",x"72",x"48"),
   949 => (x"00",x"00",x"1b",x"f4"),
   950 => (x"26",x"48",x"c1",x"58"),
   951 => (x"26",x"4c",x"26",x"4d"),
   952 => (x"26",x"4a",x"26",x"4b"),
   953 => (x"5a",x"5e",x"0e",x"4f"),
   954 => (x"0e",x"5d",x"5c",x"5b"),
   955 => (x"00",x"1b",x"e0",x"27"),
   956 => (x"c0",x"02",x"bf",x"00"),
   957 => (x"66",x"d4",x"87",x"cf"),
   958 => (x"2c",x"b7",x"c7",x"4c"),
   959 => (x"c1",x"4b",x"66",x"d4"),
   960 => (x"cc",x"c0",x"9b",x"ff"),
   961 => (x"4c",x"66",x"d4",x"87"),
   962 => (x"d4",x"2c",x"b7",x"c8"),
   963 => (x"ff",x"c3",x"4b",x"66"),
   964 => (x"19",x"d8",x"27",x"9b"),
   965 => (x"27",x"1e",x"00",x"00"),
   966 => (x"00",x"00",x"1b",x"ec"),
   967 => (x"82",x"74",x"4a",x"bf"),
   968 => (x"f1",x"27",x"1e",x"72"),
   969 => (x"0f",x"00",x"00",x"07"),
   970 => (x"4a",x"70",x"86",x"c8"),
   971 => (x"c0",x"05",x"9a",x"72"),
   972 => (x"48",x"c0",x"87",x"c5"),
   973 => (x"27",x"87",x"f2",x"c0"),
   974 => (x"00",x"00",x"1b",x"e0"),
   975 => (x"d7",x"c0",x"02",x"bf"),
   976 => (x"c4",x"4a",x"73",x"87"),
   977 => (x"27",x"4a",x"72",x"92"),
   978 => (x"00",x"00",x"19",x"d8"),
   979 => (x"cf",x"4d",x"6a",x"82"),
   980 => (x"ff",x"ff",x"ff",x"ff"),
   981 => (x"87",x"cf",x"c0",x"9d"),
   982 => (x"92",x"c2",x"4a",x"73"),
   983 => (x"d8",x"27",x"4a",x"72"),
   984 => (x"82",x"00",x"00",x"19"),
   985 => (x"75",x"4d",x"6a",x"9f"),
   986 => (x"26",x"4d",x"26",x"48"),
   987 => (x"26",x"4b",x"26",x"4c"),
   988 => (x"0e",x"4f",x"26",x"4a"),
   989 => (x"5c",x"5b",x"5a",x"5e"),
   990 => (x"8e",x"cc",x"0e",x"5d"),
   991 => (x"ff",x"ff",x"ff",x"cf"),
   992 => (x"4c",x"c0",x"4d",x"f8"),
   993 => (x"f4",x"27",x"49",x"76"),
   994 => (x"bf",x"00",x"00",x"1b"),
   995 => (x"49",x"a6",x"c4",x"79"),
   996 => (x"00",x"1b",x"f8",x"27"),
   997 => (x"27",x"79",x"bf",x"00"),
   998 => (x"00",x"00",x"1b",x"e0"),
   999 => (x"cc",x"c0",x"02",x"bf"),
  1000 => (x"1b",x"d8",x"27",x"87"),
  1001 => (x"4a",x"bf",x"00",x"00"),
  1002 => (x"c9",x"c0",x"32",x"c4"),
  1003 => (x"1b",x"fc",x"27",x"87"),
  1004 => (x"4a",x"bf",x"00",x"00"),
  1005 => (x"a6",x"c8",x"32",x"c4"),
  1006 => (x"c0",x"79",x"72",x"49"),
  1007 => (x"49",x"66",x"c8",x"4b"),
  1008 => (x"c3",x"06",x"a9",x"c0"),
  1009 => (x"4a",x"73",x"87",x"d0"),
  1010 => (x"9a",x"72",x"9a",x"cf"),
  1011 => (x"87",x"e4",x"c0",x"05"),
  1012 => (x"00",x"19",x"d8",x"27"),
  1013 => (x"66",x"c8",x"1e",x"00"),
  1014 => (x"48",x"66",x"c8",x"4a"),
  1015 => (x"a6",x"cc",x"80",x"c1"),
  1016 => (x"27",x"1e",x"72",x"58"),
  1017 => (x"00",x"00",x"07",x"f1"),
  1018 => (x"27",x"86",x"c8",x"0f"),
  1019 => (x"00",x"00",x"19",x"d8"),
  1020 => (x"87",x"c3",x"c0",x"4c"),
  1021 => (x"97",x"84",x"e0",x"c0"),
  1022 => (x"9a",x"72",x"4a",x"6c"),
  1023 => (x"87",x"cd",x"c2",x"02"),
  1024 => (x"c3",x"4a",x"6c",x"97"),
  1025 => (x"02",x"aa",x"b7",x"e5"),
  1026 => (x"74",x"87",x"c2",x"c2"),
  1027 => (x"97",x"82",x"cb",x"4a"),
  1028 => (x"9a",x"d8",x"4a",x"6a"),
  1029 => (x"c1",x"05",x"9a",x"72"),
  1030 => (x"1e",x"74",x"87",x"f3"),
  1031 => (x"00",x"00",x"5e",x"27"),
  1032 => (x"86",x"c4",x"0f",x"00"),
  1033 => (x"e8",x"c0",x"1e",x"cb"),
  1034 => (x"1e",x"74",x"1e",x"66"),
  1035 => (x"00",x"0a",x"5e",x"27"),
  1036 => (x"86",x"cc",x"0f",x"00"),
  1037 => (x"9a",x"72",x"4a",x"70"),
  1038 => (x"87",x"d1",x"c1",x"05"),
  1039 => (x"83",x"dc",x"4b",x"74"),
  1040 => (x"4a",x"66",x"e0",x"c0"),
  1041 => (x"7a",x"6b",x"82",x"c4"),
  1042 => (x"83",x"da",x"4b",x"74"),
  1043 => (x"4a",x"66",x"e0",x"c0"),
  1044 => (x"6b",x"9f",x"82",x"c8"),
  1045 => (x"72",x"7a",x"70",x"48"),
  1046 => (x"1b",x"e0",x"27",x"4d"),
  1047 => (x"02",x"bf",x"00",x"00"),
  1048 => (x"74",x"87",x"d5",x"c0"),
  1049 => (x"9f",x"82",x"d4",x"4a"),
  1050 => (x"ff",x"c0",x"4a",x"6a"),
  1051 => (x"48",x"72",x"9a",x"ff"),
  1052 => (x"a6",x"c4",x"30",x"d0"),
  1053 => (x"87",x"c4",x"c0",x"58"),
  1054 => (x"79",x"c0",x"49",x"76"),
  1055 => (x"80",x"6d",x"48",x"6e"),
  1056 => (x"e0",x"c0",x"7d",x"70"),
  1057 => (x"79",x"c0",x"49",x"66"),
  1058 => (x"ce",x"c1",x"48",x"c1"),
  1059 => (x"c8",x"83",x"c1",x"87"),
  1060 => (x"fc",x"04",x"ab",x"66"),
  1061 => (x"ff",x"cf",x"87",x"f0"),
  1062 => (x"4d",x"f8",x"ff",x"ff"),
  1063 => (x"00",x"1b",x"e0",x"27"),
  1064 => (x"c0",x"02",x"bf",x"00"),
  1065 => (x"1e",x"6e",x"87",x"f3"),
  1066 => (x"00",x"0e",x"e5",x"27"),
  1067 => (x"86",x"c4",x"0f",x"00"),
  1068 => (x"6e",x"58",x"a6",x"c4"),
  1069 => (x"75",x"9a",x"75",x"4a"),
  1070 => (x"dc",x"c0",x"02",x"aa"),
  1071 => (x"c2",x"4a",x"6e",x"87"),
  1072 => (x"27",x"4a",x"72",x"8a"),
  1073 => (x"00",x"00",x"1b",x"d8"),
  1074 => (x"f0",x"27",x"92",x"bf"),
  1075 => (x"bf",x"00",x"00",x"1b"),
  1076 => (x"c8",x"80",x"72",x"48"),
  1077 => (x"e2",x"fb",x"58",x"a6"),
  1078 => (x"cf",x"48",x"c0",x"87"),
  1079 => (x"f8",x"ff",x"ff",x"ff"),
  1080 => (x"26",x"86",x"cc",x"4d"),
  1081 => (x"26",x"4c",x"26",x"4d"),
  1082 => (x"26",x"4a",x"26",x"4b"),
  1083 => (x"5a",x"5e",x"0e",x"4f"),
  1084 => (x"66",x"cc",x"0e",x"5b"),
  1085 => (x"82",x"c1",x"4a",x"bf"),
  1086 => (x"72",x"49",x"66",x"cc"),
  1087 => (x"27",x"4a",x"72",x"79"),
  1088 => (x"00",x"00",x"1b",x"dc"),
  1089 => (x"9a",x"72",x"9a",x"bf"),
  1090 => (x"87",x"d3",x"c0",x"05"),
  1091 => (x"c8",x"4a",x"66",x"cc"),
  1092 => (x"27",x"1e",x"6a",x"82"),
  1093 => (x"00",x"00",x"0e",x"e5"),
  1094 => (x"70",x"86",x"c4",x"0f"),
  1095 => (x"c1",x"7a",x"73",x"4b"),
  1096 => (x"26",x"4b",x"26",x"48"),
  1097 => (x"0e",x"4f",x"26",x"4a"),
  1098 => (x"0e",x"5b",x"5a",x"5e"),
  1099 => (x"00",x"1b",x"f0",x"27"),
  1100 => (x"cc",x"4a",x"bf",x"00"),
  1101 => (x"83",x"c8",x"4b",x"66"),
  1102 => (x"8b",x"c2",x"4b",x"6b"),
  1103 => (x"d8",x"27",x"4b",x"73"),
  1104 => (x"bf",x"00",x"00",x"1b"),
  1105 => (x"73",x"4a",x"72",x"93"),
  1106 => (x"1b",x"dc",x"27",x"82"),
  1107 => (x"4b",x"bf",x"00",x"00"),
  1108 => (x"9b",x"bf",x"66",x"cc"),
  1109 => (x"82",x"73",x"4a",x"72"),
  1110 => (x"72",x"1e",x"66",x"d0"),
  1111 => (x"07",x"f1",x"27",x"1e"),
  1112 => (x"c8",x"0f",x"00",x"00"),
  1113 => (x"72",x"4a",x"70",x"86"),
  1114 => (x"c5",x"c0",x"05",x"9a"),
  1115 => (x"c0",x"48",x"c0",x"87"),
  1116 => (x"48",x"c1",x"87",x"c2"),
  1117 => (x"4a",x"26",x"4b",x"26"),
  1118 => (x"5e",x"0e",x"4f",x"26"),
  1119 => (x"5d",x"5c",x"5b",x"5a"),
  1120 => (x"4c",x"66",x"d8",x"0e"),
  1121 => (x"27",x"1e",x"66",x"d4"),
  1122 => (x"00",x"00",x"1c",x"10"),
  1123 => (x"0f",x"73",x"27",x"1e"),
  1124 => (x"c8",x"0f",x"00",x"00"),
  1125 => (x"72",x"4a",x"70",x"86"),
  1126 => (x"df",x"c1",x"02",x"9a"),
  1127 => (x"1c",x"14",x"27",x"87"),
  1128 => (x"4a",x"bf",x"00",x"00"),
  1129 => (x"c9",x"82",x"ff",x"c7"),
  1130 => (x"c0",x"4d",x"72",x"2a"),
  1131 => (x"12",x"1e",x"27",x"4b"),
  1132 => (x"27",x"1e",x"00",x"00"),
  1133 => (x"00",x"00",x"00",x"5e"),
  1134 => (x"c0",x"86",x"c4",x"0f"),
  1135 => (x"c1",x"06",x"ad",x"b7"),
  1136 => (x"1e",x"74",x"87",x"d0"),
  1137 => (x"00",x"1c",x"10",x"27"),
  1138 => (x"27",x"27",x"1e",x"00"),
  1139 => (x"0f",x"00",x"00",x"11"),
  1140 => (x"4a",x"70",x"86",x"c8"),
  1141 => (x"c0",x"05",x"9a",x"72"),
  1142 => (x"48",x"c0",x"87",x"c5"),
  1143 => (x"27",x"87",x"f5",x"c0"),
  1144 => (x"00",x"00",x"1c",x"10"),
  1145 => (x"10",x"ed",x"27",x"1e"),
  1146 => (x"c4",x"0f",x"00",x"00"),
  1147 => (x"84",x"c0",x"c8",x"86"),
  1148 => (x"b7",x"75",x"83",x"c1"),
  1149 => (x"c9",x"ff",x"04",x"ab"),
  1150 => (x"87",x"d6",x"c0",x"87"),
  1151 => (x"27",x"1e",x"66",x"d4"),
  1152 => (x"00",x"00",x"12",x"37"),
  1153 => (x"00",x"94",x"27",x"1e"),
  1154 => (x"c8",x"0f",x"00",x"00"),
  1155 => (x"c0",x"48",x"c0",x"86"),
  1156 => (x"48",x"c1",x"87",x"c2"),
  1157 => (x"4c",x"26",x"4d",x"26"),
  1158 => (x"4a",x"26",x"4b",x"26"),
  1159 => (x"70",x"4f",x"4f",x"26"),
  1160 => (x"64",x"65",x"6e",x"65"),
  1161 => (x"6c",x"69",x"66",x"20"),
  1162 => (x"6c",x"20",x"2c",x"65"),
  1163 => (x"69",x"64",x"61",x"6f"),
  1164 => (x"2e",x"2e",x"67",x"6e"),
  1165 => (x"43",x"00",x"0a",x"2e"),
  1166 => (x"74",x"27",x"6e",x"61"),
  1167 => (x"65",x"70",x"6f",x"20"),
  1168 => (x"73",x"25",x"20",x"6e"),
  1169 => (x"5e",x"0e",x"00",x"0a"),
  1170 => (x"cc",x"0e",x"5b",x"5a"),
  1171 => (x"2a",x"d8",x"4a",x"66"),
  1172 => (x"cc",x"9a",x"ff",x"c3"),
  1173 => (x"2b",x"c8",x"4b",x"66"),
  1174 => (x"9b",x"c0",x"fc",x"cf"),
  1175 => (x"b2",x"73",x"4a",x"72"),
  1176 => (x"c8",x"4b",x"66",x"cc"),
  1177 => (x"f0",x"ff",x"c0",x"33"),
  1178 => (x"72",x"9b",x"c0",x"c0"),
  1179 => (x"cc",x"b2",x"73",x"4a"),
  1180 => (x"33",x"d8",x"4b",x"66"),
  1181 => (x"c0",x"c0",x"c0",x"ff"),
  1182 => (x"4a",x"72",x"9b",x"c0"),
  1183 => (x"48",x"72",x"b2",x"73"),
  1184 => (x"4a",x"26",x"4b",x"26"),
  1185 => (x"5e",x"0e",x"4f",x"26"),
  1186 => (x"cc",x"0e",x"5b",x"5a"),
  1187 => (x"2b",x"c8",x"4b",x"66"),
  1188 => (x"4b",x"9b",x"ff",x"c3"),
  1189 => (x"c8",x"4a",x"66",x"cc"),
  1190 => (x"c0",x"fc",x"cf",x"32"),
  1191 => (x"73",x"4a",x"72",x"9a"),
  1192 => (x"48",x"72",x"4a",x"b2"),
  1193 => (x"4a",x"26",x"4b",x"26"),
  1194 => (x"5e",x"0e",x"4f",x"26"),
  1195 => (x"cc",x"0e",x"5b",x"5a"),
  1196 => (x"2a",x"d0",x"4a",x"66"),
  1197 => (x"9a",x"ff",x"ff",x"cf"),
  1198 => (x"4b",x"66",x"cc",x"4a"),
  1199 => (x"c0",x"f0",x"33",x"d0"),
  1200 => (x"4a",x"72",x"9b",x"c0"),
  1201 => (x"48",x"72",x"b2",x"73"),
  1202 => (x"4a",x"26",x"4b",x"26"),
  1203 => (x"72",x"1e",x"4f",x"26"),
  1204 => (x"c0",x"c0",x"d0",x"1e"),
  1205 => (x"72",x"4a",x"c0",x"c0"),
  1206 => (x"87",x"fd",x"ff",x"0f"),
  1207 => (x"4f",x"26",x"4a",x"26"),
  1208 => (x"cc",x"1e",x"72",x"1e"),
  1209 => (x"df",x"c3",x"4a",x"66"),
  1210 => (x"8a",x"f7",x"c0",x"9a"),
  1211 => (x"03",x"aa",x"b7",x"c0"),
  1212 => (x"c0",x"87",x"c3",x"c0"),
  1213 => (x"66",x"c8",x"82",x"e7"),
  1214 => (x"cc",x"30",x"c4",x"48"),
  1215 => (x"66",x"c8",x"58",x"a6"),
  1216 => (x"cc",x"b0",x"72",x"48"),
  1217 => (x"66",x"c8",x"58",x"a6"),
  1218 => (x"26",x"4a",x"26",x"48"),
  1219 => (x"5a",x"5e",x"0e",x"4f"),
  1220 => (x"0e",x"5d",x"5c",x"5b"),
  1221 => (x"c0",x"c0",x"c0",x"d0"),
  1222 => (x"20",x"27",x"4d",x"c0"),
  1223 => (x"bf",x"00",x"00",x"1c"),
  1224 => (x"27",x"80",x"c1",x"48"),
  1225 => (x"00",x"00",x"1c",x"24"),
  1226 => (x"66",x"d4",x"97",x"58"),
  1227 => (x"c0",x"c0",x"c1",x"4a"),
  1228 => (x"c4",x"92",x"c0",x"c0"),
  1229 => (x"4a",x"92",x"b7",x"c0"),
  1230 => (x"aa",x"b7",x"d3",x"c1"),
  1231 => (x"87",x"e9",x"c0",x"05"),
  1232 => (x"00",x"1c",x"20",x"27"),
  1233 => (x"79",x"c0",x"49",x"00"),
  1234 => (x"00",x"1c",x"24",x"27"),
  1235 => (x"79",x"c0",x"49",x"00"),
  1236 => (x"00",x"1c",x"2c",x"27"),
  1237 => (x"79",x"c0",x"49",x"00"),
  1238 => (x"00",x"1c",x"30",x"27"),
  1239 => (x"79",x"c0",x"49",x"00"),
  1240 => (x"c1",x"49",x"c0",x"ff"),
  1241 => (x"cb",x"ca",x"79",x"d3"),
  1242 => (x"1c",x"20",x"27",x"87"),
  1243 => (x"49",x"bf",x"00",x"00"),
  1244 => (x"05",x"a9",x"b7",x"c1"),
  1245 => (x"ff",x"87",x"db",x"c1"),
  1246 => (x"f4",x"c1",x"49",x"c0"),
  1247 => (x"66",x"d4",x"97",x"79"),
  1248 => (x"c0",x"c0",x"c1",x"4a"),
  1249 => (x"c4",x"92",x"c0",x"c0"),
  1250 => (x"4a",x"92",x"b7",x"c0"),
  1251 => (x"30",x"27",x"1e",x"72"),
  1252 => (x"bf",x"00",x"00",x"1c"),
  1253 => (x"12",x"e0",x"27",x"1e"),
  1254 => (x"c8",x"0f",x"00",x"00"),
  1255 => (x"1c",x"34",x"27",x"86"),
  1256 => (x"27",x"58",x"00",x"00"),
  1257 => (x"00",x"00",x"1c",x"30"),
  1258 => (x"b7",x"c3",x"4c",x"bf"),
  1259 => (x"c6",x"c0",x"06",x"ac"),
  1260 => (x"74",x"48",x"ca",x"87"),
  1261 => (x"74",x"4c",x"70",x"88"),
  1262 => (x"72",x"82",x"c1",x"4a"),
  1263 => (x"27",x"30",x"c1",x"48"),
  1264 => (x"00",x"00",x"1c",x"2c"),
  1265 => (x"c0",x"48",x"74",x"58"),
  1266 => (x"c0",x"ff",x"80",x"f0"),
  1267 => (x"c8",x"79",x"70",x"49"),
  1268 => (x"30",x"27",x"87",x"e2"),
  1269 => (x"bf",x"00",x"00",x"1c"),
  1270 => (x"a9",x"b7",x"c9",x"49"),
  1271 => (x"87",x"d4",x"c8",x"01"),
  1272 => (x"00",x"1c",x"30",x"27"),
  1273 => (x"c0",x"49",x"bf",x"00"),
  1274 => (x"c8",x"06",x"a9",x"b7"),
  1275 => (x"30",x"27",x"87",x"c6"),
  1276 => (x"bf",x"00",x"00",x"1c"),
  1277 => (x"80",x"f0",x"c0",x"48"),
  1278 => (x"70",x"49",x"c0",x"ff"),
  1279 => (x"1c",x"20",x"27",x"79"),
  1280 => (x"49",x"bf",x"00",x"00"),
  1281 => (x"01",x"a9",x"b7",x"c3"),
  1282 => (x"97",x"87",x"e9",x"c0"),
  1283 => (x"c1",x"4a",x"66",x"d4"),
  1284 => (x"c0",x"c0",x"c0",x"c0"),
  1285 => (x"b7",x"c0",x"c4",x"92"),
  1286 => (x"1e",x"72",x"4a",x"92"),
  1287 => (x"00",x"1c",x"2c",x"27"),
  1288 => (x"27",x"1e",x"bf",x"00"),
  1289 => (x"00",x"00",x"12",x"e0"),
  1290 => (x"27",x"86",x"c8",x"0f"),
  1291 => (x"00",x"00",x"1c",x"30"),
  1292 => (x"87",x"c0",x"c7",x"58"),
  1293 => (x"00",x"1c",x"28",x"27"),
  1294 => (x"c3",x"4a",x"bf",x"00"),
  1295 => (x"1c",x"20",x"27",x"82"),
  1296 => (x"49",x"bf",x"00",x"00"),
  1297 => (x"01",x"a9",x"b7",x"72"),
  1298 => (x"97",x"87",x"f1",x"c0"),
  1299 => (x"c1",x"4a",x"66",x"d4"),
  1300 => (x"c0",x"c0",x"c0",x"c0"),
  1301 => (x"b7",x"c0",x"c4",x"92"),
  1302 => (x"1e",x"72",x"4a",x"92"),
  1303 => (x"00",x"1c",x"24",x"27"),
  1304 => (x"27",x"1e",x"bf",x"00"),
  1305 => (x"00",x"00",x"12",x"e0"),
  1306 => (x"27",x"86",x"c8",x"0f"),
  1307 => (x"00",x"00",x"1c",x"28"),
  1308 => (x"1c",x"34",x"27",x"58"),
  1309 => (x"c1",x"49",x"00",x"00"),
  1310 => (x"87",x"f8",x"c5",x"79"),
  1311 => (x"00",x"1c",x"30",x"27"),
  1312 => (x"c0",x"49",x"bf",x"00"),
  1313 => (x"c3",x"06",x"a9",x"b7"),
  1314 => (x"30",x"27",x"87",x"d0"),
  1315 => (x"bf",x"00",x"00",x"1c"),
  1316 => (x"a9",x"b7",x"c3",x"49"),
  1317 => (x"87",x"c2",x"c3",x"01"),
  1318 => (x"00",x"1c",x"2c",x"27"),
  1319 => (x"c1",x"4a",x"bf",x"00"),
  1320 => (x"27",x"82",x"c1",x"32"),
  1321 => (x"00",x"00",x"1c",x"20"),
  1322 => (x"b7",x"72",x"49",x"bf"),
  1323 => (x"c2",x"c2",x"01",x"a9"),
  1324 => (x"66",x"d4",x"97",x"87"),
  1325 => (x"c0",x"c0",x"c1",x"4a"),
  1326 => (x"c4",x"92",x"c0",x"c0"),
  1327 => (x"4a",x"92",x"b7",x"c0"),
  1328 => (x"38",x"27",x"1e",x"72"),
  1329 => (x"bf",x"00",x"00",x"1c"),
  1330 => (x"12",x"e0",x"27",x"1e"),
  1331 => (x"c8",x"0f",x"00",x"00"),
  1332 => (x"1c",x"3c",x"27",x"86"),
  1333 => (x"27",x"58",x"00",x"00"),
  1334 => (x"00",x"00",x"1c",x"34"),
  1335 => (x"8a",x"c1",x"4a",x"bf"),
  1336 => (x"00",x"1c",x"34",x"27"),
  1337 => (x"79",x"72",x"49",x"00"),
  1338 => (x"03",x"aa",x"b7",x"c0"),
  1339 => (x"27",x"87",x"c5",x"c4"),
  1340 => (x"00",x"00",x"1c",x"24"),
  1341 => (x"38",x"27",x"4a",x"bf"),
  1342 => (x"97",x"00",x"00",x"1c"),
  1343 => (x"24",x"27",x"52",x"bf"),
  1344 => (x"bf",x"00",x"00",x"1c"),
  1345 => (x"27",x"82",x"c1",x"4a"),
  1346 => (x"00",x"00",x"1c",x"24"),
  1347 => (x"27",x"79",x"72",x"49"),
  1348 => (x"00",x"00",x"1c",x"3c"),
  1349 => (x"06",x"aa",x"b7",x"bf"),
  1350 => (x"27",x"87",x"cd",x"c0"),
  1351 => (x"00",x"00",x"1c",x"3c"),
  1352 => (x"1c",x"24",x"27",x"49"),
  1353 => (x"79",x"bf",x"00",x"00"),
  1354 => (x"00",x"1c",x"34",x"27"),
  1355 => (x"79",x"c1",x"49",x"00"),
  1356 => (x"27",x"87",x"c1",x"c3"),
  1357 => (x"00",x"00",x"1c",x"34"),
  1358 => (x"f7",x"c2",x"05",x"bf"),
  1359 => (x"1c",x"38",x"27",x"87"),
  1360 => (x"4b",x"bf",x"00",x"00"),
  1361 => (x"38",x"27",x"33",x"c4"),
  1362 => (x"49",x"00",x"00",x"1c"),
  1363 => (x"24",x"27",x"79",x"73"),
  1364 => (x"bf",x"00",x"00",x"1c"),
  1365 => (x"c2",x"52",x"73",x"4a"),
  1366 => (x"30",x"27",x"87",x"da"),
  1367 => (x"bf",x"00",x"00",x"1c"),
  1368 => (x"a9",x"b7",x"c7",x"49"),
  1369 => (x"87",x"fd",x"c1",x"04"),
  1370 => (x"f4",x"fe",x"4b",x"c0"),
  1371 => (x"27",x"79",x"c1",x"49"),
  1372 => (x"00",x"00",x"1c",x"3c"),
  1373 => (x"1e",x"75",x"1e",x"bf"),
  1374 => (x"00",x"19",x"85",x"27"),
  1375 => (x"94",x"27",x"1e",x"00"),
  1376 => (x"0f",x"00",x"00",x"00"),
  1377 => (x"24",x"27",x"86",x"cc"),
  1378 => (x"49",x"00",x"00",x"1c"),
  1379 => (x"24",x"27",x"79",x"75"),
  1380 => (x"bf",x"00",x"00",x"1c"),
  1381 => (x"1c",x"3c",x"27",x"49"),
  1382 => (x"b7",x"bf",x"00",x"00"),
  1383 => (x"e5",x"c0",x"03",x"a9"),
  1384 => (x"1c",x"24",x"27",x"87"),
  1385 => (x"bf",x"bf",x"00",x"00"),
  1386 => (x"1c",x"24",x"27",x"83"),
  1387 => (x"4a",x"bf",x"00",x"00"),
  1388 => (x"24",x"27",x"82",x"c4"),
  1389 => (x"49",x"00",x"00",x"1c"),
  1390 => (x"3c",x"27",x"79",x"72"),
  1391 => (x"bf",x"00",x"00",x"1c"),
  1392 => (x"ff",x"04",x"aa",x"b7"),
  1393 => (x"1e",x"73",x"87",x"db"),
  1394 => (x"00",x"19",x"a4",x"27"),
  1395 => (x"94",x"27",x"1e",x"00"),
  1396 => (x"0f",x"00",x"00",x"00"),
  1397 => (x"c0",x"ff",x"86",x"c8"),
  1398 => (x"79",x"c2",x"c1",x"49"),
  1399 => (x"00",x"12",x"ce",x"27"),
  1400 => (x"cf",x"c0",x"0f",x"00"),
  1401 => (x"1c",x"30",x"27",x"87"),
  1402 => (x"48",x"bf",x"00",x"00"),
  1403 => (x"ff",x"80",x"f0",x"c0"),
  1404 => (x"79",x"70",x"49",x"c0"),
  1405 => (x"4c",x"26",x"4d",x"26"),
  1406 => (x"4a",x"26",x"4b",x"26"),
  1407 => (x"ff",x"1e",x"4f",x"26"),
  1408 => (x"4f",x"26",x"87",x"fd"),
  1409 => (x"5b",x"5a",x"5e",x"0e"),
  1410 => (x"27",x"0e",x"5d",x"5c"),
  1411 => (x"00",x"00",x"17",x"ec"),
  1412 => (x"00",x"5e",x"27",x"1e"),
  1413 => (x"c4",x"0f",x"00",x"00"),
  1414 => (x"04",x"fa",x"27",x"86"),
  1415 => (x"70",x"0f",x"00",x"00"),
  1416 => (x"02",x"9a",x"72",x"4a"),
  1417 => (x"27",x"87",x"ce",x"c4"),
  1418 => (x"00",x"00",x"17",x"c9"),
  1419 => (x"00",x"5e",x"27",x"1e"),
  1420 => (x"c4",x"0f",x"00",x"00"),
  1421 => (x"0a",x"bb",x"27",x"86"),
  1422 => (x"27",x"0f",x"00",x"00"),
  1423 => (x"00",x"00",x"1c",x"40"),
  1424 => (x"17",x"e0",x"27",x"1e"),
  1425 => (x"27",x"1e",x"00",x"00"),
  1426 => (x"00",x"00",x"11",x"7a"),
  1427 => (x"70",x"86",x"c8",x"0f"),
  1428 => (x"02",x"9a",x"72",x"4a"),
  1429 => (x"27",x"87",x"d0",x"c3"),
  1430 => (x"00",x"00",x"1c",x"40"),
  1431 => (x"17",x"9e",x"27",x"4b"),
  1432 => (x"27",x"1e",x"00",x"00"),
  1433 => (x"00",x"00",x"00",x"5e"),
  1434 => (x"c0",x"86",x"c4",x"0f"),
  1435 => (x"74",x"4c",x"13",x"4d"),
  1436 => (x"b7",x"e0",x"c0",x"4a"),
  1437 => (x"ed",x"c1",x"02",x"aa"),
  1438 => (x"ff",x"48",x"74",x"87"),
  1439 => (x"79",x"70",x"49",x"c0"),
  1440 => (x"e3",x"c0",x"4a",x"74"),
  1441 => (x"c1",x"02",x"aa",x"b7"),
  1442 => (x"4a",x"74",x"87",x"dc"),
  1443 => (x"aa",x"b7",x"c7",x"c1"),
  1444 => (x"87",x"c6",x"c0",x"05"),
  1445 => (x"00",x"12",x"ce",x"27"),
  1446 => (x"4a",x"74",x"0f",x"00"),
  1447 => (x"05",x"aa",x"b7",x"ca"),
  1448 => (x"27",x"87",x"c6",x"c0"),
  1449 => (x"00",x"00",x"15",x"fe"),
  1450 => (x"c1",x"4a",x"74",x"0f"),
  1451 => (x"05",x"aa",x"b7",x"cc"),
  1452 => (x"27",x"87",x"c6",x"c0"),
  1453 => (x"00",x"00",x"1c",x"40"),
  1454 => (x"ff",x"4a",x"74",x"4b"),
  1455 => (x"8a",x"d0",x"9a",x"df"),
  1456 => (x"4a",x"74",x"4c",x"72"),
  1457 => (x"aa",x"b7",x"f9",x"c0"),
  1458 => (x"87",x"c6",x"c0",x"04"),
  1459 => (x"8a",x"d1",x"4a",x"74"),
  1460 => (x"35",x"c4",x"4c",x"72"),
  1461 => (x"4d",x"75",x"4a",x"74"),
  1462 => (x"4c",x"13",x"b5",x"72"),
  1463 => (x"e0",x"c0",x"4a",x"74"),
  1464 => (x"fe",x"05",x"aa",x"b7"),
  1465 => (x"4a",x"74",x"87",x"d3"),
  1466 => (x"aa",x"b7",x"e3",x"c0"),
  1467 => (x"87",x"e2",x"c0",x"02"),
  1468 => (x"e0",x"c0",x"4a",x"13"),
  1469 => (x"c0",x"05",x"aa",x"b7"),
  1470 => (x"4a",x"13",x"87",x"ca"),
  1471 => (x"aa",x"b7",x"e0",x"c0"),
  1472 => (x"87",x"f6",x"ff",x"02"),
  1473 => (x"1e",x"75",x"8b",x"c1"),
  1474 => (x"7a",x"27",x"1e",x"73"),
  1475 => (x"0f",x"00",x"00",x"11"),
  1476 => (x"4a",x"13",x"86",x"c8"),
  1477 => (x"02",x"aa",x"b7",x"ca"),
  1478 => (x"13",x"87",x"d0",x"fd"),
  1479 => (x"aa",x"b7",x"ca",x"4a"),
  1480 => (x"87",x"f7",x"ff",x"05"),
  1481 => (x"27",x"87",x"c4",x"fd"),
  1482 => (x"00",x"00",x"17",x"b0"),
  1483 => (x"00",x"5e",x"27",x"1e"),
  1484 => (x"c4",x"0f",x"00",x"00"),
  1485 => (x"18",x"02",x"27",x"86"),
  1486 => (x"27",x"1e",x"00",x"00"),
  1487 => (x"00",x"00",x"00",x"5e"),
  1488 => (x"27",x"86",x"c4",x"0f"),
  1489 => (x"00",x"00",x"1c",x"3c"),
  1490 => (x"c3",x"79",x"c0",x"49"),
  1491 => (x"4d",x"ff",x"c8",x"f4"),
  1492 => (x"27",x"1e",x"ee",x"c0"),
  1493 => (x"00",x"00",x"00",x"3f"),
  1494 => (x"75",x"86",x"c4",x"0f"),
  1495 => (x"c9",x"f4",x"c3",x"4b"),
  1496 => (x"c0",x"ff",x"4d",x"c0"),
  1497 => (x"4a",x"74",x"4c",x"bf"),
  1498 => (x"72",x"9a",x"c0",x"c8"),
  1499 => (x"d1",x"c0",x"02",x"9a"),
  1500 => (x"c3",x"4a",x"74",x"87"),
  1501 => (x"1e",x"72",x"9a",x"ff"),
  1502 => (x"00",x"13",x"0d",x"27"),
  1503 => (x"86",x"c4",x"0f",x"00"),
  1504 => (x"4a",x"73",x"4b",x"75"),
  1505 => (x"9a",x"72",x"8b",x"c1"),
  1506 => (x"87",x"d6",x"ff",x"05"),
  1507 => (x"ff",x"c8",x"f4",x"c3"),
  1508 => (x"87",x"fc",x"fe",x"4d"),
  1509 => (x"4c",x"26",x"4d",x"26"),
  1510 => (x"4a",x"26",x"4b",x"26"),
  1511 => (x"61",x"50",x"4f",x"26"),
  1512 => (x"6e",x"69",x"73",x"72"),
  1513 => (x"61",x"6d",x"20",x"67"),
  1514 => (x"65",x"66",x"69",x"6e"),
  1515 => (x"00",x"0a",x"74",x"73"),
  1516 => (x"64",x"61",x"6f",x"4c"),
  1517 => (x"20",x"67",x"6e",x"69"),
  1518 => (x"69",x"6e",x"61",x"6d"),
  1519 => (x"74",x"73",x"65",x"66"),
  1520 => (x"69",x"61",x"66",x"20"),
  1521 => (x"0a",x"64",x"65",x"6c"),
  1522 => (x"6e",x"75",x"48",x"00"),
  1523 => (x"67",x"6e",x"69",x"74"),
  1524 => (x"72",x"6f",x"66",x"20"),
  1525 => (x"72",x"61",x"70",x"20"),
  1526 => (x"69",x"74",x"69",x"74"),
  1527 => (x"00",x"0a",x"6e",x"6f"),
  1528 => (x"49",x"4e",x"41",x"4d"),
  1529 => (x"54",x"53",x"45",x"46"),
  1530 => (x"00",x"54",x"53",x"4d"),
  1531 => (x"74",x"69",x"6e",x"49"),
  1532 => (x"69",x"6c",x"61",x"69"),
  1533 => (x"67",x"6e",x"69",x"7a"),
  1534 => (x"20",x"44",x"53",x"20"),
  1535 => (x"64",x"72",x"61",x"63"),
  1536 => (x"6f",x"42",x"00",x"0a"),
  1537 => (x"6e",x"69",x"74",x"6f"),
  1538 => (x"72",x"66",x"20",x"67"),
  1539 => (x"52",x"20",x"6d",x"6f"),
  1540 => (x"32",x"33",x"32",x"53"),
  1541 => (x"4d",x"43",x"00",x"2e"),
  1542 => (x"65",x"52",x"00",x"44"),
  1543 => (x"6f",x"20",x"64",x"61"),
  1544 => (x"42",x"4d",x"20",x"66"),
  1545 => (x"61",x"66",x"20",x"52"),
  1546 => (x"64",x"65",x"6c",x"69"),
  1547 => (x"6f",x"4e",x"00",x"0a"),
  1548 => (x"72",x"61",x"70",x"20"),
  1549 => (x"69",x"74",x"69",x"74"),
  1550 => (x"73",x"20",x"6e",x"6f"),
  1551 => (x"61",x"6e",x"67",x"69"),
  1552 => (x"65",x"72",x"75",x"74"),
  1553 => (x"75",x"6f",x"66",x"20"),
  1554 => (x"00",x"0a",x"64",x"6e"),
  1555 => (x"73",x"52",x"42",x"4d"),
  1556 => (x"3a",x"65",x"7a",x"69"),
  1557 => (x"2c",x"64",x"25",x"20"),
  1558 => (x"72",x"61",x"70",x"20"),
  1559 => (x"69",x"74",x"69",x"74"),
  1560 => (x"69",x"73",x"6e",x"6f"),
  1561 => (x"20",x"3a",x"65",x"7a"),
  1562 => (x"20",x"2c",x"64",x"25"),
  1563 => (x"73",x"66",x"66",x"6f"),
  1564 => (x"6f",x"20",x"74",x"65"),
  1565 => (x"69",x"73",x"20",x"66"),
  1566 => (x"25",x"20",x"3a",x"67"),
  1567 => (x"73",x"20",x"2c",x"64"),
  1568 => (x"30",x"20",x"67",x"69"),
  1569 => (x"0a",x"78",x"25",x"78"),
  1570 => (x"61",x"65",x"52",x"00"),
  1571 => (x"67",x"6e",x"69",x"64"),
  1572 => (x"6f",x"6f",x"62",x"20"),
  1573 => (x"65",x"73",x"20",x"74"),
  1574 => (x"72",x"6f",x"74",x"63"),
  1575 => (x"0a",x"64",x"25",x"20"),
  1576 => (x"61",x"65",x"52",x"00"),
  1577 => (x"6f",x"62",x"20",x"64"),
  1578 => (x"73",x"20",x"74",x"6f"),
  1579 => (x"6f",x"74",x"63",x"65"),
  1580 => (x"72",x"66",x"20",x"72"),
  1581 => (x"66",x"20",x"6d",x"6f"),
  1582 => (x"74",x"73",x"72",x"69"),
  1583 => (x"72",x"61",x"70",x"20"),
  1584 => (x"69",x"74",x"69",x"74"),
  1585 => (x"00",x"0a",x"6e",x"6f"),
  1586 => (x"75",x"73",x"6e",x"55"),
  1587 => (x"72",x"6f",x"70",x"70"),
  1588 => (x"20",x"64",x"65",x"74"),
  1589 => (x"74",x"72",x"61",x"70"),
  1590 => (x"6f",x"69",x"74",x"69"),
  1591 => (x"79",x"74",x"20",x"6e"),
  1592 => (x"0d",x"21",x"65",x"70"),
  1593 => (x"54",x"41",x"46",x"00"),
  1594 => (x"20",x"20",x"32",x"33"),
  1595 => (x"65",x"52",x"00",x"20"),
  1596 => (x"6e",x"69",x"64",x"61"),
  1597 => (x"42",x"4d",x"20",x"67"),
  1598 => (x"4d",x"00",x"0a",x"52"),
  1599 => (x"73",x"20",x"52",x"42"),
  1600 => (x"65",x"63",x"63",x"75"),
  1601 => (x"75",x"66",x"73",x"73"),
  1602 => (x"20",x"79",x"6c",x"6c"),
  1603 => (x"64",x"61",x"65",x"72"),
  1604 => (x"41",x"46",x"00",x"0a"),
  1605 => (x"20",x"36",x"31",x"54"),
  1606 => (x"46",x"00",x"20",x"20"),
  1607 => (x"32",x"33",x"54",x"41"),
  1608 => (x"00",x"20",x"20",x"20"),
  1609 => (x"74",x"72",x"61",x"50"),
  1610 => (x"6f",x"69",x"74",x"69"),
  1611 => (x"75",x"6f",x"63",x"6e"),
  1612 => (x"25",x"20",x"74",x"6e"),
  1613 => (x"48",x"00",x"0a",x"64"),
  1614 => (x"69",x"74",x"6e",x"75"),
  1615 => (x"66",x"20",x"67",x"6e"),
  1616 => (x"66",x"20",x"72",x"6f"),
  1617 => (x"73",x"65",x"6c",x"69"),
  1618 => (x"65",x"74",x"73",x"79"),
  1619 => (x"46",x"00",x"0a",x"6d"),
  1620 => (x"32",x"33",x"54",x"41"),
  1621 => (x"00",x"20",x"20",x"20"),
  1622 => (x"31",x"54",x"41",x"46"),
  1623 => (x"20",x"20",x"20",x"36"),
  1624 => (x"75",x"6c",x"43",x"00"),
  1625 => (x"72",x"65",x"74",x"73"),
  1626 => (x"7a",x"69",x"73",x"20"),
  1627 => (x"25",x"20",x"3a",x"65"),
  1628 => (x"43",x"20",x"2c",x"64"),
  1629 => (x"74",x"73",x"75",x"6c"),
  1630 => (x"6d",x"20",x"72",x"65"),
  1631 => (x"2c",x"6b",x"73",x"61"),
  1632 => (x"0a",x"64",x"25",x"20"),
  1633 => (x"65",x"68",x"43",x"00"),
  1634 => (x"75",x"73",x"6b",x"63"),
  1635 => (x"6e",x"69",x"6d",x"6d"),
  1636 => (x"72",x"66",x"20",x"67"),
  1637 => (x"25",x"20",x"6d",x"6f"),
  1638 => (x"6f",x"74",x"20",x"64"),
  1639 => (x"2e",x"64",x"25",x"20"),
  1640 => (x"00",x"20",x"2e",x"2e"),
  1641 => (x"00",x"0a",x"64",x"25"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
