
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"d4",x"01"),
     1 => (x"18",x"0e",x"87",x"d7"),
     2 => (x"3e",x"27",x"0e",x"1e"),
     3 => (x"0f",x"00",x"00",x"00"),
     4 => (x"80",x"ff",x"48",x"26"),
     5 => (x"27",x"4f",x"08",x"26"),
     6 => (x"00",x"00",x"00",x"23"),
     7 => (x"00",x"30",x"27",x"4f"),
     8 => (x"c2",x"4f",x"00",x"00"),
     9 => (x"27",x"4e",x"c0",x"c0"),
    10 => (x"00",x"00",x"16",x"03"),
    11 => (x"87",x"fd",x"00",x"0f"),
    12 => (x"4e",x"c0",x"f0",x"c1"),
    13 => (x"00",x"00",x"3d",x"27"),
    14 => (x"fd",x"00",x"0f",x"00"),
    15 => (x"1e",x"4f",x"4f",x"87"),
    16 => (x"ff",x"1e",x"1e",x"72"),
    17 => (x"48",x"6a",x"4a",x"c0"),
    18 => (x"c4",x"98",x"c0",x"c4"),
    19 => (x"02",x"6e",x"58",x"a6"),
    20 => (x"cc",x"87",x"f3",x"ff"),
    21 => (x"66",x"cc",x"7a",x"66"),
    22 => (x"4a",x"26",x"26",x"48"),
    23 => (x"5e",x"0e",x"4f",x"26"),
    24 => (x"5d",x"5c",x"5b",x"5a"),
    25 => (x"4b",x"66",x"d4",x"0e"),
    26 => (x"4c",x"13",x"4d",x"c0"),
    27 => (x"c0",x"02",x"9c",x"74"),
    28 => (x"4a",x"74",x"87",x"d6"),
    29 => (x"3f",x"27",x"1e",x"72"),
    30 => (x"0f",x"00",x"00",x"00"),
    31 => (x"85",x"c1",x"86",x"c4"),
    32 => (x"9c",x"74",x"4c",x"13"),
    33 => (x"87",x"ea",x"ff",x"05"),
    34 => (x"4d",x"26",x"48",x"75"),
    35 => (x"4b",x"26",x"4c",x"26"),
    36 => (x"4f",x"26",x"4a",x"26"),
    37 => (x"5b",x"5a",x"5e",x"0e"),
    38 => (x"d0",x"0e",x"5d",x"5c"),
    39 => (x"c4",x"4c",x"c0",x"8e"),
    40 => (x"79",x"c0",x"49",x"a6"),
    41 => (x"4b",x"a6",x"e8",x"c0"),
    42 => (x"4a",x"66",x"e4",x"c0"),
    43 => (x"48",x"66",x"e4",x"c0"),
    44 => (x"e8",x"c0",x"80",x"c1"),
    45 => (x"48",x"12",x"58",x"a6"),
    46 => (x"c0",x"c0",x"c0",x"c1"),
    47 => (x"c0",x"c4",x"90",x"c0"),
    48 => (x"c4",x"48",x"90",x"b7"),
    49 => (x"02",x"6e",x"58",x"a6"),
    50 => (x"c4",x"87",x"c2",x"c5"),
    51 => (x"fe",x"c3",x"02",x"66"),
    52 => (x"49",x"a6",x"c4",x"87"),
    53 => (x"4a",x"6e",x"79",x"c0"),
    54 => (x"f0",x"c0",x"49",x"6e"),
    55 => (x"c4",x"c3",x"02",x"a9"),
    56 => (x"aa",x"e3",x"c1",x"87"),
    57 => (x"87",x"c5",x"c3",x"02"),
    58 => (x"02",x"aa",x"e4",x"c1"),
    59 => (x"c1",x"87",x"e3",x"c0"),
    60 => (x"c2",x"02",x"aa",x"ec"),
    61 => (x"f0",x"c1",x"87",x"ef"),
    62 => (x"d5",x"c0",x"02",x"aa"),
    63 => (x"aa",x"f3",x"c1",x"87"),
    64 => (x"87",x"c8",x"c2",x"02"),
    65 => (x"02",x"aa",x"f5",x"c1"),
    66 => (x"c1",x"87",x"c7",x"c0"),
    67 => (x"c2",x"05",x"aa",x"f8"),
    68 => (x"83",x"c4",x"87",x"f0"),
    69 => (x"8a",x"c4",x"4a",x"73"),
    70 => (x"79",x"6a",x"49",x"76"),
    71 => (x"db",x"c1",x"02",x"6e"),
    72 => (x"49",x"a6",x"c8",x"87"),
    73 => (x"a6",x"cc",x"79",x"c0"),
    74 => (x"6e",x"79",x"c0",x"49"),
    75 => (x"2a",x"b7",x"dc",x"4a"),
    76 => (x"9d",x"cf",x"4d",x"72"),
    77 => (x"30",x"c4",x"48",x"6e"),
    78 => (x"75",x"58",x"a6",x"c4"),
    79 => (x"c5",x"c0",x"02",x"9d"),
    80 => (x"49",x"a6",x"c8",x"87"),
    81 => (x"ad",x"c9",x"79",x"c1"),
    82 => (x"87",x"c6",x"c0",x"06"),
    83 => (x"c0",x"85",x"f7",x"c0"),
    84 => (x"f0",x"c0",x"87",x"c3"),
    85 => (x"02",x"66",x"c8",x"85"),
    86 => (x"75",x"87",x"cc",x"c0"),
    87 => (x"00",x"3f",x"27",x"1e"),
    88 => (x"c4",x"0f",x"00",x"00"),
    89 => (x"cc",x"84",x"c1",x"86"),
    90 => (x"80",x"c1",x"48",x"66"),
    91 => (x"cc",x"58",x"a6",x"d0"),
    92 => (x"b7",x"c8",x"49",x"66"),
    93 => (x"f2",x"fe",x"04",x"a9"),
    94 => (x"87",x"ee",x"c1",x"87"),
    95 => (x"27",x"1e",x"f0",x"c0"),
    96 => (x"00",x"00",x"00",x"3f"),
    97 => (x"c1",x"86",x"c4",x"0f"),
    98 => (x"87",x"de",x"c1",x"84"),
    99 => (x"4a",x"73",x"83",x"c4"),
   100 => (x"1e",x"6a",x"8a",x"c4"),
   101 => (x"00",x"00",x"5e",x"27"),
   102 => (x"86",x"c4",x"0f",x"00"),
   103 => (x"4c",x"74",x"4a",x"70"),
   104 => (x"c5",x"c1",x"84",x"72"),
   105 => (x"49",x"a6",x"c4",x"87"),
   106 => (x"fd",x"c0",x"79",x"c1"),
   107 => (x"73",x"83",x"c4",x"87"),
   108 => (x"6a",x"8a",x"c4",x"4a"),
   109 => (x"00",x"3f",x"27",x"1e"),
   110 => (x"c4",x"0f",x"00",x"00"),
   111 => (x"c0",x"84",x"c1",x"86"),
   112 => (x"1e",x"6e",x"87",x"e8"),
   113 => (x"00",x"00",x"3f",x"27"),
   114 => (x"86",x"c4",x"0f",x"00"),
   115 => (x"6e",x"87",x"db",x"c0"),
   116 => (x"a9",x"e5",x"c0",x"49"),
   117 => (x"87",x"c8",x"c0",x"05"),
   118 => (x"c1",x"49",x"a6",x"c4"),
   119 => (x"87",x"ca",x"c0",x"79"),
   120 => (x"3f",x"27",x"1e",x"6e"),
   121 => (x"0f",x"00",x"00",x"00"),
   122 => (x"e4",x"c0",x"86",x"c4"),
   123 => (x"e4",x"c0",x"4a",x"66"),
   124 => (x"80",x"c1",x"48",x"66"),
   125 => (x"58",x"a6",x"e8",x"c0"),
   126 => (x"c0",x"c1",x"48",x"12"),
   127 => (x"90",x"c0",x"c0",x"c0"),
   128 => (x"90",x"b7",x"c0",x"c4"),
   129 => (x"58",x"a6",x"c4",x"48"),
   130 => (x"fe",x"fa",x"05",x"6e"),
   131 => (x"d0",x"48",x"74",x"87"),
   132 => (x"26",x"4d",x"26",x"86"),
   133 => (x"26",x"4b",x"26",x"4c"),
   134 => (x"00",x"4f",x"26",x"4a"),
   135 => (x"1e",x"00",x"00",x"00"),
   136 => (x"d4",x"ff",x"1e",x"75"),
   137 => (x"49",x"ff",x"c3",x"4d"),
   138 => (x"c8",x"48",x"6d",x"7d"),
   139 => (x"6d",x"7d",x"71",x"38"),
   140 => (x"71",x"38",x"c8",x"b0"),
   141 => (x"c8",x"b0",x"6d",x"7d"),
   142 => (x"6d",x"7d",x"71",x"38"),
   143 => (x"26",x"38",x"c8",x"b0"),
   144 => (x"1e",x"4f",x"26",x"4d"),
   145 => (x"d4",x"ff",x"1e",x"75"),
   146 => (x"49",x"ff",x"c3",x"4d"),
   147 => (x"c8",x"48",x"6d",x"7d"),
   148 => (x"6d",x"7d",x"71",x"30"),
   149 => (x"71",x"30",x"c8",x"b0"),
   150 => (x"c8",x"b0",x"6d",x"7d"),
   151 => (x"6d",x"7d",x"71",x"30"),
   152 => (x"26",x"4d",x"26",x"b0"),
   153 => (x"1e",x"75",x"1e",x"4f"),
   154 => (x"cc",x"4d",x"d4",x"ff"),
   155 => (x"66",x"c8",x"49",x"66"),
   156 => (x"e6",x"fe",x"7d",x"48"),
   157 => (x"31",x"c9",x"02",x"67"),
   158 => (x"09",x"39",x"d8",x"07"),
   159 => (x"09",x"39",x"09",x"7d"),
   160 => (x"09",x"39",x"09",x"7d"),
   161 => (x"09",x"39",x"09",x"7d"),
   162 => (x"70",x"38",x"d0",x"7d"),
   163 => (x"c0",x"f1",x"c9",x"7d"),
   164 => (x"48",x"ff",x"c3",x"49"),
   165 => (x"05",x"a8",x"08",x"6d"),
   166 => (x"7d",x"08",x"87",x"c7"),
   167 => (x"f3",x"05",x"89",x"c1"),
   168 => (x"26",x"4d",x"26",x"87"),
   169 => (x"d4",x"ff",x"1e",x"4f"),
   170 => (x"48",x"c8",x"c3",x"49"),
   171 => (x"05",x"80",x"79",x"ff"),
   172 => (x"4f",x"26",x"87",x"fa"),
   173 => (x"5b",x"5a",x"5e",x"0e"),
   174 => (x"c0",x"0e",x"5d",x"5c"),
   175 => (x"f7",x"c1",x"f0",x"ff"),
   176 => (x"c0",x"c0",x"c1",x"4d"),
   177 => (x"4b",x"c0",x"c0",x"c0"),
   178 => (x"00",x"02",x"a5",x"27"),
   179 => (x"f8",x"c4",x"0f",x"00"),
   180 => (x"1e",x"c0",x"4c",x"df"),
   181 => (x"65",x"27",x"1e",x"75"),
   182 => (x"0f",x"00",x"00",x"02"),
   183 => (x"4a",x"70",x"86",x"c8"),
   184 => (x"05",x"aa",x"b7",x"c1"),
   185 => (x"ff",x"87",x"ef",x"c0"),
   186 => (x"ff",x"c3",x"49",x"d4"),
   187 => (x"c0",x"1e",x"73",x"79"),
   188 => (x"e9",x"c1",x"f0",x"e1"),
   189 => (x"02",x"65",x"27",x"1e"),
   190 => (x"c8",x"0f",x"00",x"00"),
   191 => (x"72",x"4a",x"70",x"86"),
   192 => (x"cb",x"c0",x"05",x"9a"),
   193 => (x"49",x"d4",x"ff",x"87"),
   194 => (x"c1",x"79",x"ff",x"c3"),
   195 => (x"87",x"d0",x"c0",x"48"),
   196 => (x"00",x"02",x"a5",x"27"),
   197 => (x"8c",x"c1",x"0f",x"00"),
   198 => (x"fe",x"05",x"9c",x"74"),
   199 => (x"48",x"c0",x"87",x"f4"),
   200 => (x"4c",x"26",x"4d",x"26"),
   201 => (x"4a",x"26",x"4b",x"26"),
   202 => (x"5e",x"0e",x"4f",x"26"),
   203 => (x"0e",x"5c",x"5b",x"5a"),
   204 => (x"c1",x"f0",x"ff",x"c0"),
   205 => (x"d4",x"ff",x"4c",x"c1"),
   206 => (x"79",x"ff",x"c3",x"49"),
   207 => (x"00",x"18",x"15",x"27"),
   208 => (x"5e",x"27",x"1e",x"00"),
   209 => (x"0f",x"00",x"00",x"00"),
   210 => (x"4b",x"d3",x"86",x"c4"),
   211 => (x"1e",x"74",x"1e",x"c0"),
   212 => (x"00",x"02",x"65",x"27"),
   213 => (x"86",x"c8",x"0f",x"00"),
   214 => (x"9a",x"72",x"4a",x"70"),
   215 => (x"87",x"cb",x"c0",x"05"),
   216 => (x"c3",x"49",x"d4",x"ff"),
   217 => (x"48",x"c1",x"79",x"ff"),
   218 => (x"27",x"87",x"d0",x"c0"),
   219 => (x"00",x"00",x"02",x"a5"),
   220 => (x"73",x"8b",x"c1",x"0f"),
   221 => (x"d3",x"ff",x"05",x"9b"),
   222 => (x"26",x"48",x"c0",x"87"),
   223 => (x"26",x"4b",x"26",x"4c"),
   224 => (x"0e",x"4f",x"26",x"4a"),
   225 => (x"5c",x"5b",x"5a",x"5e"),
   226 => (x"c3",x"1e",x"0e",x"5d"),
   227 => (x"d4",x"ff",x"4d",x"ff"),
   228 => (x"02",x"a5",x"27",x"4c"),
   229 => (x"c6",x"0f",x"00",x"00"),
   230 => (x"e1",x"c0",x"1e",x"ea"),
   231 => (x"1e",x"c8",x"c1",x"f0"),
   232 => (x"00",x"02",x"65",x"27"),
   233 => (x"86",x"c8",x"0f",x"00"),
   234 => (x"1e",x"72",x"4a",x"70"),
   235 => (x"00",x"04",x"e2",x"27"),
   236 => (x"94",x"27",x"1e",x"00"),
   237 => (x"0f",x"00",x"00",x"00"),
   238 => (x"b7",x"c1",x"86",x"c8"),
   239 => (x"cb",x"c0",x"02",x"aa"),
   240 => (x"03",x"2a",x"27",x"87"),
   241 => (x"c0",x"0f",x"00",x"00"),
   242 => (x"87",x"c9",x"c3",x"48"),
   243 => (x"00",x"02",x"43",x"27"),
   244 => (x"4a",x"70",x"0f",x"00"),
   245 => (x"9a",x"ff",x"ff",x"cf"),
   246 => (x"aa",x"b7",x"ea",x"c6"),
   247 => (x"87",x"cb",x"c0",x"02"),
   248 => (x"00",x"03",x"2a",x"27"),
   249 => (x"48",x"c0",x"0f",x"00"),
   250 => (x"75",x"87",x"ea",x"c2"),
   251 => (x"c0",x"49",x"76",x"7c"),
   252 => (x"b4",x"27",x"79",x"f1"),
   253 => (x"0f",x"00",x"00",x"02"),
   254 => (x"9a",x"72",x"4a",x"70"),
   255 => (x"87",x"eb",x"c1",x"02"),
   256 => (x"ff",x"c0",x"1e",x"c0"),
   257 => (x"1e",x"fa",x"c1",x"f0"),
   258 => (x"00",x"02",x"65",x"27"),
   259 => (x"86",x"c8",x"0f",x"00"),
   260 => (x"9b",x"73",x"4b",x"70"),
   261 => (x"87",x"c3",x"c1",x"05"),
   262 => (x"a0",x"27",x"1e",x"73"),
   263 => (x"1e",x"00",x"00",x"04"),
   264 => (x"00",x"00",x"94",x"27"),
   265 => (x"86",x"c8",x"0f",x"00"),
   266 => (x"4b",x"6c",x"7c",x"75"),
   267 => (x"1e",x"73",x"9b",x"75"),
   268 => (x"00",x"04",x"ac",x"27"),
   269 => (x"94",x"27",x"1e",x"00"),
   270 => (x"0f",x"00",x"00",x"00"),
   271 => (x"7c",x"75",x"86",x"c8"),
   272 => (x"7c",x"75",x"7c",x"75"),
   273 => (x"4a",x"73",x"7c",x"75"),
   274 => (x"72",x"9a",x"c0",x"c1"),
   275 => (x"c5",x"c0",x"02",x"9a"),
   276 => (x"c0",x"48",x"c1",x"87"),
   277 => (x"48",x"c0",x"87",x"ff"),
   278 => (x"73",x"87",x"fa",x"c0"),
   279 => (x"04",x"ba",x"27",x"1e"),
   280 => (x"27",x"1e",x"00",x"00"),
   281 => (x"00",x"00",x"00",x"94"),
   282 => (x"6e",x"86",x"c8",x"0f"),
   283 => (x"a9",x"b7",x"c2",x"49"),
   284 => (x"87",x"d3",x"c0",x"05"),
   285 => (x"00",x"04",x"c6",x"27"),
   286 => (x"94",x"27",x"1e",x"00"),
   287 => (x"0f",x"00",x"00",x"00"),
   288 => (x"48",x"c0",x"86",x"c4"),
   289 => (x"6e",x"87",x"ce",x"c0"),
   290 => (x"c4",x"88",x"c1",x"48"),
   291 => (x"05",x"6e",x"58",x"a6"),
   292 => (x"c0",x"87",x"df",x"fd"),
   293 => (x"4d",x"26",x"26",x"48"),
   294 => (x"4b",x"26",x"4c",x"26"),
   295 => (x"4f",x"26",x"4a",x"26"),
   296 => (x"35",x"44",x"4d",x"43"),
   297 => (x"64",x"25",x"20",x"38"),
   298 => (x"00",x"20",x"20",x"0a"),
   299 => (x"35",x"44",x"4d",x"43"),
   300 => (x"20",x"32",x"5f",x"38"),
   301 => (x"20",x"0a",x"64",x"25"),
   302 => (x"4d",x"43",x"00",x"20"),
   303 => (x"20",x"38",x"35",x"44"),
   304 => (x"20",x"0a",x"64",x"25"),
   305 => (x"44",x"53",x"00",x"20"),
   306 => (x"49",x"20",x"43",x"48"),
   307 => (x"69",x"74",x"69",x"6e"),
   308 => (x"7a",x"69",x"6c",x"61"),
   309 => (x"6f",x"69",x"74",x"61"),
   310 => (x"72",x"65",x"20",x"6e"),
   311 => (x"21",x"72",x"6f",x"72"),
   312 => (x"6d",x"63",x"00",x"0a"),
   313 => (x"4d",x"43",x"5f",x"64"),
   314 => (x"72",x"20",x"38",x"44"),
   315 => (x"6f",x"70",x"73",x"65"),
   316 => (x"3a",x"65",x"73",x"6e"),
   317 => (x"0a",x"64",x"25",x"20"),
   318 => (x"5a",x"5e",x"0e",x"00"),
   319 => (x"0e",x"5d",x"5c",x"5b"),
   320 => (x"4c",x"d0",x"ff",x"1e"),
   321 => (x"4b",x"c0",x"c0",x"c8"),
   322 => (x"00",x"02",x"1b",x"27"),
   323 => (x"79",x"c1",x"49",x"00"),
   324 => (x"00",x"06",x"16",x"27"),
   325 => (x"5e",x"27",x"1e",x"00"),
   326 => (x"0f",x"00",x"00",x"00"),
   327 => (x"4d",x"c7",x"86",x"c4"),
   328 => (x"98",x"73",x"48",x"6c"),
   329 => (x"6e",x"58",x"a6",x"c4"),
   330 => (x"87",x"cc",x"c0",x"02"),
   331 => (x"98",x"73",x"48",x"6c"),
   332 => (x"6e",x"58",x"a6",x"c4"),
   333 => (x"87",x"f4",x"ff",x"05"),
   334 => (x"a5",x"27",x"7c",x"c0"),
   335 => (x"0f",x"00",x"00",x"02"),
   336 => (x"98",x"73",x"48",x"6c"),
   337 => (x"6e",x"58",x"a6",x"c4"),
   338 => (x"87",x"cc",x"c0",x"02"),
   339 => (x"98",x"73",x"48",x"6c"),
   340 => (x"6e",x"58",x"a6",x"c4"),
   341 => (x"87",x"f4",x"ff",x"05"),
   342 => (x"1e",x"c0",x"7c",x"c1"),
   343 => (x"c1",x"d0",x"e5",x"c0"),
   344 => (x"65",x"27",x"1e",x"c0"),
   345 => (x"0f",x"00",x"00",x"02"),
   346 => (x"4a",x"70",x"86",x"c8"),
   347 => (x"05",x"aa",x"b7",x"c1"),
   348 => (x"c1",x"87",x"c2",x"c0"),
   349 => (x"ad",x"b7",x"c2",x"4d"),
   350 => (x"87",x"d3",x"c0",x"05"),
   351 => (x"00",x"06",x"11",x"27"),
   352 => (x"5e",x"27",x"1e",x"00"),
   353 => (x"0f",x"00",x"00",x"00"),
   354 => (x"48",x"c0",x"86",x"c4"),
   355 => (x"c1",x"87",x"f7",x"c1"),
   356 => (x"05",x"9d",x"75",x"8d"),
   357 => (x"27",x"87",x"c9",x"fe"),
   358 => (x"00",x"00",x"03",x"83"),
   359 => (x"02",x"1f",x"27",x"0f"),
   360 => (x"27",x"58",x"00",x"00"),
   361 => (x"00",x"00",x"02",x"1b"),
   362 => (x"d0",x"c0",x"05",x"bf"),
   363 => (x"c0",x"1e",x"c1",x"87"),
   364 => (x"d0",x"c1",x"f0",x"ff"),
   365 => (x"02",x"65",x"27",x"1e"),
   366 => (x"c8",x"0f",x"00",x"00"),
   367 => (x"49",x"d4",x"ff",x"86"),
   368 => (x"27",x"79",x"ff",x"c3"),
   369 => (x"00",x"00",x"08",x"ac"),
   370 => (x"19",x"b0",x"27",x"0f"),
   371 => (x"27",x"58",x"00",x"00"),
   372 => (x"00",x"00",x"19",x"ac"),
   373 => (x"1a",x"27",x"1e",x"bf"),
   374 => (x"1e",x"00",x"00",x"06"),
   375 => (x"00",x"00",x"94",x"27"),
   376 => (x"86",x"c8",x"0f",x"00"),
   377 => (x"98",x"73",x"48",x"6c"),
   378 => (x"6e",x"58",x"a6",x"c4"),
   379 => (x"87",x"cc",x"c0",x"02"),
   380 => (x"98",x"73",x"48",x"6c"),
   381 => (x"6e",x"58",x"a6",x"c4"),
   382 => (x"87",x"f4",x"ff",x"05"),
   383 => (x"d4",x"ff",x"7c",x"c0"),
   384 => (x"79",x"ff",x"c3",x"49"),
   385 => (x"26",x"26",x"48",x"c1"),
   386 => (x"26",x"4c",x"26",x"4d"),
   387 => (x"26",x"4a",x"26",x"4b"),
   388 => (x"52",x"45",x"49",x"4f"),
   389 => (x"50",x"53",x"00",x"52"),
   390 => (x"44",x"53",x"00",x"49"),
   391 => (x"72",x"61",x"63",x"20"),
   392 => (x"69",x"73",x"20",x"64"),
   393 => (x"69",x"20",x"65",x"7a"),
   394 => (x"64",x"25",x"20",x"73"),
   395 => (x"5e",x"0e",x"00",x"0a"),
   396 => (x"5d",x"5c",x"5b",x"5a"),
   397 => (x"ff",x"c3",x"1e",x"0e"),
   398 => (x"4c",x"d4",x"ff",x"4d"),
   399 => (x"d0",x"ff",x"7c",x"75"),
   400 => (x"c0",x"c8",x"48",x"bf"),
   401 => (x"a6",x"c4",x"98",x"c0"),
   402 => (x"c0",x"02",x"6e",x"58"),
   403 => (x"c0",x"c8",x"87",x"d2"),
   404 => (x"d0",x"ff",x"4a",x"c0"),
   405 => (x"98",x"72",x"48",x"bf"),
   406 => (x"6e",x"58",x"a6",x"c4"),
   407 => (x"87",x"f2",x"ff",x"05"),
   408 => (x"c4",x"49",x"d0",x"ff"),
   409 => (x"7c",x"75",x"79",x"c1"),
   410 => (x"c0",x"1e",x"66",x"d8"),
   411 => (x"d8",x"c1",x"f0",x"ff"),
   412 => (x"02",x"65",x"27",x"1e"),
   413 => (x"c8",x"0f",x"00",x"00"),
   414 => (x"72",x"4a",x"70",x"86"),
   415 => (x"d3",x"c0",x"02",x"9a"),
   416 => (x"07",x"36",x"27",x"87"),
   417 => (x"27",x"1e",x"00",x"00"),
   418 => (x"00",x"00",x"00",x"5e"),
   419 => (x"c1",x"86",x"c4",x"0f"),
   420 => (x"87",x"d7",x"c2",x"48"),
   421 => (x"fe",x"c3",x"7c",x"75"),
   422 => (x"c0",x"49",x"76",x"7c"),
   423 => (x"bf",x"66",x"dc",x"79"),
   424 => (x"d8",x"4b",x"72",x"4a"),
   425 => (x"48",x"73",x"2b",x"b7"),
   426 => (x"7c",x"70",x"98",x"75"),
   427 => (x"b7",x"d0",x"4b",x"72"),
   428 => (x"75",x"48",x"73",x"2b"),
   429 => (x"72",x"7c",x"70",x"98"),
   430 => (x"2b",x"b7",x"c8",x"4b"),
   431 => (x"98",x"75",x"48",x"73"),
   432 => (x"48",x"72",x"7c",x"70"),
   433 => (x"7c",x"70",x"98",x"75"),
   434 => (x"c4",x"48",x"66",x"dc"),
   435 => (x"a6",x"e0",x"c0",x"80"),
   436 => (x"c1",x"48",x"6e",x"58"),
   437 => (x"58",x"a6",x"c4",x"80"),
   438 => (x"c0",x"c2",x"49",x"6e"),
   439 => (x"fe",x"04",x"a9",x"b7"),
   440 => (x"7c",x"75",x"87",x"fb"),
   441 => (x"7c",x"75",x"7c",x"75"),
   442 => (x"4b",x"e0",x"da",x"d8"),
   443 => (x"4a",x"6c",x"7c",x"75"),
   444 => (x"9a",x"72",x"9a",x"75"),
   445 => (x"87",x"c8",x"c0",x"05"),
   446 => (x"9b",x"73",x"8b",x"c1"),
   447 => (x"87",x"ec",x"ff",x"05"),
   448 => (x"d0",x"ff",x"7c",x"75"),
   449 => (x"c0",x"c8",x"48",x"bf"),
   450 => (x"a6",x"c4",x"98",x"c0"),
   451 => (x"c0",x"02",x"6e",x"58"),
   452 => (x"c0",x"c8",x"87",x"d2"),
   453 => (x"d0",x"ff",x"4a",x"c0"),
   454 => (x"98",x"72",x"48",x"bf"),
   455 => (x"6e",x"58",x"a6",x"c4"),
   456 => (x"87",x"f2",x"ff",x"05"),
   457 => (x"c0",x"49",x"d0",x"ff"),
   458 => (x"26",x"48",x"c0",x"79"),
   459 => (x"4c",x"26",x"4d",x"26"),
   460 => (x"4a",x"26",x"4b",x"26"),
   461 => (x"72",x"57",x"4f",x"26"),
   462 => (x"20",x"65",x"74",x"69"),
   463 => (x"6c",x"69",x"61",x"66"),
   464 => (x"00",x"0a",x"64",x"65"),
   465 => (x"5b",x"5a",x"5e",x"0e"),
   466 => (x"1e",x"0e",x"5d",x"5c"),
   467 => (x"dc",x"4c",x"66",x"d8"),
   468 => (x"49",x"76",x"4b",x"66"),
   469 => (x"ee",x"c5",x"79",x"c0"),
   470 => (x"ff",x"4d",x"df",x"cd"),
   471 => (x"ff",x"c3",x"49",x"d4"),
   472 => (x"bf",x"d4",x"ff",x"79"),
   473 => (x"9a",x"ff",x"c3",x"4a"),
   474 => (x"aa",x"b7",x"fe",x"c3"),
   475 => (x"87",x"e5",x"c1",x"05"),
   476 => (x"00",x"19",x"a8",x"27"),
   477 => (x"79",x"c0",x"49",x"00"),
   478 => (x"04",x"ab",x"b7",x"c4"),
   479 => (x"27",x"87",x"e4",x"c0"),
   480 => (x"00",x"00",x"02",x"1f"),
   481 => (x"72",x"4a",x"70",x"0f"),
   482 => (x"27",x"84",x"c4",x"7c"),
   483 => (x"00",x"00",x"19",x"a8"),
   484 => (x"80",x"72",x"48",x"bf"),
   485 => (x"00",x"19",x"ac",x"27"),
   486 => (x"8b",x"c4",x"58",x"00"),
   487 => (x"03",x"ab",x"b7",x"c4"),
   488 => (x"c0",x"87",x"dc",x"ff"),
   489 => (x"c0",x"06",x"ab",x"b7"),
   490 => (x"d4",x"ff",x"87",x"e5"),
   491 => (x"7d",x"ff",x"c3",x"4d"),
   492 => (x"97",x"72",x"4a",x"6d"),
   493 => (x"27",x"84",x"c1",x"7c"),
   494 => (x"00",x"00",x"19",x"a8"),
   495 => (x"80",x"72",x"48",x"bf"),
   496 => (x"00",x"19",x"ac",x"27"),
   497 => (x"8b",x"c1",x"58",x"00"),
   498 => (x"01",x"ab",x"b7",x"c0"),
   499 => (x"c1",x"87",x"de",x"ff"),
   500 => (x"c1",x"49",x"76",x"4d"),
   501 => (x"75",x"8d",x"c1",x"79"),
   502 => (x"fe",x"fd",x"05",x"9d"),
   503 => (x"49",x"d4",x"ff",x"87"),
   504 => (x"6e",x"79",x"ff",x"c3"),
   505 => (x"4d",x"26",x"26",x"48"),
   506 => (x"4b",x"26",x"4c",x"26"),
   507 => (x"4f",x"26",x"4a",x"26"),
   508 => (x"5b",x"5a",x"5e",x"0e"),
   509 => (x"1e",x"0e",x"5d",x"5c"),
   510 => (x"c8",x"4b",x"d0",x"ff"),
   511 => (x"c0",x"4a",x"c0",x"c0"),
   512 => (x"49",x"d4",x"ff",x"4c"),
   513 => (x"6b",x"79",x"ff",x"c3"),
   514 => (x"c4",x"98",x"72",x"48"),
   515 => (x"02",x"6e",x"58",x"a6"),
   516 => (x"6b",x"87",x"cc",x"c0"),
   517 => (x"c4",x"98",x"72",x"48"),
   518 => (x"05",x"6e",x"58",x"a6"),
   519 => (x"c4",x"87",x"f4",x"ff"),
   520 => (x"d4",x"ff",x"7b",x"c1"),
   521 => (x"79",x"ff",x"c3",x"49"),
   522 => (x"c0",x"1e",x"66",x"d8"),
   523 => (x"d1",x"c1",x"f0",x"ff"),
   524 => (x"02",x"65",x"27",x"1e"),
   525 => (x"c8",x"0f",x"00",x"00"),
   526 => (x"75",x"4d",x"70",x"86"),
   527 => (x"d6",x"c0",x"02",x"9d"),
   528 => (x"dc",x"1e",x"75",x"87"),
   529 => (x"8c",x"27",x"1e",x"66"),
   530 => (x"1e",x"00",x"00",x"08"),
   531 => (x"00",x"00",x"94",x"27"),
   532 => (x"86",x"cc",x"0f",x"00"),
   533 => (x"c8",x"87",x"e8",x"c0"),
   534 => (x"e0",x"c0",x"1e",x"c0"),
   535 => (x"e3",x"fb",x"1e",x"66"),
   536 => (x"70",x"86",x"c8",x"87"),
   537 => (x"72",x"48",x"6b",x"4c"),
   538 => (x"58",x"a6",x"c4",x"98"),
   539 => (x"cc",x"c0",x"02",x"6e"),
   540 => (x"72",x"48",x"6b",x"87"),
   541 => (x"58",x"a6",x"c4",x"98"),
   542 => (x"f4",x"ff",x"05",x"6e"),
   543 => (x"74",x"7b",x"c0",x"87"),
   544 => (x"4d",x"26",x"26",x"48"),
   545 => (x"4b",x"26",x"4c",x"26"),
   546 => (x"4f",x"26",x"4a",x"26"),
   547 => (x"64",x"61",x"65",x"52"),
   548 => (x"6d",x"6f",x"63",x"20"),
   549 => (x"64",x"6e",x"61",x"6d"),
   550 => (x"69",x"61",x"66",x"20"),
   551 => (x"20",x"64",x"65",x"6c"),
   552 => (x"25",x"20",x"74",x"61"),
   553 => (x"25",x"28",x"20",x"64"),
   554 => (x"00",x"0a",x"29",x"64"),
   555 => (x"5b",x"5a",x"5e",x"0e"),
   556 => (x"1e",x"0e",x"5d",x"5c"),
   557 => (x"ff",x"c0",x"1e",x"c0"),
   558 => (x"1e",x"c9",x"c1",x"f0"),
   559 => (x"00",x"02",x"65",x"27"),
   560 => (x"86",x"c8",x"0f",x"00"),
   561 => (x"b8",x"27",x"1e",x"d2"),
   562 => (x"1e",x"00",x"00",x"19"),
   563 => (x"c8",x"87",x"f5",x"f9"),
   564 => (x"c1",x"4d",x"c0",x"86"),
   565 => (x"ad",x"b7",x"d2",x"85"),
   566 => (x"87",x"f7",x"ff",x"04"),
   567 => (x"00",x"19",x"b8",x"27"),
   568 => (x"4a",x"bf",x"97",x"00"),
   569 => (x"c1",x"9a",x"c0",x"c3"),
   570 => (x"05",x"aa",x"b7",x"c0"),
   571 => (x"27",x"87",x"f2",x"c0"),
   572 => (x"00",x"00",x"19",x"bf"),
   573 => (x"d0",x"4a",x"bf",x"97"),
   574 => (x"19",x"c0",x"27",x"32"),
   575 => (x"bf",x"97",x"00",x"00"),
   576 => (x"72",x"33",x"c8",x"4b"),
   577 => (x"27",x"b2",x"73",x"4a"),
   578 => (x"00",x"00",x"19",x"c1"),
   579 => (x"72",x"4b",x"bf",x"97"),
   580 => (x"cf",x"b2",x"73",x"4a"),
   581 => (x"9a",x"ff",x"ff",x"ff"),
   582 => (x"85",x"c1",x"4d",x"72"),
   583 => (x"cb",x"c3",x"35",x"ca"),
   584 => (x"19",x"c1",x"27",x"87"),
   585 => (x"bf",x"97",x"00",x"00"),
   586 => (x"c6",x"32",x"c1",x"4a"),
   587 => (x"19",x"c2",x"27",x"9a"),
   588 => (x"bf",x"97",x"00",x"00"),
   589 => (x"2b",x"b7",x"c7",x"4b"),
   590 => (x"b2",x"73",x"4a",x"72"),
   591 => (x"00",x"19",x"bd",x"27"),
   592 => (x"4b",x"bf",x"97",x"00"),
   593 => (x"98",x"cf",x"48",x"73"),
   594 => (x"27",x"58",x"a6",x"c4"),
   595 => (x"00",x"00",x"19",x"be"),
   596 => (x"c3",x"4b",x"bf",x"97"),
   597 => (x"27",x"33",x"ca",x"9b"),
   598 => (x"00",x"00",x"19",x"bf"),
   599 => (x"c2",x"4c",x"bf",x"97"),
   600 => (x"74",x"4b",x"73",x"34"),
   601 => (x"19",x"c0",x"27",x"b3"),
   602 => (x"bf",x"97",x"00",x"00"),
   603 => (x"9c",x"c0",x"c3",x"4c"),
   604 => (x"73",x"2c",x"b7",x"c6"),
   605 => (x"73",x"b3",x"74",x"4b"),
   606 => (x"1e",x"66",x"c4",x"1e"),
   607 => (x"f9",x"27",x"1e",x"72"),
   608 => (x"1e",x"00",x"00",x"09"),
   609 => (x"00",x"00",x"94",x"27"),
   610 => (x"86",x"d0",x"0f",x"00"),
   611 => (x"48",x"c1",x"82",x"c2"),
   612 => (x"4a",x"70",x"30",x"72"),
   613 => (x"26",x"27",x"1e",x"72"),
   614 => (x"1e",x"00",x"00",x"0a"),
   615 => (x"00",x"00",x"94",x"27"),
   616 => (x"86",x"c8",x"0f",x"00"),
   617 => (x"30",x"6e",x"48",x"c1"),
   618 => (x"c1",x"58",x"a6",x"c4"),
   619 => (x"72",x"4d",x"73",x"83"),
   620 => (x"75",x"1e",x"6e",x"95"),
   621 => (x"0a",x"2f",x"27",x"1e"),
   622 => (x"27",x"1e",x"00",x"00"),
   623 => (x"00",x"00",x"00",x"94"),
   624 => (x"6e",x"86",x"cc",x"0f"),
   625 => (x"b7",x"c0",x"c8",x"49"),
   626 => (x"cf",x"c0",x"06",x"a9"),
   627 => (x"c1",x"4a",x"6e",x"87"),
   628 => (x"2a",x"b7",x"c1",x"35"),
   629 => (x"aa",x"b7",x"c0",x"c8"),
   630 => (x"87",x"f3",x"ff",x"01"),
   631 => (x"45",x"27",x"1e",x"75"),
   632 => (x"1e",x"00",x"00",x"0a"),
   633 => (x"00",x"00",x"94",x"27"),
   634 => (x"86",x"c8",x"0f",x"00"),
   635 => (x"26",x"26",x"48",x"75"),
   636 => (x"26",x"4c",x"26",x"4d"),
   637 => (x"26",x"4a",x"26",x"4b"),
   638 => (x"73",x"5f",x"63",x"4f"),
   639 => (x"5f",x"65",x"7a",x"69"),
   640 => (x"74",x"6c",x"75",x"6d"),
   641 => (x"64",x"25",x"20",x"3a"),
   642 => (x"65",x"72",x"20",x"2c"),
   643 => (x"62",x"5f",x"64",x"61"),
   644 => (x"65",x"6c",x"5f",x"6c"),
   645 => (x"25",x"20",x"3a",x"6e"),
   646 => (x"63",x"20",x"2c",x"64"),
   647 => (x"65",x"7a",x"69",x"73"),
   648 => (x"64",x"25",x"20",x"3a"),
   649 => (x"75",x"4d",x"00",x"0a"),
   650 => (x"25",x"20",x"74",x"6c"),
   651 => (x"25",x"00",x"0a",x"64"),
   652 => (x"6c",x"62",x"20",x"64"),
   653 => (x"73",x"6b",x"63",x"6f"),
   654 => (x"20",x"66",x"6f",x"20"),
   655 => (x"65",x"7a",x"69",x"73"),
   656 => (x"0a",x"64",x"25",x"20"),
   657 => (x"20",x"64",x"25",x"00"),
   658 => (x"63",x"6f",x"6c",x"62"),
   659 => (x"6f",x"20",x"73",x"6b"),
   660 => (x"31",x"35",x"20",x"66"),
   661 => (x"79",x"62",x"20",x"32"),
   662 => (x"0a",x"73",x"65",x"74"),
   663 => (x"5a",x"5e",x"0e",x"00"),
   664 => (x"0e",x"5d",x"5c",x"5b"),
   665 => (x"c0",x"4d",x"66",x"d4"),
   666 => (x"49",x"66",x"dc",x"4c"),
   667 => (x"06",x"a9",x"b7",x"c0"),
   668 => (x"15",x"87",x"fb",x"c0"),
   669 => (x"c0",x"c0",x"c1",x"4b"),
   670 => (x"c4",x"93",x"c0",x"c0"),
   671 => (x"4b",x"93",x"b7",x"c0"),
   672 => (x"bf",x"97",x"66",x"d8"),
   673 => (x"c0",x"c0",x"c1",x"4a"),
   674 => (x"c4",x"92",x"c0",x"c0"),
   675 => (x"4a",x"92",x"b7",x"c0"),
   676 => (x"c1",x"48",x"66",x"d8"),
   677 => (x"58",x"a6",x"dc",x"80"),
   678 => (x"02",x"ab",x"b7",x"72"),
   679 => (x"c1",x"87",x"c5",x"c0"),
   680 => (x"87",x"cc",x"c0",x"48"),
   681 => (x"66",x"dc",x"84",x"c1"),
   682 => (x"ff",x"04",x"ac",x"b7"),
   683 => (x"48",x"c0",x"87",x"c5"),
   684 => (x"4c",x"26",x"4d",x"26"),
   685 => (x"4a",x"26",x"4b",x"26"),
   686 => (x"5e",x"0e",x"4f",x"26"),
   687 => (x"5d",x"5c",x"5b",x"5a"),
   688 => (x"1b",x"d8",x"27",x"0e"),
   689 => (x"c0",x"49",x"00",x"00"),
   690 => (x"18",x"ed",x"27",x"79"),
   691 => (x"27",x"1e",x"00",x"00"),
   692 => (x"00",x"00",x"00",x"5e"),
   693 => (x"27",x"86",x"c4",x"0f"),
   694 => (x"00",x"00",x"19",x"d0"),
   695 => (x"27",x"1e",x"c0",x"1e"),
   696 => (x"00",x"00",x"07",x"f0"),
   697 => (x"70",x"86",x"c8",x"0f"),
   698 => (x"05",x"9a",x"72",x"4a"),
   699 => (x"27",x"87",x"d3",x"c0"),
   700 => (x"00",x"00",x"18",x"19"),
   701 => (x"00",x"5e",x"27",x"1e"),
   702 => (x"c4",x"0f",x"00",x"00"),
   703 => (x"cf",x"48",x"c0",x"86"),
   704 => (x"fa",x"27",x"87",x"d8"),
   705 => (x"1e",x"00",x"00",x"18"),
   706 => (x"00",x"00",x"5e",x"27"),
   707 => (x"86",x"c4",x"0f",x"00"),
   708 => (x"04",x"27",x"4c",x"c0"),
   709 => (x"49",x"00",x"00",x"1c"),
   710 => (x"1e",x"c8",x"79",x"c1"),
   711 => (x"00",x"19",x"11",x"27"),
   712 => (x"06",x"27",x"1e",x"00"),
   713 => (x"1e",x"00",x"00",x"1a"),
   714 => (x"00",x"0a",x"5d",x"27"),
   715 => (x"86",x"cc",x"0f",x"00"),
   716 => (x"9a",x"72",x"4a",x"70"),
   717 => (x"87",x"c8",x"c0",x"05"),
   718 => (x"00",x"1c",x"04",x"27"),
   719 => (x"79",x"c0",x"49",x"00"),
   720 => (x"1a",x"27",x"1e",x"c8"),
   721 => (x"1e",x"00",x"00",x"19"),
   722 => (x"00",x"1a",x"22",x"27"),
   723 => (x"5d",x"27",x"1e",x"00"),
   724 => (x"0f",x"00",x"00",x"0a"),
   725 => (x"4a",x"70",x"86",x"cc"),
   726 => (x"c0",x"05",x"9a",x"72"),
   727 => (x"04",x"27",x"87",x"c8"),
   728 => (x"49",x"00",x"00",x"1c"),
   729 => (x"04",x"27",x"79",x"c0"),
   730 => (x"bf",x"00",x"00",x"1c"),
   731 => (x"19",x"23",x"27",x"1e"),
   732 => (x"27",x"1e",x"00",x"00"),
   733 => (x"00",x"00",x"00",x"94"),
   734 => (x"27",x"86",x"c8",x"0f"),
   735 => (x"00",x"00",x"1c",x"04"),
   736 => (x"c0",x"c3",x"02",x"bf"),
   737 => (x"19",x"d0",x"27",x"87"),
   738 => (x"27",x"4d",x"00",x"00"),
   739 => (x"00",x"00",x"1b",x"8e"),
   740 => (x"1b",x"ce",x"27",x"4b"),
   741 => (x"bf",x"9f",x"00",x"00"),
   742 => (x"27",x"1e",x"72",x"4a"),
   743 => (x"00",x"00",x"1b",x"ce"),
   744 => (x"19",x"d0",x"27",x"4a"),
   745 => (x"72",x"8a",x"00",x"00"),
   746 => (x"c8",x"1e",x"d0",x"1e"),
   747 => (x"4b",x"27",x"1e",x"c0"),
   748 => (x"1e",x"00",x"00",x"18"),
   749 => (x"00",x"00",x"94",x"27"),
   750 => (x"86",x"d4",x"0f",x"00"),
   751 => (x"82",x"c8",x"4a",x"73"),
   752 => (x"ce",x"27",x"4c",x"6a"),
   753 => (x"9f",x"00",x"00",x"1b"),
   754 => (x"d6",x"c5",x"4a",x"bf"),
   755 => (x"05",x"aa",x"b7",x"ea"),
   756 => (x"73",x"87",x"d3",x"c0"),
   757 => (x"6a",x"82",x"c8",x"4a"),
   758 => (x"12",x"45",x"27",x"1e"),
   759 => (x"c4",x"0f",x"00",x"00"),
   760 => (x"c0",x"4c",x"70",x"86"),
   761 => (x"4a",x"75",x"87",x"e4"),
   762 => (x"9f",x"82",x"fe",x"c7"),
   763 => (x"e9",x"ca",x"4a",x"6a"),
   764 => (x"02",x"aa",x"b7",x"d5"),
   765 => (x"27",x"87",x"d3",x"c0"),
   766 => (x"00",x"00",x"18",x"2d"),
   767 => (x"00",x"5e",x"27",x"1e"),
   768 => (x"c4",x"0f",x"00",x"00"),
   769 => (x"cb",x"48",x"c0",x"86"),
   770 => (x"1e",x"74",x"87",x"d0"),
   771 => (x"00",x"18",x"88",x"27"),
   772 => (x"94",x"27",x"1e",x"00"),
   773 => (x"0f",x"00",x"00",x"00"),
   774 => (x"d0",x"27",x"86",x"c8"),
   775 => (x"1e",x"00",x"00",x"19"),
   776 => (x"f0",x"27",x"1e",x"74"),
   777 => (x"0f",x"00",x"00",x"07"),
   778 => (x"4a",x"70",x"86",x"c8"),
   779 => (x"c0",x"05",x"9a",x"72"),
   780 => (x"48",x"c0",x"87",x"c5"),
   781 => (x"27",x"87",x"e3",x"ca"),
   782 => (x"00",x"00",x"18",x"a0"),
   783 => (x"00",x"5e",x"27",x"1e"),
   784 => (x"c4",x"0f",x"00",x"00"),
   785 => (x"19",x"36",x"27",x"86"),
   786 => (x"27",x"1e",x"00",x"00"),
   787 => (x"00",x"00",x"00",x"94"),
   788 => (x"c8",x"86",x"c4",x"0f"),
   789 => (x"19",x"4e",x"27",x"1e"),
   790 => (x"27",x"1e",x"00",x"00"),
   791 => (x"00",x"00",x"1a",x"22"),
   792 => (x"0a",x"5d",x"27",x"1e"),
   793 => (x"cc",x"0f",x"00",x"00"),
   794 => (x"72",x"4a",x"70",x"86"),
   795 => (x"cb",x"c0",x"05",x"9a"),
   796 => (x"1b",x"d8",x"27",x"87"),
   797 => (x"c1",x"49",x"00",x"00"),
   798 => (x"87",x"f1",x"c0",x"79"),
   799 => (x"57",x"27",x"1e",x"c8"),
   800 => (x"1e",x"00",x"00",x"19"),
   801 => (x"00",x"1a",x"06",x"27"),
   802 => (x"5d",x"27",x"1e",x"00"),
   803 => (x"0f",x"00",x"00",x"0a"),
   804 => (x"4a",x"70",x"86",x"cc"),
   805 => (x"c0",x"02",x"9a",x"72"),
   806 => (x"c7",x"27",x"87",x"d3"),
   807 => (x"1e",x"00",x"00",x"18"),
   808 => (x"00",x"00",x"94",x"27"),
   809 => (x"86",x"c4",x"0f",x"00"),
   810 => (x"ed",x"c8",x"48",x"c0"),
   811 => (x"1b",x"ce",x"27",x"87"),
   812 => (x"bf",x"97",x"00",x"00"),
   813 => (x"b7",x"d5",x"c1",x"4a"),
   814 => (x"d0",x"c0",x"05",x"aa"),
   815 => (x"1b",x"cf",x"27",x"87"),
   816 => (x"bf",x"97",x"00",x"00"),
   817 => (x"b7",x"ea",x"c2",x"4a"),
   818 => (x"c5",x"c0",x"02",x"aa"),
   819 => (x"c8",x"48",x"c0",x"87"),
   820 => (x"d0",x"27",x"87",x"c8"),
   821 => (x"97",x"00",x"00",x"19"),
   822 => (x"e9",x"c3",x"4a",x"bf"),
   823 => (x"c0",x"02",x"aa",x"b7"),
   824 => (x"d0",x"27",x"87",x"d5"),
   825 => (x"97",x"00",x"00",x"19"),
   826 => (x"eb",x"c3",x"4a",x"bf"),
   827 => (x"c0",x"02",x"aa",x"b7"),
   828 => (x"48",x"c0",x"87",x"c5"),
   829 => (x"27",x"87",x"e3",x"c7"),
   830 => (x"00",x"00",x"19",x"db"),
   831 => (x"72",x"4a",x"bf",x"97"),
   832 => (x"cf",x"c0",x"05",x"9a"),
   833 => (x"19",x"dc",x"27",x"87"),
   834 => (x"bf",x"97",x"00",x"00"),
   835 => (x"aa",x"b7",x"c2",x"4a"),
   836 => (x"87",x"c5",x"c0",x"02"),
   837 => (x"c1",x"c7",x"48",x"c0"),
   838 => (x"19",x"dd",x"27",x"87"),
   839 => (x"bf",x"97",x"00",x"00"),
   840 => (x"1b",x"d4",x"27",x"48"),
   841 => (x"27",x"58",x"00",x"00"),
   842 => (x"00",x"00",x"1b",x"d0"),
   843 => (x"4b",x"72",x"4a",x"bf"),
   844 => (x"d4",x"27",x"8b",x"c1"),
   845 => (x"49",x"00",x"00",x"1b"),
   846 => (x"1e",x"73",x"79",x"73"),
   847 => (x"60",x"27",x"1e",x"72"),
   848 => (x"1e",x"00",x"00",x"19"),
   849 => (x"00",x"00",x"94",x"27"),
   850 => (x"86",x"cc",x"0f",x"00"),
   851 => (x"00",x"19",x"de",x"27"),
   852 => (x"4a",x"bf",x"97",x"00"),
   853 => (x"df",x"27",x"82",x"74"),
   854 => (x"97",x"00",x"00",x"19"),
   855 => (x"33",x"c8",x"4b",x"bf"),
   856 => (x"80",x"72",x"48",x"73"),
   857 => (x"00",x"1b",x"e8",x"27"),
   858 => (x"e0",x"27",x"58",x"00"),
   859 => (x"97",x"00",x"00",x"19"),
   860 => (x"fc",x"27",x"48",x"bf"),
   861 => (x"58",x"00",x"00",x"1b"),
   862 => (x"00",x"1b",x"d8",x"27"),
   863 => (x"c3",x"02",x"bf",x"00"),
   864 => (x"1e",x"c8",x"87",x"df"),
   865 => (x"00",x"18",x"e4",x"27"),
   866 => (x"22",x"27",x"1e",x"00"),
   867 => (x"1e",x"00",x"00",x"1a"),
   868 => (x"00",x"0a",x"5d",x"27"),
   869 => (x"86",x"cc",x"0f",x"00"),
   870 => (x"9a",x"72",x"4a",x"70"),
   871 => (x"87",x"c5",x"c0",x"02"),
   872 => (x"f5",x"c4",x"48",x"c0"),
   873 => (x"1b",x"d0",x"27",x"87"),
   874 => (x"4b",x"bf",x"00",x"00"),
   875 => (x"30",x"c4",x"48",x"73"),
   876 => (x"00",x"1c",x"00",x"27"),
   877 => (x"f4",x"27",x"58",x"00"),
   878 => (x"49",x"00",x"00",x"1b"),
   879 => (x"f5",x"27",x"79",x"73"),
   880 => (x"97",x"00",x"00",x"19"),
   881 => (x"32",x"c8",x"4a",x"bf"),
   882 => (x"00",x"19",x"f4",x"27"),
   883 => (x"4c",x"bf",x"97",x"00"),
   884 => (x"82",x"74",x"4a",x"72"),
   885 => (x"00",x"19",x"f6",x"27"),
   886 => (x"4c",x"bf",x"97",x"00"),
   887 => (x"4a",x"72",x"34",x"d0"),
   888 => (x"f7",x"27",x"82",x"74"),
   889 => (x"97",x"00",x"00",x"19"),
   890 => (x"34",x"d8",x"4c",x"bf"),
   891 => (x"82",x"74",x"4a",x"72"),
   892 => (x"00",x"1c",x"00",x"27"),
   893 => (x"79",x"72",x"49",x"00"),
   894 => (x"f8",x"27",x"4a",x"72"),
   895 => (x"bf",x"00",x"00",x"1b"),
   896 => (x"27",x"4a",x"72",x"92"),
   897 => (x"00",x"00",x"1b",x"e4"),
   898 => (x"e8",x"27",x"82",x"bf"),
   899 => (x"49",x"00",x"00",x"1b"),
   900 => (x"fd",x"27",x"79",x"72"),
   901 => (x"97",x"00",x"00",x"19"),
   902 => (x"34",x"c8",x"4c",x"bf"),
   903 => (x"00",x"19",x"fc",x"27"),
   904 => (x"4d",x"bf",x"97",x"00"),
   905 => (x"84",x"75",x"4c",x"74"),
   906 => (x"00",x"19",x"fe",x"27"),
   907 => (x"4d",x"bf",x"97",x"00"),
   908 => (x"4c",x"74",x"35",x"d0"),
   909 => (x"ff",x"27",x"84",x"75"),
   910 => (x"97",x"00",x"00",x"19"),
   911 => (x"9d",x"cf",x"4d",x"bf"),
   912 => (x"4c",x"74",x"35",x"d8"),
   913 => (x"ec",x"27",x"84",x"75"),
   914 => (x"49",x"00",x"00",x"1b"),
   915 => (x"8c",x"c2",x"79",x"74"),
   916 => (x"93",x"74",x"4b",x"73"),
   917 => (x"80",x"72",x"48",x"73"),
   918 => (x"00",x"1b",x"f4",x"27"),
   919 => (x"f7",x"c1",x"58",x"00"),
   920 => (x"19",x"e2",x"27",x"87"),
   921 => (x"bf",x"97",x"00",x"00"),
   922 => (x"27",x"32",x"c8",x"4a"),
   923 => (x"00",x"00",x"19",x"e1"),
   924 => (x"72",x"4b",x"bf",x"97"),
   925 => (x"27",x"82",x"73",x"4a"),
   926 => (x"00",x"00",x"1b",x"fc"),
   927 => (x"c5",x"79",x"72",x"49"),
   928 => (x"82",x"ff",x"c7",x"32"),
   929 => (x"f4",x"27",x"2a",x"c9"),
   930 => (x"49",x"00",x"00",x"1b"),
   931 => (x"e7",x"27",x"79",x"72"),
   932 => (x"97",x"00",x"00",x"19"),
   933 => (x"33",x"c8",x"4b",x"bf"),
   934 => (x"00",x"19",x"e6",x"27"),
   935 => (x"4c",x"bf",x"97",x"00"),
   936 => (x"83",x"74",x"4b",x"73"),
   937 => (x"00",x"1c",x"00",x"27"),
   938 => (x"79",x"73",x"49",x"00"),
   939 => (x"f8",x"27",x"4b",x"73"),
   940 => (x"bf",x"00",x"00",x"1b"),
   941 => (x"27",x"4b",x"73",x"93"),
   942 => (x"00",x"00",x"1b",x"e4"),
   943 => (x"f0",x"27",x"83",x"bf"),
   944 => (x"49",x"00",x"00",x"1b"),
   945 => (x"ec",x"27",x"79",x"73"),
   946 => (x"49",x"00",x"00",x"1b"),
   947 => (x"48",x"73",x"79",x"c0"),
   948 => (x"ec",x"27",x"80",x"72"),
   949 => (x"58",x"00",x"00",x"1b"),
   950 => (x"4d",x"26",x"48",x"c1"),
   951 => (x"4b",x"26",x"4c",x"26"),
   952 => (x"4f",x"26",x"4a",x"26"),
   953 => (x"5b",x"5a",x"5e",x"0e"),
   954 => (x"27",x"0e",x"5d",x"5c"),
   955 => (x"00",x"00",x"1b",x"d8"),
   956 => (x"cf",x"c0",x"02",x"bf"),
   957 => (x"4c",x"66",x"d4",x"87"),
   958 => (x"d4",x"2c",x"b7",x"c7"),
   959 => (x"ff",x"c1",x"4b",x"66"),
   960 => (x"87",x"cc",x"c0",x"9b"),
   961 => (x"c8",x"4c",x"66",x"d4"),
   962 => (x"66",x"d4",x"2c",x"b7"),
   963 => (x"9b",x"ff",x"c3",x"4b"),
   964 => (x"00",x"19",x"d0",x"27"),
   965 => (x"e4",x"27",x"1e",x"00"),
   966 => (x"bf",x"00",x"00",x"1b"),
   967 => (x"72",x"82",x"74",x"4a"),
   968 => (x"07",x"f0",x"27",x"1e"),
   969 => (x"c8",x"0f",x"00",x"00"),
   970 => (x"72",x"4a",x"70",x"86"),
   971 => (x"c5",x"c0",x"05",x"9a"),
   972 => (x"c0",x"48",x"c0",x"87"),
   973 => (x"d8",x"27",x"87",x"f2"),
   974 => (x"bf",x"00",x"00",x"1b"),
   975 => (x"87",x"d7",x"c0",x"02"),
   976 => (x"92",x"c4",x"4a",x"73"),
   977 => (x"d0",x"27",x"4a",x"72"),
   978 => (x"82",x"00",x"00",x"19"),
   979 => (x"ff",x"cf",x"4d",x"6a"),
   980 => (x"9d",x"ff",x"ff",x"ff"),
   981 => (x"73",x"87",x"cf",x"c0"),
   982 => (x"72",x"92",x"c2",x"4a"),
   983 => (x"19",x"d0",x"27",x"4a"),
   984 => (x"9f",x"82",x"00",x"00"),
   985 => (x"48",x"75",x"4d",x"6a"),
   986 => (x"4c",x"26",x"4d",x"26"),
   987 => (x"4a",x"26",x"4b",x"26"),
   988 => (x"5e",x"0e",x"4f",x"26"),
   989 => (x"5d",x"5c",x"5b",x"5a"),
   990 => (x"cf",x"8e",x"cc",x"0e"),
   991 => (x"f8",x"ff",x"ff",x"ff"),
   992 => (x"76",x"4c",x"c0",x"4d"),
   993 => (x"1b",x"ec",x"27",x"49"),
   994 => (x"79",x"bf",x"00",x"00"),
   995 => (x"27",x"49",x"a6",x"c4"),
   996 => (x"00",x"00",x"1b",x"f0"),
   997 => (x"d8",x"27",x"79",x"bf"),
   998 => (x"bf",x"00",x"00",x"1b"),
   999 => (x"87",x"cc",x"c0",x"02"),
  1000 => (x"00",x"1b",x"d0",x"27"),
  1001 => (x"c4",x"4a",x"bf",x"00"),
  1002 => (x"87",x"c9",x"c0",x"32"),
  1003 => (x"00",x"1b",x"f4",x"27"),
  1004 => (x"c4",x"4a",x"bf",x"00"),
  1005 => (x"49",x"a6",x"c8",x"32"),
  1006 => (x"4b",x"c0",x"79",x"72"),
  1007 => (x"c0",x"49",x"66",x"c8"),
  1008 => (x"d0",x"c3",x"06",x"a9"),
  1009 => (x"cf",x"4a",x"73",x"87"),
  1010 => (x"05",x"9a",x"72",x"9a"),
  1011 => (x"27",x"87",x"e4",x"c0"),
  1012 => (x"00",x"00",x"19",x"d0"),
  1013 => (x"4a",x"66",x"c8",x"1e"),
  1014 => (x"c1",x"48",x"66",x"c8"),
  1015 => (x"58",x"a6",x"cc",x"80"),
  1016 => (x"f0",x"27",x"1e",x"72"),
  1017 => (x"0f",x"00",x"00",x"07"),
  1018 => (x"d0",x"27",x"86",x"c8"),
  1019 => (x"4c",x"00",x"00",x"19"),
  1020 => (x"c0",x"87",x"c3",x"c0"),
  1021 => (x"6c",x"97",x"84",x"e0"),
  1022 => (x"02",x"9a",x"72",x"4a"),
  1023 => (x"97",x"87",x"cd",x"c2"),
  1024 => (x"e5",x"c3",x"4a",x"6c"),
  1025 => (x"c2",x"02",x"aa",x"b7"),
  1026 => (x"4a",x"74",x"87",x"c2"),
  1027 => (x"6a",x"97",x"82",x"cb"),
  1028 => (x"72",x"9a",x"d8",x"4a"),
  1029 => (x"f3",x"c1",x"05",x"9a"),
  1030 => (x"27",x"1e",x"74",x"87"),
  1031 => (x"00",x"00",x"00",x"5e"),
  1032 => (x"cb",x"86",x"c4",x"0f"),
  1033 => (x"66",x"e8",x"c0",x"1e"),
  1034 => (x"27",x"1e",x"74",x"1e"),
  1035 => (x"00",x"00",x"0a",x"5d"),
  1036 => (x"70",x"86",x"cc",x"0f"),
  1037 => (x"05",x"9a",x"72",x"4a"),
  1038 => (x"74",x"87",x"d1",x"c1"),
  1039 => (x"c0",x"83",x"dc",x"4b"),
  1040 => (x"c4",x"4a",x"66",x"e0"),
  1041 => (x"74",x"7a",x"6b",x"82"),
  1042 => (x"c0",x"83",x"da",x"4b"),
  1043 => (x"c8",x"4a",x"66",x"e0"),
  1044 => (x"48",x"6b",x"9f",x"82"),
  1045 => (x"4d",x"72",x"7a",x"70"),
  1046 => (x"00",x"1b",x"d8",x"27"),
  1047 => (x"c0",x"02",x"bf",x"00"),
  1048 => (x"4a",x"74",x"87",x"d5"),
  1049 => (x"6a",x"9f",x"82",x"d4"),
  1050 => (x"ff",x"ff",x"c0",x"4a"),
  1051 => (x"d0",x"48",x"72",x"9a"),
  1052 => (x"58",x"a6",x"c4",x"30"),
  1053 => (x"76",x"87",x"c4",x"c0"),
  1054 => (x"6e",x"79",x"c0",x"49"),
  1055 => (x"70",x"80",x"6d",x"48"),
  1056 => (x"66",x"e0",x"c0",x"7d"),
  1057 => (x"c1",x"79",x"c0",x"49"),
  1058 => (x"87",x"ce",x"c1",x"48"),
  1059 => (x"66",x"c8",x"83",x"c1"),
  1060 => (x"f0",x"fc",x"04",x"ab"),
  1061 => (x"ff",x"ff",x"cf",x"87"),
  1062 => (x"27",x"4d",x"f8",x"ff"),
  1063 => (x"00",x"00",x"1b",x"d8"),
  1064 => (x"f3",x"c0",x"02",x"bf"),
  1065 => (x"27",x"1e",x"6e",x"87"),
  1066 => (x"00",x"00",x"0e",x"e4"),
  1067 => (x"c4",x"86",x"c4",x"0f"),
  1068 => (x"4a",x"6e",x"58",x"a6"),
  1069 => (x"aa",x"75",x"9a",x"75"),
  1070 => (x"87",x"dc",x"c0",x"02"),
  1071 => (x"8a",x"c2",x"4a",x"6e"),
  1072 => (x"d0",x"27",x"4a",x"72"),
  1073 => (x"bf",x"00",x"00",x"1b"),
  1074 => (x"1b",x"e8",x"27",x"92"),
  1075 => (x"48",x"bf",x"00",x"00"),
  1076 => (x"a6",x"c8",x"80",x"72"),
  1077 => (x"87",x"e2",x"fb",x"58"),
  1078 => (x"ff",x"cf",x"48",x"c0"),
  1079 => (x"4d",x"f8",x"ff",x"ff"),
  1080 => (x"4d",x"26",x"86",x"cc"),
  1081 => (x"4b",x"26",x"4c",x"26"),
  1082 => (x"4f",x"26",x"4a",x"26"),
  1083 => (x"5b",x"5a",x"5e",x"0e"),
  1084 => (x"bf",x"66",x"cc",x"0e"),
  1085 => (x"cc",x"82",x"c1",x"4a"),
  1086 => (x"79",x"72",x"49",x"66"),
  1087 => (x"d4",x"27",x"4a",x"72"),
  1088 => (x"bf",x"00",x"00",x"1b"),
  1089 => (x"05",x"9a",x"72",x"9a"),
  1090 => (x"cc",x"87",x"d3",x"c0"),
  1091 => (x"82",x"c8",x"4a",x"66"),
  1092 => (x"e4",x"27",x"1e",x"6a"),
  1093 => (x"0f",x"00",x"00",x"0e"),
  1094 => (x"4b",x"70",x"86",x"c4"),
  1095 => (x"48",x"c1",x"7a",x"73"),
  1096 => (x"4a",x"26",x"4b",x"26"),
  1097 => (x"5e",x"0e",x"4f",x"26"),
  1098 => (x"27",x"0e",x"5b",x"5a"),
  1099 => (x"00",x"00",x"1b",x"e8"),
  1100 => (x"66",x"cc",x"4a",x"bf"),
  1101 => (x"6b",x"83",x"c8",x"4b"),
  1102 => (x"73",x"8b",x"c2",x"4b"),
  1103 => (x"1b",x"d0",x"27",x"4b"),
  1104 => (x"93",x"bf",x"00",x"00"),
  1105 => (x"82",x"73",x"4a",x"72"),
  1106 => (x"00",x"1b",x"d4",x"27"),
  1107 => (x"cc",x"4b",x"bf",x"00"),
  1108 => (x"72",x"9b",x"bf",x"66"),
  1109 => (x"d0",x"82",x"73",x"4a"),
  1110 => (x"1e",x"72",x"1e",x"66"),
  1111 => (x"00",x"07",x"f0",x"27"),
  1112 => (x"86",x"c8",x"0f",x"00"),
  1113 => (x"9a",x"72",x"4a",x"70"),
  1114 => (x"87",x"c5",x"c0",x"05"),
  1115 => (x"c2",x"c0",x"48",x"c0"),
  1116 => (x"26",x"48",x"c1",x"87"),
  1117 => (x"26",x"4a",x"26",x"4b"),
  1118 => (x"5a",x"5e",x"0e",x"4f"),
  1119 => (x"0e",x"5d",x"5c",x"5b"),
  1120 => (x"d4",x"4c",x"66",x"d8"),
  1121 => (x"08",x"27",x"1e",x"66"),
  1122 => (x"1e",x"00",x"00",x"1c"),
  1123 => (x"00",x"0f",x"72",x"27"),
  1124 => (x"86",x"c8",x"0f",x"00"),
  1125 => (x"9a",x"72",x"4a",x"70"),
  1126 => (x"87",x"df",x"c1",x"02"),
  1127 => (x"00",x"1c",x"0c",x"27"),
  1128 => (x"c7",x"4a",x"bf",x"00"),
  1129 => (x"2a",x"c9",x"82",x"ff"),
  1130 => (x"4b",x"c0",x"4d",x"72"),
  1131 => (x"00",x"12",x"1d",x"27"),
  1132 => (x"5e",x"27",x"1e",x"00"),
  1133 => (x"0f",x"00",x"00",x"00"),
  1134 => (x"b7",x"c0",x"86",x"c4"),
  1135 => (x"d0",x"c1",x"06",x"ad"),
  1136 => (x"27",x"1e",x"74",x"87"),
  1137 => (x"00",x"00",x"1c",x"08"),
  1138 => (x"11",x"26",x"27",x"1e"),
  1139 => (x"c8",x"0f",x"00",x"00"),
  1140 => (x"72",x"4a",x"70",x"86"),
  1141 => (x"c5",x"c0",x"05",x"9a"),
  1142 => (x"c0",x"48",x"c0",x"87"),
  1143 => (x"08",x"27",x"87",x"f5"),
  1144 => (x"1e",x"00",x"00",x"1c"),
  1145 => (x"00",x"10",x"ec",x"27"),
  1146 => (x"86",x"c4",x"0f",x"00"),
  1147 => (x"c1",x"84",x"c0",x"c8"),
  1148 => (x"ab",x"b7",x"75",x"83"),
  1149 => (x"87",x"c9",x"ff",x"04"),
  1150 => (x"d4",x"87",x"d6",x"c0"),
  1151 => (x"36",x"27",x"1e",x"66"),
  1152 => (x"1e",x"00",x"00",x"12"),
  1153 => (x"00",x"00",x"94",x"27"),
  1154 => (x"86",x"c8",x"0f",x"00"),
  1155 => (x"c2",x"c0",x"48",x"c0"),
  1156 => (x"26",x"48",x"c1",x"87"),
  1157 => (x"26",x"4c",x"26",x"4d"),
  1158 => (x"26",x"4a",x"26",x"4b"),
  1159 => (x"65",x"70",x"4f",x"4f"),
  1160 => (x"20",x"64",x"65",x"6e"),
  1161 => (x"65",x"6c",x"69",x"66"),
  1162 => (x"6f",x"6c",x"20",x"2c"),
  1163 => (x"6e",x"69",x"64",x"61"),
  1164 => (x"2e",x"2e",x"2e",x"67"),
  1165 => (x"61",x"43",x"00",x"0a"),
  1166 => (x"20",x"74",x"27",x"6e"),
  1167 => (x"6e",x"65",x"70",x"6f"),
  1168 => (x"0a",x"73",x"25",x"20"),
  1169 => (x"5a",x"5e",x"0e",x"00"),
  1170 => (x"66",x"cc",x"0e",x"5b"),
  1171 => (x"c3",x"2a",x"d8",x"4a"),
  1172 => (x"66",x"cc",x"9a",x"ff"),
  1173 => (x"cf",x"2b",x"c8",x"4b"),
  1174 => (x"72",x"9b",x"c0",x"fc"),
  1175 => (x"cc",x"b2",x"73",x"4a"),
  1176 => (x"33",x"c8",x"4b",x"66"),
  1177 => (x"c0",x"f0",x"ff",x"c0"),
  1178 => (x"4a",x"72",x"9b",x"c0"),
  1179 => (x"66",x"cc",x"b2",x"73"),
  1180 => (x"ff",x"33",x"d8",x"4b"),
  1181 => (x"c0",x"c0",x"c0",x"c0"),
  1182 => (x"73",x"4a",x"72",x"9b"),
  1183 => (x"26",x"48",x"72",x"b2"),
  1184 => (x"26",x"4a",x"26",x"4b"),
  1185 => (x"5a",x"5e",x"0e",x"4f"),
  1186 => (x"66",x"cc",x"0e",x"5b"),
  1187 => (x"c3",x"2b",x"c8",x"4b"),
  1188 => (x"cc",x"4b",x"9b",x"ff"),
  1189 => (x"32",x"c8",x"4a",x"66"),
  1190 => (x"9a",x"c0",x"fc",x"cf"),
  1191 => (x"b2",x"73",x"4a",x"72"),
  1192 => (x"26",x"48",x"72",x"4a"),
  1193 => (x"26",x"4a",x"26",x"4b"),
  1194 => (x"5a",x"5e",x"0e",x"4f"),
  1195 => (x"66",x"cc",x"0e",x"5b"),
  1196 => (x"cf",x"2a",x"d0",x"4a"),
  1197 => (x"4a",x"9a",x"ff",x"ff"),
  1198 => (x"d0",x"4b",x"66",x"cc"),
  1199 => (x"c0",x"c0",x"f0",x"33"),
  1200 => (x"73",x"4a",x"72",x"9b"),
  1201 => (x"26",x"48",x"72",x"b2"),
  1202 => (x"26",x"4a",x"26",x"4b"),
  1203 => (x"1e",x"72",x"1e",x"4f"),
  1204 => (x"c0",x"c0",x"c0",x"d0"),
  1205 => (x"0f",x"72",x"4a",x"c0"),
  1206 => (x"26",x"87",x"fd",x"ff"),
  1207 => (x"1e",x"4f",x"26",x"4a"),
  1208 => (x"66",x"cc",x"1e",x"72"),
  1209 => (x"9a",x"df",x"c3",x"4a"),
  1210 => (x"c0",x"8a",x"f7",x"c0"),
  1211 => (x"c0",x"03",x"aa",x"b7"),
  1212 => (x"e7",x"c0",x"87",x"c3"),
  1213 => (x"48",x"66",x"c8",x"82"),
  1214 => (x"a6",x"cc",x"30",x"c4"),
  1215 => (x"48",x"66",x"c8",x"58"),
  1216 => (x"a6",x"cc",x"b0",x"72"),
  1217 => (x"48",x"66",x"c8",x"58"),
  1218 => (x"4f",x"26",x"4a",x"26"),
  1219 => (x"5b",x"5a",x"5e",x"0e"),
  1220 => (x"d0",x"0e",x"5d",x"5c"),
  1221 => (x"c0",x"c0",x"c0",x"c0"),
  1222 => (x"1c",x"18",x"27",x"4d"),
  1223 => (x"48",x"bf",x"00",x"00"),
  1224 => (x"1c",x"27",x"80",x"c1"),
  1225 => (x"58",x"00",x"00",x"1c"),
  1226 => (x"4a",x"66",x"d4",x"97"),
  1227 => (x"c0",x"c0",x"c0",x"c1"),
  1228 => (x"c0",x"c4",x"92",x"c0"),
  1229 => (x"c1",x"4a",x"92",x"b7"),
  1230 => (x"05",x"aa",x"b7",x"d3"),
  1231 => (x"27",x"87",x"e9",x"c0"),
  1232 => (x"00",x"00",x"1c",x"18"),
  1233 => (x"27",x"79",x"c0",x"49"),
  1234 => (x"00",x"00",x"1c",x"1c"),
  1235 => (x"27",x"79",x"c0",x"49"),
  1236 => (x"00",x"00",x"1c",x"24"),
  1237 => (x"27",x"79",x"c0",x"49"),
  1238 => (x"00",x"00",x"1c",x"28"),
  1239 => (x"ff",x"79",x"c0",x"49"),
  1240 => (x"d3",x"c1",x"49",x"c0"),
  1241 => (x"87",x"cb",x"ca",x"79"),
  1242 => (x"00",x"1c",x"18",x"27"),
  1243 => (x"c1",x"49",x"bf",x"00"),
  1244 => (x"c1",x"05",x"a9",x"b7"),
  1245 => (x"c0",x"ff",x"87",x"db"),
  1246 => (x"79",x"f4",x"c1",x"49"),
  1247 => (x"4a",x"66",x"d4",x"97"),
  1248 => (x"c0",x"c0",x"c0",x"c1"),
  1249 => (x"c0",x"c4",x"92",x"c0"),
  1250 => (x"72",x"4a",x"92",x"b7"),
  1251 => (x"1c",x"28",x"27",x"1e"),
  1252 => (x"1e",x"bf",x"00",x"00"),
  1253 => (x"00",x"12",x"df",x"27"),
  1254 => (x"86",x"c8",x"0f",x"00"),
  1255 => (x"00",x"1c",x"2c",x"27"),
  1256 => (x"28",x"27",x"58",x"00"),
  1257 => (x"bf",x"00",x"00",x"1c"),
  1258 => (x"ac",x"b7",x"c3",x"4c"),
  1259 => (x"87",x"c6",x"c0",x"06"),
  1260 => (x"88",x"74",x"48",x"ca"),
  1261 => (x"4a",x"74",x"4c",x"70"),
  1262 => (x"48",x"72",x"82",x"c1"),
  1263 => (x"24",x"27",x"30",x"c1"),
  1264 => (x"58",x"00",x"00",x"1c"),
  1265 => (x"f0",x"c0",x"48",x"74"),
  1266 => (x"49",x"c0",x"ff",x"80"),
  1267 => (x"e2",x"c8",x"79",x"70"),
  1268 => (x"1c",x"28",x"27",x"87"),
  1269 => (x"49",x"bf",x"00",x"00"),
  1270 => (x"01",x"a9",x"b7",x"c9"),
  1271 => (x"27",x"87",x"d4",x"c8"),
  1272 => (x"00",x"00",x"1c",x"28"),
  1273 => (x"b7",x"c0",x"49",x"bf"),
  1274 => (x"c6",x"c8",x"06",x"a9"),
  1275 => (x"1c",x"28",x"27",x"87"),
  1276 => (x"48",x"bf",x"00",x"00"),
  1277 => (x"ff",x"80",x"f0",x"c0"),
  1278 => (x"79",x"70",x"49",x"c0"),
  1279 => (x"00",x"1c",x"18",x"27"),
  1280 => (x"c3",x"49",x"bf",x"00"),
  1281 => (x"c0",x"01",x"a9",x"b7"),
  1282 => (x"d4",x"97",x"87",x"e9"),
  1283 => (x"c0",x"c1",x"4a",x"66"),
  1284 => (x"92",x"c0",x"c0",x"c0"),
  1285 => (x"92",x"b7",x"c0",x"c4"),
  1286 => (x"27",x"1e",x"72",x"4a"),
  1287 => (x"00",x"00",x"1c",x"24"),
  1288 => (x"df",x"27",x"1e",x"bf"),
  1289 => (x"0f",x"00",x"00",x"12"),
  1290 => (x"28",x"27",x"86",x"c8"),
  1291 => (x"58",x"00",x"00",x"1c"),
  1292 => (x"27",x"87",x"c0",x"c7"),
  1293 => (x"00",x"00",x"1c",x"20"),
  1294 => (x"82",x"c3",x"4a",x"bf"),
  1295 => (x"00",x"1c",x"18",x"27"),
  1296 => (x"72",x"49",x"bf",x"00"),
  1297 => (x"c0",x"01",x"a9",x"b7"),
  1298 => (x"d4",x"97",x"87",x"f1"),
  1299 => (x"c0",x"c1",x"4a",x"66"),
  1300 => (x"92",x"c0",x"c0",x"c0"),
  1301 => (x"92",x"b7",x"c0",x"c4"),
  1302 => (x"27",x"1e",x"72",x"4a"),
  1303 => (x"00",x"00",x"1c",x"1c"),
  1304 => (x"df",x"27",x"1e",x"bf"),
  1305 => (x"0f",x"00",x"00",x"12"),
  1306 => (x"20",x"27",x"86",x"c8"),
  1307 => (x"58",x"00",x"00",x"1c"),
  1308 => (x"00",x"1c",x"2c",x"27"),
  1309 => (x"79",x"c1",x"49",x"00"),
  1310 => (x"27",x"87",x"f8",x"c5"),
  1311 => (x"00",x"00",x"1c",x"28"),
  1312 => (x"b7",x"c0",x"49",x"bf"),
  1313 => (x"d0",x"c3",x"06",x"a9"),
  1314 => (x"1c",x"28",x"27",x"87"),
  1315 => (x"49",x"bf",x"00",x"00"),
  1316 => (x"01",x"a9",x"b7",x"c3"),
  1317 => (x"27",x"87",x"c2",x"c3"),
  1318 => (x"00",x"00",x"1c",x"24"),
  1319 => (x"32",x"c1",x"4a",x"bf"),
  1320 => (x"18",x"27",x"82",x"c1"),
  1321 => (x"bf",x"00",x"00",x"1c"),
  1322 => (x"a9",x"b7",x"72",x"49"),
  1323 => (x"87",x"c2",x"c2",x"01"),
  1324 => (x"4a",x"66",x"d4",x"97"),
  1325 => (x"c0",x"c0",x"c0",x"c1"),
  1326 => (x"c0",x"c4",x"92",x"c0"),
  1327 => (x"72",x"4a",x"92",x"b7"),
  1328 => (x"1c",x"30",x"27",x"1e"),
  1329 => (x"1e",x"bf",x"00",x"00"),
  1330 => (x"00",x"12",x"df",x"27"),
  1331 => (x"86",x"c8",x"0f",x"00"),
  1332 => (x"00",x"1c",x"34",x"27"),
  1333 => (x"2c",x"27",x"58",x"00"),
  1334 => (x"bf",x"00",x"00",x"1c"),
  1335 => (x"27",x"8a",x"c1",x"4a"),
  1336 => (x"00",x"00",x"1c",x"2c"),
  1337 => (x"c0",x"79",x"72",x"49"),
  1338 => (x"c4",x"03",x"aa",x"b7"),
  1339 => (x"1c",x"27",x"87",x"c5"),
  1340 => (x"bf",x"00",x"00",x"1c"),
  1341 => (x"1c",x"30",x"27",x"4a"),
  1342 => (x"bf",x"97",x"00",x"00"),
  1343 => (x"1c",x"1c",x"27",x"52"),
  1344 => (x"4a",x"bf",x"00",x"00"),
  1345 => (x"1c",x"27",x"82",x"c1"),
  1346 => (x"49",x"00",x"00",x"1c"),
  1347 => (x"34",x"27",x"79",x"72"),
  1348 => (x"bf",x"00",x"00",x"1c"),
  1349 => (x"c0",x"06",x"aa",x"b7"),
  1350 => (x"34",x"27",x"87",x"cd"),
  1351 => (x"49",x"00",x"00",x"1c"),
  1352 => (x"00",x"1c",x"1c",x"27"),
  1353 => (x"27",x"79",x"bf",x"00"),
  1354 => (x"00",x"00",x"1c",x"2c"),
  1355 => (x"c3",x"79",x"c1",x"49"),
  1356 => (x"2c",x"27",x"87",x"c1"),
  1357 => (x"bf",x"00",x"00",x"1c"),
  1358 => (x"87",x"f7",x"c2",x"05"),
  1359 => (x"00",x"1c",x"30",x"27"),
  1360 => (x"c4",x"4b",x"bf",x"00"),
  1361 => (x"1c",x"30",x"27",x"33"),
  1362 => (x"73",x"49",x"00",x"00"),
  1363 => (x"1c",x"1c",x"27",x"79"),
  1364 => (x"4a",x"bf",x"00",x"00"),
  1365 => (x"da",x"c2",x"52",x"73"),
  1366 => (x"1c",x"28",x"27",x"87"),
  1367 => (x"49",x"bf",x"00",x"00"),
  1368 => (x"04",x"a9",x"b7",x"c7"),
  1369 => (x"c0",x"87",x"fd",x"c1"),
  1370 => (x"49",x"f4",x"fe",x"4b"),
  1371 => (x"34",x"27",x"79",x"c1"),
  1372 => (x"bf",x"00",x"00",x"1c"),
  1373 => (x"27",x"1e",x"75",x"1e"),
  1374 => (x"00",x"00",x"19",x"84"),
  1375 => (x"00",x"94",x"27",x"1e"),
  1376 => (x"cc",x"0f",x"00",x"00"),
  1377 => (x"1c",x"1c",x"27",x"86"),
  1378 => (x"75",x"49",x"00",x"00"),
  1379 => (x"1c",x"1c",x"27",x"79"),
  1380 => (x"49",x"bf",x"00",x"00"),
  1381 => (x"00",x"1c",x"34",x"27"),
  1382 => (x"a9",x"b7",x"bf",x"00"),
  1383 => (x"87",x"e5",x"c0",x"03"),
  1384 => (x"00",x"1c",x"1c",x"27"),
  1385 => (x"83",x"bf",x"bf",x"00"),
  1386 => (x"00",x"1c",x"1c",x"27"),
  1387 => (x"c4",x"4a",x"bf",x"00"),
  1388 => (x"1c",x"1c",x"27",x"82"),
  1389 => (x"72",x"49",x"00",x"00"),
  1390 => (x"1c",x"34",x"27",x"79"),
  1391 => (x"b7",x"bf",x"00",x"00"),
  1392 => (x"db",x"ff",x"04",x"aa"),
  1393 => (x"27",x"1e",x"73",x"87"),
  1394 => (x"00",x"00",x"19",x"a3"),
  1395 => (x"00",x"94",x"27",x"1e"),
  1396 => (x"c8",x"0f",x"00",x"00"),
  1397 => (x"49",x"c0",x"ff",x"86"),
  1398 => (x"27",x"79",x"c2",x"c1"),
  1399 => (x"00",x"00",x"12",x"cd"),
  1400 => (x"87",x"cf",x"c0",x"0f"),
  1401 => (x"00",x"1c",x"28",x"27"),
  1402 => (x"c0",x"48",x"bf",x"00"),
  1403 => (x"c0",x"ff",x"80",x"f0"),
  1404 => (x"26",x"79",x"70",x"49"),
  1405 => (x"26",x"4c",x"26",x"4d"),
  1406 => (x"26",x"4a",x"26",x"4b"),
  1407 => (x"fd",x"ff",x"1e",x"4f"),
  1408 => (x"0e",x"4f",x"26",x"87"),
  1409 => (x"5c",x"5b",x"5a",x"5e"),
  1410 => (x"eb",x"27",x"0e",x"5d"),
  1411 => (x"1e",x"00",x"00",x"17"),
  1412 => (x"00",x"00",x"5e",x"27"),
  1413 => (x"86",x"c4",x"0f",x"00"),
  1414 => (x"00",x"04",x"f9",x"27"),
  1415 => (x"4a",x"70",x"0f",x"00"),
  1416 => (x"c4",x"02",x"9a",x"72"),
  1417 => (x"c8",x"27",x"87",x"ce"),
  1418 => (x"1e",x"00",x"00",x"17"),
  1419 => (x"00",x"00",x"5e",x"27"),
  1420 => (x"86",x"c4",x"0f",x"00"),
  1421 => (x"00",x"0a",x"ba",x"27"),
  1422 => (x"38",x"27",x"0f",x"00"),
  1423 => (x"1e",x"00",x"00",x"1c"),
  1424 => (x"00",x"17",x"df",x"27"),
  1425 => (x"79",x"27",x"1e",x"00"),
  1426 => (x"0f",x"00",x"00",x"11"),
  1427 => (x"4a",x"70",x"86",x"c8"),
  1428 => (x"c3",x"02",x"9a",x"72"),
  1429 => (x"38",x"27",x"87",x"d0"),
  1430 => (x"4b",x"00",x"00",x"1c"),
  1431 => (x"00",x"17",x"9d",x"27"),
  1432 => (x"5e",x"27",x"1e",x"00"),
  1433 => (x"0f",x"00",x"00",x"00"),
  1434 => (x"4d",x"c0",x"86",x"c4"),
  1435 => (x"4a",x"74",x"4c",x"13"),
  1436 => (x"aa",x"b7",x"e0",x"c0"),
  1437 => (x"87",x"ed",x"c1",x"02"),
  1438 => (x"c0",x"ff",x"48",x"74"),
  1439 => (x"74",x"79",x"70",x"49"),
  1440 => (x"b7",x"e3",x"c0",x"4a"),
  1441 => (x"dc",x"c1",x"02",x"aa"),
  1442 => (x"c1",x"4a",x"74",x"87"),
  1443 => (x"05",x"aa",x"b7",x"c7"),
  1444 => (x"27",x"87",x"c6",x"c0"),
  1445 => (x"00",x"00",x"12",x"cd"),
  1446 => (x"ca",x"4a",x"74",x"0f"),
  1447 => (x"c0",x"05",x"aa",x"b7"),
  1448 => (x"fd",x"27",x"87",x"c6"),
  1449 => (x"0f",x"00",x"00",x"15"),
  1450 => (x"cc",x"c1",x"4a",x"74"),
  1451 => (x"c0",x"05",x"aa",x"b7"),
  1452 => (x"38",x"27",x"87",x"c6"),
  1453 => (x"4b",x"00",x"00",x"1c"),
  1454 => (x"df",x"ff",x"4a",x"74"),
  1455 => (x"72",x"8a",x"d0",x"9a"),
  1456 => (x"c0",x"4a",x"74",x"4c"),
  1457 => (x"04",x"aa",x"b7",x"f9"),
  1458 => (x"74",x"87",x"c6",x"c0"),
  1459 => (x"72",x"8a",x"d1",x"4a"),
  1460 => (x"74",x"35",x"c4",x"4c"),
  1461 => (x"72",x"4d",x"75",x"4a"),
  1462 => (x"74",x"4c",x"13",x"b5"),
  1463 => (x"b7",x"e0",x"c0",x"4a"),
  1464 => (x"d3",x"fe",x"05",x"aa"),
  1465 => (x"c0",x"4a",x"74",x"87"),
  1466 => (x"02",x"aa",x"b7",x"e3"),
  1467 => (x"13",x"87",x"e2",x"c0"),
  1468 => (x"b7",x"e0",x"c0",x"4a"),
  1469 => (x"ca",x"c0",x"05",x"aa"),
  1470 => (x"c0",x"4a",x"13",x"87"),
  1471 => (x"02",x"aa",x"b7",x"e0"),
  1472 => (x"c1",x"87",x"f6",x"ff"),
  1473 => (x"73",x"1e",x"75",x"8b"),
  1474 => (x"11",x"79",x"27",x"1e"),
  1475 => (x"c8",x"0f",x"00",x"00"),
  1476 => (x"ca",x"4a",x"13",x"86"),
  1477 => (x"fd",x"02",x"aa",x"b7"),
  1478 => (x"4a",x"13",x"87",x"d0"),
  1479 => (x"05",x"aa",x"b7",x"ca"),
  1480 => (x"fd",x"87",x"f7",x"ff"),
  1481 => (x"af",x"27",x"87",x"c4"),
  1482 => (x"1e",x"00",x"00",x"17"),
  1483 => (x"00",x"00",x"5e",x"27"),
  1484 => (x"86",x"c4",x"0f",x"00"),
  1485 => (x"00",x"18",x"01",x"27"),
  1486 => (x"5e",x"27",x"1e",x"00"),
  1487 => (x"0f",x"00",x"00",x"00"),
  1488 => (x"34",x"27",x"86",x"c4"),
  1489 => (x"49",x"00",x"00",x"1c"),
  1490 => (x"f4",x"c3",x"79",x"c0"),
  1491 => (x"c0",x"4d",x"ff",x"c8"),
  1492 => (x"3f",x"27",x"1e",x"ee"),
  1493 => (x"0f",x"00",x"00",x"00"),
  1494 => (x"4b",x"75",x"86",x"c4"),
  1495 => (x"c0",x"c9",x"f4",x"c3"),
  1496 => (x"bf",x"c0",x"ff",x"4d"),
  1497 => (x"c8",x"4a",x"74",x"4c"),
  1498 => (x"9a",x"72",x"9a",x"c0"),
  1499 => (x"87",x"d1",x"c0",x"02"),
  1500 => (x"ff",x"c3",x"4a",x"74"),
  1501 => (x"27",x"1e",x"72",x"9a"),
  1502 => (x"00",x"00",x"13",x"0c"),
  1503 => (x"75",x"86",x"c4",x"0f"),
  1504 => (x"c1",x"4a",x"73",x"4b"),
  1505 => (x"05",x"9a",x"72",x"8b"),
  1506 => (x"c3",x"87",x"d6",x"ff"),
  1507 => (x"4d",x"ff",x"c8",x"f4"),
  1508 => (x"26",x"87",x"fc",x"fe"),
  1509 => (x"26",x"4c",x"26",x"4d"),
  1510 => (x"26",x"4a",x"26",x"4b"),
  1511 => (x"72",x"61",x"50",x"4f"),
  1512 => (x"67",x"6e",x"69",x"73"),
  1513 => (x"6e",x"61",x"6d",x"20"),
  1514 => (x"73",x"65",x"66",x"69"),
  1515 => (x"4c",x"00",x"0a",x"74"),
  1516 => (x"69",x"64",x"61",x"6f"),
  1517 => (x"6d",x"20",x"67",x"6e"),
  1518 => (x"66",x"69",x"6e",x"61"),
  1519 => (x"20",x"74",x"73",x"65"),
  1520 => (x"6c",x"69",x"61",x"66"),
  1521 => (x"00",x"0a",x"64",x"65"),
  1522 => (x"74",x"6e",x"75",x"48"),
  1523 => (x"20",x"67",x"6e",x"69"),
  1524 => (x"20",x"72",x"6f",x"66"),
  1525 => (x"74",x"72",x"61",x"70"),
  1526 => (x"6f",x"69",x"74",x"69"),
  1527 => (x"4d",x"00",x"0a",x"6e"),
  1528 => (x"46",x"49",x"4e",x"41"),
  1529 => (x"4d",x"54",x"53",x"45"),
  1530 => (x"49",x"00",x"54",x"53"),
  1531 => (x"69",x"74",x"69",x"6e"),
  1532 => (x"7a",x"69",x"6c",x"61"),
  1533 => (x"20",x"67",x"6e",x"69"),
  1534 => (x"63",x"20",x"44",x"53"),
  1535 => (x"0a",x"64",x"72",x"61"),
  1536 => (x"6f",x"6f",x"42",x"00"),
  1537 => (x"67",x"6e",x"69",x"74"),
  1538 => (x"6f",x"72",x"66",x"20"),
  1539 => (x"53",x"52",x"20",x"6d"),
  1540 => (x"2e",x"32",x"33",x"32"),
  1541 => (x"44",x"4d",x"43",x"00"),
  1542 => (x"61",x"65",x"52",x"00"),
  1543 => (x"66",x"6f",x"20",x"64"),
  1544 => (x"52",x"42",x"4d",x"20"),
  1545 => (x"69",x"61",x"66",x"20"),
  1546 => (x"0a",x"64",x"65",x"6c"),
  1547 => (x"20",x"6f",x"4e",x"00"),
  1548 => (x"74",x"72",x"61",x"70"),
  1549 => (x"6f",x"69",x"74",x"69"),
  1550 => (x"69",x"73",x"20",x"6e"),
  1551 => (x"74",x"61",x"6e",x"67"),
  1552 => (x"20",x"65",x"72",x"75"),
  1553 => (x"6e",x"75",x"6f",x"66"),
  1554 => (x"4d",x"00",x"0a",x"64"),
  1555 => (x"69",x"73",x"52",x"42"),
  1556 => (x"20",x"3a",x"65",x"7a"),
  1557 => (x"20",x"2c",x"64",x"25"),
  1558 => (x"74",x"72",x"61",x"70"),
  1559 => (x"6f",x"69",x"74",x"69"),
  1560 => (x"7a",x"69",x"73",x"6e"),
  1561 => (x"25",x"20",x"3a",x"65"),
  1562 => (x"6f",x"20",x"2c",x"64"),
  1563 => (x"65",x"73",x"66",x"66"),
  1564 => (x"66",x"6f",x"20",x"74"),
  1565 => (x"67",x"69",x"73",x"20"),
  1566 => (x"64",x"25",x"20",x"3a"),
  1567 => (x"69",x"73",x"20",x"2c"),
  1568 => (x"78",x"30",x"20",x"67"),
  1569 => (x"00",x"0a",x"78",x"25"),
  1570 => (x"64",x"61",x"65",x"52"),
  1571 => (x"20",x"67",x"6e",x"69"),
  1572 => (x"74",x"6f",x"6f",x"62"),
  1573 => (x"63",x"65",x"73",x"20"),
  1574 => (x"20",x"72",x"6f",x"74"),
  1575 => (x"00",x"0a",x"64",x"25"),
  1576 => (x"64",x"61",x"65",x"52"),
  1577 => (x"6f",x"6f",x"62",x"20"),
  1578 => (x"65",x"73",x"20",x"74"),
  1579 => (x"72",x"6f",x"74",x"63"),
  1580 => (x"6f",x"72",x"66",x"20"),
  1581 => (x"69",x"66",x"20",x"6d"),
  1582 => (x"20",x"74",x"73",x"72"),
  1583 => (x"74",x"72",x"61",x"70"),
  1584 => (x"6f",x"69",x"74",x"69"),
  1585 => (x"55",x"00",x"0a",x"6e"),
  1586 => (x"70",x"75",x"73",x"6e"),
  1587 => (x"74",x"72",x"6f",x"70"),
  1588 => (x"70",x"20",x"64",x"65"),
  1589 => (x"69",x"74",x"72",x"61"),
  1590 => (x"6e",x"6f",x"69",x"74"),
  1591 => (x"70",x"79",x"74",x"20"),
  1592 => (x"00",x"0d",x"21",x"65"),
  1593 => (x"33",x"54",x"41",x"46"),
  1594 => (x"20",x"20",x"20",x"32"),
  1595 => (x"61",x"65",x"52",x"00"),
  1596 => (x"67",x"6e",x"69",x"64"),
  1597 => (x"52",x"42",x"4d",x"20"),
  1598 => (x"42",x"4d",x"00",x"0a"),
  1599 => (x"75",x"73",x"20",x"52"),
  1600 => (x"73",x"65",x"63",x"63"),
  1601 => (x"6c",x"75",x"66",x"73"),
  1602 => (x"72",x"20",x"79",x"6c"),
  1603 => (x"0a",x"64",x"61",x"65"),
  1604 => (x"54",x"41",x"46",x"00"),
  1605 => (x"20",x"20",x"36",x"31"),
  1606 => (x"41",x"46",x"00",x"20"),
  1607 => (x"20",x"32",x"33",x"54"),
  1608 => (x"50",x"00",x"20",x"20"),
  1609 => (x"69",x"74",x"72",x"61"),
  1610 => (x"6e",x"6f",x"69",x"74"),
  1611 => (x"6e",x"75",x"6f",x"63"),
  1612 => (x"64",x"25",x"20",x"74"),
  1613 => (x"75",x"48",x"00",x"0a"),
  1614 => (x"6e",x"69",x"74",x"6e"),
  1615 => (x"6f",x"66",x"20",x"67"),
  1616 => (x"69",x"66",x"20",x"72"),
  1617 => (x"79",x"73",x"65",x"6c"),
  1618 => (x"6d",x"65",x"74",x"73"),
  1619 => (x"41",x"46",x"00",x"0a"),
  1620 => (x"20",x"32",x"33",x"54"),
  1621 => (x"46",x"00",x"20",x"20"),
  1622 => (x"36",x"31",x"54",x"41"),
  1623 => (x"00",x"20",x"20",x"20"),
  1624 => (x"73",x"75",x"6c",x"43"),
  1625 => (x"20",x"72",x"65",x"74"),
  1626 => (x"65",x"7a",x"69",x"73"),
  1627 => (x"64",x"25",x"20",x"3a"),
  1628 => (x"6c",x"43",x"20",x"2c"),
  1629 => (x"65",x"74",x"73",x"75"),
  1630 => (x"61",x"6d",x"20",x"72"),
  1631 => (x"20",x"2c",x"6b",x"73"),
  1632 => (x"00",x"0a",x"64",x"25"),
  1633 => (x"63",x"65",x"68",x"43"),
  1634 => (x"6d",x"75",x"73",x"6b"),
  1635 => (x"67",x"6e",x"69",x"6d"),
  1636 => (x"6f",x"72",x"66",x"20"),
  1637 => (x"64",x"25",x"20",x"6d"),
  1638 => (x"20",x"6f",x"74",x"20"),
  1639 => (x"2e",x"2e",x"64",x"25"),
  1640 => (x"25",x"00",x"20",x"2e"),
  1641 => (x"25",x"00",x"0a",x"64"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
