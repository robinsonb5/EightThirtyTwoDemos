library ieee;
use ieee.std_logic_1164.all;

package SoC_Peripheral_config is
	constant SoC_PeripheralBit : integer := 31;
	constant SoC_BlockBits : integer := 4;
	constant SoC_Block_HighBit : integer := 11;
	constant SoC_Block_LowBit : integer := 8;
end package;

