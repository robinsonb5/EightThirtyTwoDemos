
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"d4",x"01"),
     1 => (x"18",x"0e",x"87",x"d7"),
     2 => (x"3e",x"27",x"0e",x"1e"),
     3 => (x"0f",x"00",x"00",x"00"),
     4 => (x"80",x"ff",x"48",x"26"),
     5 => (x"27",x"4f",x"08",x"26"),
     6 => (x"00",x"00",x"00",x"23"),
     7 => (x"00",x"30",x"27",x"4f"),
     8 => (x"c2",x"4f",x"00",x"00"),
     9 => (x"27",x"4e",x"c0",x"c0"),
    10 => (x"00",x"00",x"16",x"23"),
    11 => (x"87",x"fd",x"00",x"0f"),
    12 => (x"4e",x"c0",x"f0",x"c1"),
    13 => (x"00",x"00",x"3d",x"27"),
    14 => (x"fd",x"00",x"0f",x"00"),
    15 => (x"1e",x"4f",x"4f",x"87"),
    16 => (x"ff",x"1e",x"1e",x"72"),
    17 => (x"48",x"6a",x"4a",x"c0"),
    18 => (x"c4",x"98",x"c0",x"c4"),
    19 => (x"02",x"6e",x"58",x"a6"),
    20 => (x"cc",x"87",x"f3",x"ff"),
    21 => (x"66",x"cc",x"7a",x"66"),
    22 => (x"4a",x"26",x"26",x"48"),
    23 => (x"5e",x"0e",x"4f",x"26"),
    24 => (x"5d",x"5c",x"5b",x"5a"),
    25 => (x"4b",x"66",x"d4",x"0e"),
    26 => (x"4c",x"13",x"4d",x"c0"),
    27 => (x"c0",x"02",x"9c",x"74"),
    28 => (x"4a",x"74",x"87",x"d6"),
    29 => (x"3f",x"27",x"1e",x"72"),
    30 => (x"0f",x"00",x"00",x"00"),
    31 => (x"85",x"c1",x"86",x"c4"),
    32 => (x"9c",x"74",x"4c",x"13"),
    33 => (x"87",x"ea",x"ff",x"05"),
    34 => (x"4d",x"26",x"48",x"75"),
    35 => (x"4b",x"26",x"4c",x"26"),
    36 => (x"4f",x"26",x"4a",x"26"),
    37 => (x"5b",x"5a",x"5e",x"0e"),
    38 => (x"1e",x"0e",x"5d",x"5c"),
    39 => (x"76",x"4d",x"66",x"d8"),
    40 => (x"c0",x"79",x"c0",x"49"),
    41 => (x"c0",x"03",x"ad",x"b7"),
    42 => (x"ed",x"c0",x"87",x"cd"),
    43 => (x"00",x"3f",x"27",x"1e"),
    44 => (x"c4",x"0f",x"00",x"00"),
    45 => (x"75",x"8d",x"0d",x"86"),
    46 => (x"c2",x"c1",x"02",x"9d"),
    47 => (x"75",x"4c",x"c0",x"87"),
    48 => (x"2a",x"b7",x"dc",x"4a"),
    49 => (x"9b",x"cf",x"4b",x"72"),
    50 => (x"9b",x"73",x"35",x"c4"),
    51 => (x"87",x"c4",x"c0",x"02"),
    52 => (x"79",x"c1",x"49",x"76"),
    53 => (x"06",x"ab",x"b7",x"c9"),
    54 => (x"c0",x"87",x"c6",x"c0"),
    55 => (x"c3",x"c0",x"83",x"f7"),
    56 => (x"83",x"f0",x"c0",x"87"),
    57 => (x"ca",x"c0",x"02",x"6e"),
    58 => (x"27",x"1e",x"73",x"87"),
    59 => (x"00",x"00",x"00",x"3f"),
    60 => (x"c1",x"86",x"c4",x"0f"),
    61 => (x"ac",x"b7",x"c8",x"84"),
    62 => (x"87",x"c3",x"ff",x"04"),
    63 => (x"c0",x"87",x"cb",x"c0"),
    64 => (x"3f",x"27",x"1e",x"f0"),
    65 => (x"0f",x"00",x"00",x"00"),
    66 => (x"48",x"c0",x"86",x"c4"),
    67 => (x"26",x"4d",x"26",x"26"),
    68 => (x"26",x"4b",x"26",x"4c"),
    69 => (x"0e",x"4f",x"26",x"4a"),
    70 => (x"5c",x"5b",x"5a",x"5e"),
    71 => (x"c0",x"1e",x"0e",x"5d"),
    72 => (x"c0",x"49",x"76",x"4c"),
    73 => (x"4b",x"a6",x"dc",x"79"),
    74 => (x"d8",x"4a",x"66",x"d8"),
    75 => (x"80",x"c1",x"48",x"66"),
    76 => (x"12",x"58",x"a6",x"dc"),
    77 => (x"c0",x"c0",x"c1",x"4d"),
    78 => (x"c4",x"95",x"c0",x"c0"),
    79 => (x"4d",x"95",x"b7",x"c0"),
    80 => (x"c4",x"02",x"9d",x"75"),
    81 => (x"02",x"6e",x"87",x"d2"),
    82 => (x"76",x"87",x"d7",x"c3"),
    83 => (x"75",x"79",x"c0",x"49"),
    84 => (x"ad",x"e3",x"c1",x"4a"),
    85 => (x"87",x"dd",x"c2",x"02"),
    86 => (x"02",x"aa",x"e4",x"c1"),
    87 => (x"c1",x"87",x"d8",x"c0"),
    88 => (x"c2",x"02",x"aa",x"ec"),
    89 => (x"f3",x"c1",x"87",x"c8"),
    90 => (x"e8",x"c1",x"02",x"aa"),
    91 => (x"aa",x"f8",x"c1",x"87"),
    92 => (x"87",x"f2",x"c0",x"02"),
    93 => (x"ca",x"87",x"d3",x"c2"),
    94 => (x"1a",x"08",x"27",x"1e"),
    95 => (x"c4",x"1e",x"00",x"00"),
    96 => (x"c4",x"4a",x"73",x"83"),
    97 => (x"27",x"1e",x"6a",x"8a"),
    98 => (x"00",x"00",x"00",x"94"),
    99 => (x"70",x"86",x"cc",x"0f"),
   100 => (x"72",x"4c",x"74",x"4a"),
   101 => (x"1a",x"08",x"27",x"84"),
   102 => (x"27",x"1e",x"00",x"00"),
   103 => (x"00",x"00",x"00",x"5e"),
   104 => (x"c2",x"86",x"c4",x"0f"),
   105 => (x"1e",x"d0",x"87",x"d4"),
   106 => (x"00",x"1a",x"08",x"27"),
   107 => (x"83",x"c4",x"1e",x"00"),
   108 => (x"8a",x"c4",x"4a",x"73"),
   109 => (x"94",x"27",x"1e",x"6a"),
   110 => (x"0f",x"00",x"00",x"00"),
   111 => (x"4a",x"70",x"86",x"cc"),
   112 => (x"84",x"72",x"4c",x"74"),
   113 => (x"00",x"1a",x"08",x"27"),
   114 => (x"5e",x"27",x"1e",x"00"),
   115 => (x"0f",x"00",x"00",x"00"),
   116 => (x"e5",x"c1",x"86",x"c4"),
   117 => (x"73",x"83",x"c4",x"87"),
   118 => (x"6a",x"8a",x"c4",x"4a"),
   119 => (x"00",x"5e",x"27",x"1e"),
   120 => (x"c4",x"0f",x"00",x"00"),
   121 => (x"74",x"4a",x"70",x"86"),
   122 => (x"c1",x"84",x"72",x"4c"),
   123 => (x"49",x"76",x"87",x"cc"),
   124 => (x"c5",x"c1",x"79",x"c1"),
   125 => (x"73",x"83",x"c4",x"87"),
   126 => (x"6a",x"8a",x"c4",x"4a"),
   127 => (x"00",x"3f",x"27",x"1e"),
   128 => (x"c4",x"0f",x"00",x"00"),
   129 => (x"c0",x"84",x"c1",x"86"),
   130 => (x"e5",x"c0",x"87",x"f0"),
   131 => (x"00",x"3f",x"27",x"1e"),
   132 => (x"c4",x"0f",x"00",x"00"),
   133 => (x"27",x"1e",x"75",x"86"),
   134 => (x"00",x"00",x"00",x"3f"),
   135 => (x"c0",x"86",x"c4",x"0f"),
   136 => (x"e5",x"c0",x"87",x"d8"),
   137 => (x"c7",x"c0",x"05",x"ad"),
   138 => (x"c1",x"49",x"76",x"87"),
   139 => (x"87",x"ca",x"c0",x"79"),
   140 => (x"3f",x"27",x"1e",x"75"),
   141 => (x"0f",x"00",x"00",x"00"),
   142 => (x"66",x"d8",x"86",x"c4"),
   143 => (x"48",x"66",x"d8",x"4a"),
   144 => (x"a6",x"dc",x"80",x"c1"),
   145 => (x"c1",x"4d",x"12",x"58"),
   146 => (x"c0",x"c0",x"c0",x"c0"),
   147 => (x"b7",x"c0",x"c4",x"95"),
   148 => (x"9d",x"75",x"4d",x"95"),
   149 => (x"87",x"ee",x"fb",x"05"),
   150 => (x"26",x"26",x"48",x"74"),
   151 => (x"26",x"4c",x"26",x"4d"),
   152 => (x"26",x"4a",x"26",x"4b"),
   153 => (x"00",x"00",x"00",x"4f"),
   154 => (x"1e",x"75",x"1e",x"00"),
   155 => (x"c3",x"4d",x"d4",x"ff"),
   156 => (x"6d",x"7d",x"49",x"ff"),
   157 => (x"71",x"38",x"c8",x"48"),
   158 => (x"c8",x"b0",x"6d",x"7d"),
   159 => (x"6d",x"7d",x"71",x"38"),
   160 => (x"71",x"38",x"c8",x"b0"),
   161 => (x"c8",x"b0",x"6d",x"7d"),
   162 => (x"26",x"4d",x"26",x"38"),
   163 => (x"1e",x"75",x"1e",x"4f"),
   164 => (x"c3",x"4d",x"d4",x"ff"),
   165 => (x"6d",x"7d",x"49",x"ff"),
   166 => (x"71",x"30",x"c8",x"48"),
   167 => (x"c8",x"b0",x"6d",x"7d"),
   168 => (x"6d",x"7d",x"71",x"30"),
   169 => (x"71",x"30",x"c8",x"b0"),
   170 => (x"26",x"b0",x"6d",x"7d"),
   171 => (x"1e",x"4f",x"26",x"4d"),
   172 => (x"d4",x"ff",x"1e",x"75"),
   173 => (x"49",x"66",x"cc",x"4d"),
   174 => (x"7d",x"48",x"66",x"c8"),
   175 => (x"02",x"67",x"e6",x"fe"),
   176 => (x"d8",x"07",x"31",x"c9"),
   177 => (x"09",x"7d",x"09",x"39"),
   178 => (x"09",x"7d",x"09",x"39"),
   179 => (x"09",x"7d",x"09",x"39"),
   180 => (x"d0",x"7d",x"09",x"39"),
   181 => (x"c9",x"7d",x"70",x"38"),
   182 => (x"c3",x"49",x"c0",x"f1"),
   183 => (x"08",x"6d",x"48",x"ff"),
   184 => (x"87",x"c7",x"05",x"a8"),
   185 => (x"89",x"c1",x"7d",x"08"),
   186 => (x"26",x"87",x"f3",x"05"),
   187 => (x"1e",x"4f",x"26",x"4d"),
   188 => (x"c3",x"49",x"d4",x"ff"),
   189 => (x"79",x"ff",x"48",x"c8"),
   190 => (x"87",x"fa",x"05",x"80"),
   191 => (x"5e",x"0e",x"4f",x"26"),
   192 => (x"5d",x"5c",x"5b",x"5a"),
   193 => (x"f0",x"ff",x"c0",x"0e"),
   194 => (x"c1",x"4d",x"f7",x"c1"),
   195 => (x"c0",x"c0",x"c0",x"c0"),
   196 => (x"ef",x"27",x"4b",x"c0"),
   197 => (x"0f",x"00",x"00",x"02"),
   198 => (x"4c",x"df",x"f8",x"c4"),
   199 => (x"1e",x"75",x"1e",x"c0"),
   200 => (x"00",x"02",x"af",x"27"),
   201 => (x"86",x"c8",x"0f",x"00"),
   202 => (x"b7",x"c1",x"4a",x"70"),
   203 => (x"ef",x"c0",x"05",x"aa"),
   204 => (x"49",x"d4",x"ff",x"87"),
   205 => (x"73",x"79",x"ff",x"c3"),
   206 => (x"f0",x"e1",x"c0",x"1e"),
   207 => (x"27",x"1e",x"e9",x"c1"),
   208 => (x"00",x"00",x"02",x"af"),
   209 => (x"70",x"86",x"c8",x"0f"),
   210 => (x"05",x"9a",x"72",x"4a"),
   211 => (x"ff",x"87",x"cb",x"c0"),
   212 => (x"ff",x"c3",x"49",x"d4"),
   213 => (x"c0",x"48",x"c1",x"79"),
   214 => (x"ef",x"27",x"87",x"d0"),
   215 => (x"0f",x"00",x"00",x"02"),
   216 => (x"9c",x"74",x"8c",x"c1"),
   217 => (x"87",x"f4",x"fe",x"05"),
   218 => (x"4d",x"26",x"48",x"c0"),
   219 => (x"4b",x"26",x"4c",x"26"),
   220 => (x"4f",x"26",x"4a",x"26"),
   221 => (x"5b",x"5a",x"5e",x"0e"),
   222 => (x"ff",x"c0",x"0e",x"5c"),
   223 => (x"4c",x"c1",x"c1",x"f0"),
   224 => (x"c3",x"49",x"d4",x"ff"),
   225 => (x"35",x"27",x"79",x"ff"),
   226 => (x"1e",x"00",x"00",x"18"),
   227 => (x"00",x"00",x"5e",x"27"),
   228 => (x"86",x"c4",x"0f",x"00"),
   229 => (x"1e",x"c0",x"4b",x"d3"),
   230 => (x"af",x"27",x"1e",x"74"),
   231 => (x"0f",x"00",x"00",x"02"),
   232 => (x"4a",x"70",x"86",x"c8"),
   233 => (x"c0",x"05",x"9a",x"72"),
   234 => (x"d4",x"ff",x"87",x"cb"),
   235 => (x"79",x"ff",x"c3",x"49"),
   236 => (x"d0",x"c0",x"48",x"c1"),
   237 => (x"02",x"ef",x"27",x"87"),
   238 => (x"c1",x"0f",x"00",x"00"),
   239 => (x"05",x"9b",x"73",x"8b"),
   240 => (x"c0",x"87",x"d3",x"ff"),
   241 => (x"26",x"4c",x"26",x"48"),
   242 => (x"26",x"4a",x"26",x"4b"),
   243 => (x"5a",x"5e",x"0e",x"4f"),
   244 => (x"0e",x"5d",x"5c",x"5b"),
   245 => (x"4d",x"ff",x"c3",x"1e"),
   246 => (x"27",x"4c",x"d4",x"ff"),
   247 => (x"00",x"00",x"02",x"ef"),
   248 => (x"1e",x"ea",x"c6",x"0f"),
   249 => (x"c1",x"f0",x"e1",x"c0"),
   250 => (x"af",x"27",x"1e",x"c8"),
   251 => (x"0f",x"00",x"00",x"02"),
   252 => (x"4a",x"70",x"86",x"c8"),
   253 => (x"2c",x"27",x"1e",x"72"),
   254 => (x"1e",x"00",x"00",x"05"),
   255 => (x"00",x"01",x"17",x"27"),
   256 => (x"86",x"c8",x"0f",x"00"),
   257 => (x"02",x"aa",x"b7",x"c1"),
   258 => (x"27",x"87",x"cb",x"c0"),
   259 => (x"00",x"00",x"03",x"74"),
   260 => (x"c3",x"48",x"c0",x"0f"),
   261 => (x"8d",x"27",x"87",x"c9"),
   262 => (x"0f",x"00",x"00",x"02"),
   263 => (x"ff",x"cf",x"4a",x"70"),
   264 => (x"ea",x"c6",x"9a",x"ff"),
   265 => (x"c0",x"02",x"aa",x"b7"),
   266 => (x"74",x"27",x"87",x"cb"),
   267 => (x"0f",x"00",x"00",x"03"),
   268 => (x"ea",x"c2",x"48",x"c0"),
   269 => (x"76",x"7c",x"75",x"87"),
   270 => (x"79",x"f1",x"c0",x"49"),
   271 => (x"00",x"02",x"fe",x"27"),
   272 => (x"4a",x"70",x"0f",x"00"),
   273 => (x"c1",x"02",x"9a",x"72"),
   274 => (x"1e",x"c0",x"87",x"eb"),
   275 => (x"c1",x"f0",x"ff",x"c0"),
   276 => (x"af",x"27",x"1e",x"fa"),
   277 => (x"0f",x"00",x"00",x"02"),
   278 => (x"4b",x"70",x"86",x"c8"),
   279 => (x"c1",x"05",x"9b",x"73"),
   280 => (x"1e",x"73",x"87",x"c3"),
   281 => (x"00",x"04",x"ea",x"27"),
   282 => (x"17",x"27",x"1e",x"00"),
   283 => (x"0f",x"00",x"00",x"01"),
   284 => (x"7c",x"75",x"86",x"c8"),
   285 => (x"9b",x"75",x"4b",x"6c"),
   286 => (x"f6",x"27",x"1e",x"73"),
   287 => (x"1e",x"00",x"00",x"04"),
   288 => (x"00",x"01",x"17",x"27"),
   289 => (x"86",x"c8",x"0f",x"00"),
   290 => (x"7c",x"75",x"7c",x"75"),
   291 => (x"7c",x"75",x"7c",x"75"),
   292 => (x"c0",x"c1",x"4a",x"73"),
   293 => (x"02",x"9a",x"72",x"9a"),
   294 => (x"c1",x"87",x"c5",x"c0"),
   295 => (x"87",x"ff",x"c0",x"48"),
   296 => (x"fa",x"c0",x"48",x"c0"),
   297 => (x"27",x"1e",x"73",x"87"),
   298 => (x"00",x"00",x"05",x"04"),
   299 => (x"01",x"17",x"27",x"1e"),
   300 => (x"c8",x"0f",x"00",x"00"),
   301 => (x"c2",x"49",x"6e",x"86"),
   302 => (x"c0",x"05",x"a9",x"b7"),
   303 => (x"10",x"27",x"87",x"d3"),
   304 => (x"1e",x"00",x"00",x"05"),
   305 => (x"00",x"01",x"17",x"27"),
   306 => (x"86",x"c4",x"0f",x"00"),
   307 => (x"ce",x"c0",x"48",x"c0"),
   308 => (x"c1",x"48",x"6e",x"87"),
   309 => (x"58",x"a6",x"c4",x"88"),
   310 => (x"df",x"fd",x"05",x"6e"),
   311 => (x"26",x"48",x"c0",x"87"),
   312 => (x"4c",x"26",x"4d",x"26"),
   313 => (x"4a",x"26",x"4b",x"26"),
   314 => (x"4d",x"43",x"4f",x"26"),
   315 => (x"20",x"38",x"35",x"44"),
   316 => (x"20",x"0a",x"64",x"25"),
   317 => (x"4d",x"43",x"00",x"20"),
   318 => (x"5f",x"38",x"35",x"44"),
   319 => (x"64",x"25",x"20",x"32"),
   320 => (x"00",x"20",x"20",x"0a"),
   321 => (x"35",x"44",x"4d",x"43"),
   322 => (x"64",x"25",x"20",x"38"),
   323 => (x"00",x"20",x"20",x"0a"),
   324 => (x"43",x"48",x"44",x"53"),
   325 => (x"69",x"6e",x"49",x"20"),
   326 => (x"6c",x"61",x"69",x"74"),
   327 => (x"74",x"61",x"7a",x"69"),
   328 => (x"20",x"6e",x"6f",x"69"),
   329 => (x"6f",x"72",x"72",x"65"),
   330 => (x"00",x"0a",x"21",x"72"),
   331 => (x"5f",x"64",x"6d",x"63"),
   332 => (x"38",x"44",x"4d",x"43"),
   333 => (x"73",x"65",x"72",x"20"),
   334 => (x"73",x"6e",x"6f",x"70"),
   335 => (x"25",x"20",x"3a",x"65"),
   336 => (x"0e",x"00",x"0a",x"64"),
   337 => (x"5c",x"5b",x"5a",x"5e"),
   338 => (x"ff",x"1e",x"0e",x"5d"),
   339 => (x"c0",x"c8",x"4c",x"d0"),
   340 => (x"65",x"27",x"4b",x"c0"),
   341 => (x"49",x"00",x"00",x"02"),
   342 => (x"60",x"27",x"79",x"c1"),
   343 => (x"1e",x"00",x"00",x"06"),
   344 => (x"00",x"00",x"5e",x"27"),
   345 => (x"86",x"c4",x"0f",x"00"),
   346 => (x"48",x"6c",x"4d",x"c7"),
   347 => (x"a6",x"c4",x"98",x"73"),
   348 => (x"c0",x"02",x"6e",x"58"),
   349 => (x"48",x"6c",x"87",x"cc"),
   350 => (x"a6",x"c4",x"98",x"73"),
   351 => (x"ff",x"05",x"6e",x"58"),
   352 => (x"7c",x"c0",x"87",x"f4"),
   353 => (x"00",x"02",x"ef",x"27"),
   354 => (x"48",x"6c",x"0f",x"00"),
   355 => (x"a6",x"c4",x"98",x"73"),
   356 => (x"c0",x"02",x"6e",x"58"),
   357 => (x"48",x"6c",x"87",x"cc"),
   358 => (x"a6",x"c4",x"98",x"73"),
   359 => (x"ff",x"05",x"6e",x"58"),
   360 => (x"7c",x"c1",x"87",x"f4"),
   361 => (x"e5",x"c0",x"1e",x"c0"),
   362 => (x"1e",x"c0",x"c1",x"d0"),
   363 => (x"00",x"02",x"af",x"27"),
   364 => (x"86",x"c8",x"0f",x"00"),
   365 => (x"b7",x"c1",x"4a",x"70"),
   366 => (x"c2",x"c0",x"05",x"aa"),
   367 => (x"c2",x"4d",x"c1",x"87"),
   368 => (x"c0",x"05",x"ad",x"b7"),
   369 => (x"5b",x"27",x"87",x"d3"),
   370 => (x"1e",x"00",x"00",x"06"),
   371 => (x"00",x"00",x"5e",x"27"),
   372 => (x"86",x"c4",x"0f",x"00"),
   373 => (x"f7",x"c1",x"48",x"c0"),
   374 => (x"75",x"8d",x"c1",x"87"),
   375 => (x"c9",x"fe",x"05",x"9d"),
   376 => (x"03",x"cd",x"27",x"87"),
   377 => (x"27",x"0f",x"00",x"00"),
   378 => (x"00",x"00",x"02",x"69"),
   379 => (x"02",x"65",x"27",x"58"),
   380 => (x"05",x"bf",x"00",x"00"),
   381 => (x"c1",x"87",x"d0",x"c0"),
   382 => (x"f0",x"ff",x"c0",x"1e"),
   383 => (x"27",x"1e",x"d0",x"c1"),
   384 => (x"00",x"00",x"02",x"af"),
   385 => (x"ff",x"86",x"c8",x"0f"),
   386 => (x"ff",x"c3",x"49",x"d4"),
   387 => (x"08",x"f6",x"27",x"79"),
   388 => (x"27",x"0f",x"00",x"00"),
   389 => (x"00",x"00",x"1a",x"30"),
   390 => (x"1a",x"2c",x"27",x"58"),
   391 => (x"1e",x"bf",x"00",x"00"),
   392 => (x"00",x"06",x"64",x"27"),
   393 => (x"17",x"27",x"1e",x"00"),
   394 => (x"0f",x"00",x"00",x"01"),
   395 => (x"48",x"6c",x"86",x"c8"),
   396 => (x"a6",x"c4",x"98",x"73"),
   397 => (x"c0",x"02",x"6e",x"58"),
   398 => (x"48",x"6c",x"87",x"cc"),
   399 => (x"a6",x"c4",x"98",x"73"),
   400 => (x"ff",x"05",x"6e",x"58"),
   401 => (x"7c",x"c0",x"87",x"f4"),
   402 => (x"c3",x"49",x"d4",x"ff"),
   403 => (x"48",x"c1",x"79",x"ff"),
   404 => (x"26",x"4d",x"26",x"26"),
   405 => (x"26",x"4b",x"26",x"4c"),
   406 => (x"49",x"4f",x"26",x"4a"),
   407 => (x"00",x"52",x"52",x"45"),
   408 => (x"00",x"49",x"50",x"53"),
   409 => (x"63",x"20",x"44",x"53"),
   410 => (x"20",x"64",x"72",x"61"),
   411 => (x"65",x"7a",x"69",x"73"),
   412 => (x"20",x"73",x"69",x"20"),
   413 => (x"00",x"0a",x"64",x"25"),
   414 => (x"5b",x"5a",x"5e",x"0e"),
   415 => (x"1e",x"0e",x"5d",x"5c"),
   416 => (x"ff",x"4d",x"ff",x"c3"),
   417 => (x"7c",x"75",x"4c",x"d4"),
   418 => (x"48",x"bf",x"d0",x"ff"),
   419 => (x"98",x"c0",x"c0",x"c8"),
   420 => (x"6e",x"58",x"a6",x"c4"),
   421 => (x"87",x"d2",x"c0",x"02"),
   422 => (x"4a",x"c0",x"c0",x"c8"),
   423 => (x"48",x"bf",x"d0",x"ff"),
   424 => (x"a6",x"c4",x"98",x"72"),
   425 => (x"ff",x"05",x"6e",x"58"),
   426 => (x"d0",x"ff",x"87",x"f2"),
   427 => (x"79",x"c1",x"c4",x"49"),
   428 => (x"66",x"d8",x"7c",x"75"),
   429 => (x"f0",x"ff",x"c0",x"1e"),
   430 => (x"27",x"1e",x"d8",x"c1"),
   431 => (x"00",x"00",x"02",x"af"),
   432 => (x"70",x"86",x"c8",x"0f"),
   433 => (x"02",x"9a",x"72",x"4a"),
   434 => (x"27",x"87",x"d3",x"c0"),
   435 => (x"00",x"00",x"07",x"80"),
   436 => (x"00",x"5e",x"27",x"1e"),
   437 => (x"c4",x"0f",x"00",x"00"),
   438 => (x"c2",x"48",x"c1",x"86"),
   439 => (x"7c",x"75",x"87",x"d7"),
   440 => (x"76",x"7c",x"fe",x"c3"),
   441 => (x"dc",x"79",x"c0",x"49"),
   442 => (x"72",x"4a",x"bf",x"66"),
   443 => (x"2b",x"b7",x"d8",x"4b"),
   444 => (x"98",x"75",x"48",x"73"),
   445 => (x"4b",x"72",x"7c",x"70"),
   446 => (x"73",x"2b",x"b7",x"d0"),
   447 => (x"70",x"98",x"75",x"48"),
   448 => (x"c8",x"4b",x"72",x"7c"),
   449 => (x"48",x"73",x"2b",x"b7"),
   450 => (x"7c",x"70",x"98",x"75"),
   451 => (x"98",x"75",x"48",x"72"),
   452 => (x"66",x"dc",x"7c",x"70"),
   453 => (x"c0",x"80",x"c4",x"48"),
   454 => (x"6e",x"58",x"a6",x"e0"),
   455 => (x"c4",x"80",x"c1",x"48"),
   456 => (x"49",x"6e",x"58",x"a6"),
   457 => (x"a9",x"b7",x"c0",x"c2"),
   458 => (x"87",x"fb",x"fe",x"04"),
   459 => (x"7c",x"75",x"7c",x"75"),
   460 => (x"da",x"d8",x"7c",x"75"),
   461 => (x"7c",x"75",x"4b",x"e0"),
   462 => (x"9a",x"75",x"4a",x"6c"),
   463 => (x"c0",x"05",x"9a",x"72"),
   464 => (x"8b",x"c1",x"87",x"c8"),
   465 => (x"ff",x"05",x"9b",x"73"),
   466 => (x"7c",x"75",x"87",x"ec"),
   467 => (x"48",x"bf",x"d0",x"ff"),
   468 => (x"98",x"c0",x"c0",x"c8"),
   469 => (x"6e",x"58",x"a6",x"c4"),
   470 => (x"87",x"d2",x"c0",x"02"),
   471 => (x"4a",x"c0",x"c0",x"c8"),
   472 => (x"48",x"bf",x"d0",x"ff"),
   473 => (x"a6",x"c4",x"98",x"72"),
   474 => (x"ff",x"05",x"6e",x"58"),
   475 => (x"d0",x"ff",x"87",x"f2"),
   476 => (x"c0",x"79",x"c0",x"49"),
   477 => (x"4d",x"26",x"26",x"48"),
   478 => (x"4b",x"26",x"4c",x"26"),
   479 => (x"4f",x"26",x"4a",x"26"),
   480 => (x"74",x"69",x"72",x"57"),
   481 => (x"61",x"66",x"20",x"65"),
   482 => (x"64",x"65",x"6c",x"69"),
   483 => (x"5e",x"0e",x"00",x"0a"),
   484 => (x"5d",x"5c",x"5b",x"5a"),
   485 => (x"66",x"d8",x"1e",x"0e"),
   486 => (x"4b",x"66",x"dc",x"4c"),
   487 => (x"79",x"c0",x"49",x"76"),
   488 => (x"df",x"cd",x"ee",x"c5"),
   489 => (x"49",x"d4",x"ff",x"4d"),
   490 => (x"ff",x"79",x"ff",x"c3"),
   491 => (x"c3",x"4a",x"bf",x"d4"),
   492 => (x"fe",x"c3",x"9a",x"ff"),
   493 => (x"c1",x"05",x"aa",x"b7"),
   494 => (x"28",x"27",x"87",x"e5"),
   495 => (x"49",x"00",x"00",x"1a"),
   496 => (x"b7",x"c4",x"79",x"c0"),
   497 => (x"e4",x"c0",x"04",x"ab"),
   498 => (x"02",x"69",x"27",x"87"),
   499 => (x"70",x"0f",x"00",x"00"),
   500 => (x"c4",x"7c",x"72",x"4a"),
   501 => (x"1a",x"28",x"27",x"84"),
   502 => (x"48",x"bf",x"00",x"00"),
   503 => (x"2c",x"27",x"80",x"72"),
   504 => (x"58",x"00",x"00",x"1a"),
   505 => (x"b7",x"c4",x"8b",x"c4"),
   506 => (x"dc",x"ff",x"03",x"ab"),
   507 => (x"ab",x"b7",x"c0",x"87"),
   508 => (x"87",x"e5",x"c0",x"06"),
   509 => (x"c3",x"4d",x"d4",x"ff"),
   510 => (x"4a",x"6d",x"7d",x"ff"),
   511 => (x"c1",x"7c",x"97",x"72"),
   512 => (x"1a",x"28",x"27",x"84"),
   513 => (x"48",x"bf",x"00",x"00"),
   514 => (x"2c",x"27",x"80",x"72"),
   515 => (x"58",x"00",x"00",x"1a"),
   516 => (x"b7",x"c0",x"8b",x"c1"),
   517 => (x"de",x"ff",x"01",x"ab"),
   518 => (x"76",x"4d",x"c1",x"87"),
   519 => (x"c1",x"79",x"c1",x"49"),
   520 => (x"05",x"9d",x"75",x"8d"),
   521 => (x"ff",x"87",x"fe",x"fd"),
   522 => (x"ff",x"c3",x"49",x"d4"),
   523 => (x"26",x"48",x"6e",x"79"),
   524 => (x"4c",x"26",x"4d",x"26"),
   525 => (x"4a",x"26",x"4b",x"26"),
   526 => (x"5e",x"0e",x"4f",x"26"),
   527 => (x"5d",x"5c",x"5b",x"5a"),
   528 => (x"d0",x"ff",x"1e",x"0e"),
   529 => (x"c0",x"c0",x"c8",x"4b"),
   530 => (x"ff",x"4c",x"c0",x"4a"),
   531 => (x"ff",x"c3",x"49",x"d4"),
   532 => (x"72",x"48",x"6b",x"79"),
   533 => (x"58",x"a6",x"c4",x"98"),
   534 => (x"cc",x"c0",x"02",x"6e"),
   535 => (x"72",x"48",x"6b",x"87"),
   536 => (x"58",x"a6",x"c4",x"98"),
   537 => (x"f4",x"ff",x"05",x"6e"),
   538 => (x"7b",x"c1",x"c4",x"87"),
   539 => (x"c3",x"49",x"d4",x"ff"),
   540 => (x"66",x"d8",x"79",x"ff"),
   541 => (x"f0",x"ff",x"c0",x"1e"),
   542 => (x"27",x"1e",x"d1",x"c1"),
   543 => (x"00",x"00",x"02",x"af"),
   544 => (x"70",x"86",x"c8",x"0f"),
   545 => (x"02",x"9d",x"75",x"4d"),
   546 => (x"75",x"87",x"d6",x"c0"),
   547 => (x"1e",x"66",x"dc",x"1e"),
   548 => (x"00",x"08",x"d6",x"27"),
   549 => (x"17",x"27",x"1e",x"00"),
   550 => (x"0f",x"00",x"00",x"01"),
   551 => (x"e8",x"c0",x"86",x"cc"),
   552 => (x"1e",x"c0",x"c8",x"87"),
   553 => (x"1e",x"66",x"e0",x"c0"),
   554 => (x"c8",x"87",x"e3",x"fb"),
   555 => (x"6b",x"4c",x"70",x"86"),
   556 => (x"c4",x"98",x"72",x"48"),
   557 => (x"02",x"6e",x"58",x"a6"),
   558 => (x"6b",x"87",x"cc",x"c0"),
   559 => (x"c4",x"98",x"72",x"48"),
   560 => (x"05",x"6e",x"58",x"a6"),
   561 => (x"c0",x"87",x"f4",x"ff"),
   562 => (x"26",x"48",x"74",x"7b"),
   563 => (x"4c",x"26",x"4d",x"26"),
   564 => (x"4a",x"26",x"4b",x"26"),
   565 => (x"65",x"52",x"4f",x"26"),
   566 => (x"63",x"20",x"64",x"61"),
   567 => (x"61",x"6d",x"6d",x"6f"),
   568 => (x"66",x"20",x"64",x"6e"),
   569 => (x"65",x"6c",x"69",x"61"),
   570 => (x"74",x"61",x"20",x"64"),
   571 => (x"20",x"64",x"25",x"20"),
   572 => (x"29",x"64",x"25",x"28"),
   573 => (x"5e",x"0e",x"00",x"0a"),
   574 => (x"5d",x"5c",x"5b",x"5a"),
   575 => (x"1e",x"c0",x"1e",x"0e"),
   576 => (x"c1",x"f0",x"ff",x"c0"),
   577 => (x"af",x"27",x"1e",x"c9"),
   578 => (x"0f",x"00",x"00",x"02"),
   579 => (x"1e",x"d2",x"86",x"c8"),
   580 => (x"00",x"1a",x"38",x"27"),
   581 => (x"f5",x"f9",x"1e",x"00"),
   582 => (x"c0",x"86",x"c8",x"87"),
   583 => (x"d2",x"85",x"c1",x"4d"),
   584 => (x"ff",x"04",x"ad",x"b7"),
   585 => (x"38",x"27",x"87",x"f7"),
   586 => (x"97",x"00",x"00",x"1a"),
   587 => (x"c0",x"c3",x"4a",x"bf"),
   588 => (x"b7",x"c0",x"c1",x"9a"),
   589 => (x"f2",x"c0",x"05",x"aa"),
   590 => (x"1a",x"3f",x"27",x"87"),
   591 => (x"bf",x"97",x"00",x"00"),
   592 => (x"27",x"32",x"d0",x"4a"),
   593 => (x"00",x"00",x"1a",x"40"),
   594 => (x"c8",x"4b",x"bf",x"97"),
   595 => (x"73",x"4a",x"72",x"33"),
   596 => (x"1a",x"41",x"27",x"b2"),
   597 => (x"bf",x"97",x"00",x"00"),
   598 => (x"73",x"4a",x"72",x"4b"),
   599 => (x"ff",x"ff",x"cf",x"b2"),
   600 => (x"4d",x"72",x"9a",x"ff"),
   601 => (x"35",x"ca",x"85",x"c1"),
   602 => (x"27",x"87",x"cb",x"c3"),
   603 => (x"00",x"00",x"1a",x"41"),
   604 => (x"c1",x"4a",x"bf",x"97"),
   605 => (x"27",x"9a",x"c6",x"32"),
   606 => (x"00",x"00",x"1a",x"42"),
   607 => (x"c7",x"4b",x"bf",x"97"),
   608 => (x"4a",x"72",x"2b",x"b7"),
   609 => (x"3d",x"27",x"b2",x"73"),
   610 => (x"97",x"00",x"00",x"1a"),
   611 => (x"48",x"73",x"4b",x"bf"),
   612 => (x"a6",x"c4",x"98",x"cf"),
   613 => (x"1a",x"3e",x"27",x"58"),
   614 => (x"bf",x"97",x"00",x"00"),
   615 => (x"ca",x"9b",x"c3",x"4b"),
   616 => (x"1a",x"3f",x"27",x"33"),
   617 => (x"bf",x"97",x"00",x"00"),
   618 => (x"73",x"34",x"c2",x"4c"),
   619 => (x"27",x"b3",x"74",x"4b"),
   620 => (x"00",x"00",x"1a",x"40"),
   621 => (x"c3",x"4c",x"bf",x"97"),
   622 => (x"b7",x"c6",x"9c",x"c0"),
   623 => (x"74",x"4b",x"73",x"2c"),
   624 => (x"c4",x"1e",x"73",x"b3"),
   625 => (x"1e",x"72",x"1e",x"66"),
   626 => (x"00",x"0a",x"43",x"27"),
   627 => (x"17",x"27",x"1e",x"00"),
   628 => (x"0f",x"00",x"00",x"01"),
   629 => (x"82",x"c2",x"86",x"d0"),
   630 => (x"30",x"72",x"48",x"c1"),
   631 => (x"1e",x"72",x"4a",x"70"),
   632 => (x"00",x"0a",x"70",x"27"),
   633 => (x"17",x"27",x"1e",x"00"),
   634 => (x"0f",x"00",x"00",x"01"),
   635 => (x"48",x"c1",x"86",x"c8"),
   636 => (x"a6",x"c4",x"30",x"6e"),
   637 => (x"73",x"83",x"c1",x"58"),
   638 => (x"6e",x"95",x"72",x"4d"),
   639 => (x"27",x"1e",x"75",x"1e"),
   640 => (x"00",x"00",x"0a",x"79"),
   641 => (x"01",x"17",x"27",x"1e"),
   642 => (x"cc",x"0f",x"00",x"00"),
   643 => (x"c8",x"49",x"6e",x"86"),
   644 => (x"06",x"a9",x"b7",x"c0"),
   645 => (x"6e",x"87",x"cf",x"c0"),
   646 => (x"c1",x"35",x"c1",x"4a"),
   647 => (x"c0",x"c8",x"2a",x"b7"),
   648 => (x"ff",x"01",x"aa",x"b7"),
   649 => (x"1e",x"75",x"87",x"f3"),
   650 => (x"00",x"0a",x"8f",x"27"),
   651 => (x"17",x"27",x"1e",x"00"),
   652 => (x"0f",x"00",x"00",x"01"),
   653 => (x"48",x"75",x"86",x"c8"),
   654 => (x"26",x"4d",x"26",x"26"),
   655 => (x"26",x"4b",x"26",x"4c"),
   656 => (x"63",x"4f",x"26",x"4a"),
   657 => (x"7a",x"69",x"73",x"5f"),
   658 => (x"75",x"6d",x"5f",x"65"),
   659 => (x"20",x"3a",x"74",x"6c"),
   660 => (x"20",x"2c",x"64",x"25"),
   661 => (x"64",x"61",x"65",x"72"),
   662 => (x"5f",x"6c",x"62",x"5f"),
   663 => (x"3a",x"6e",x"65",x"6c"),
   664 => (x"2c",x"64",x"25",x"20"),
   665 => (x"69",x"73",x"63",x"20"),
   666 => (x"20",x"3a",x"65",x"7a"),
   667 => (x"00",x"0a",x"64",x"25"),
   668 => (x"74",x"6c",x"75",x"4d"),
   669 => (x"0a",x"64",x"25",x"20"),
   670 => (x"20",x"64",x"25",x"00"),
   671 => (x"63",x"6f",x"6c",x"62"),
   672 => (x"6f",x"20",x"73",x"6b"),
   673 => (x"69",x"73",x"20",x"66"),
   674 => (x"25",x"20",x"65",x"7a"),
   675 => (x"25",x"00",x"0a",x"64"),
   676 => (x"6c",x"62",x"20",x"64"),
   677 => (x"73",x"6b",x"63",x"6f"),
   678 => (x"20",x"66",x"6f",x"20"),
   679 => (x"20",x"32",x"31",x"35"),
   680 => (x"65",x"74",x"79",x"62"),
   681 => (x"0e",x"00",x"0a",x"73"),
   682 => (x"5c",x"5b",x"5a",x"5e"),
   683 => (x"66",x"d4",x"0e",x"5d"),
   684 => (x"dc",x"4c",x"c0",x"4d"),
   685 => (x"b7",x"c0",x"49",x"66"),
   686 => (x"fb",x"c0",x"06",x"a9"),
   687 => (x"c1",x"4b",x"15",x"87"),
   688 => (x"c0",x"c0",x"c0",x"c0"),
   689 => (x"b7",x"c0",x"c4",x"93"),
   690 => (x"66",x"d8",x"4b",x"93"),
   691 => (x"c1",x"4a",x"bf",x"97"),
   692 => (x"c0",x"c0",x"c0",x"c0"),
   693 => (x"b7",x"c0",x"c4",x"92"),
   694 => (x"66",x"d8",x"4a",x"92"),
   695 => (x"dc",x"80",x"c1",x"48"),
   696 => (x"b7",x"72",x"58",x"a6"),
   697 => (x"c5",x"c0",x"02",x"ab"),
   698 => (x"c0",x"48",x"c1",x"87"),
   699 => (x"84",x"c1",x"87",x"cc"),
   700 => (x"ac",x"b7",x"66",x"dc"),
   701 => (x"87",x"c5",x"ff",x"04"),
   702 => (x"4d",x"26",x"48",x"c0"),
   703 => (x"4b",x"26",x"4c",x"26"),
   704 => (x"4f",x"26",x"4a",x"26"),
   705 => (x"5b",x"5a",x"5e",x"0e"),
   706 => (x"27",x"0e",x"5d",x"5c"),
   707 => (x"00",x"00",x"1c",x"60"),
   708 => (x"27",x"79",x"c0",x"49"),
   709 => (x"00",x"00",x"19",x"0d"),
   710 => (x"00",x"5e",x"27",x"1e"),
   711 => (x"c4",x"0f",x"00",x"00"),
   712 => (x"1a",x"58",x"27",x"86"),
   713 => (x"c0",x"1e",x"00",x"00"),
   714 => (x"08",x"3a",x"27",x"1e"),
   715 => (x"c8",x"0f",x"00",x"00"),
   716 => (x"72",x"4a",x"70",x"86"),
   717 => (x"d3",x"c0",x"05",x"9a"),
   718 => (x"18",x"39",x"27",x"87"),
   719 => (x"27",x"1e",x"00",x"00"),
   720 => (x"00",x"00",x"00",x"5e"),
   721 => (x"c0",x"86",x"c4",x"0f"),
   722 => (x"87",x"d8",x"cf",x"48"),
   723 => (x"00",x"19",x"1a",x"27"),
   724 => (x"5e",x"27",x"1e",x"00"),
   725 => (x"0f",x"00",x"00",x"00"),
   726 => (x"4c",x"c0",x"86",x"c4"),
   727 => (x"00",x"1c",x"8c",x"27"),
   728 => (x"79",x"c1",x"49",x"00"),
   729 => (x"31",x"27",x"1e",x"c8"),
   730 => (x"1e",x"00",x"00",x"19"),
   731 => (x"00",x"1a",x"8e",x"27"),
   732 => (x"a7",x"27",x"1e",x"00"),
   733 => (x"0f",x"00",x"00",x"0a"),
   734 => (x"4a",x"70",x"86",x"cc"),
   735 => (x"c0",x"05",x"9a",x"72"),
   736 => (x"8c",x"27",x"87",x"c8"),
   737 => (x"49",x"00",x"00",x"1c"),
   738 => (x"1e",x"c8",x"79",x"c0"),
   739 => (x"00",x"19",x"3a",x"27"),
   740 => (x"aa",x"27",x"1e",x"00"),
   741 => (x"1e",x"00",x"00",x"1a"),
   742 => (x"00",x"0a",x"a7",x"27"),
   743 => (x"86",x"cc",x"0f",x"00"),
   744 => (x"9a",x"72",x"4a",x"70"),
   745 => (x"87",x"c8",x"c0",x"05"),
   746 => (x"00",x"1c",x"8c",x"27"),
   747 => (x"79",x"c0",x"49",x"00"),
   748 => (x"00",x"1c",x"8c",x"27"),
   749 => (x"27",x"1e",x"bf",x"00"),
   750 => (x"00",x"00",x"19",x"43"),
   751 => (x"01",x"17",x"27",x"1e"),
   752 => (x"c8",x"0f",x"00",x"00"),
   753 => (x"1c",x"8c",x"27",x"86"),
   754 => (x"02",x"bf",x"00",x"00"),
   755 => (x"27",x"87",x"c0",x"c3"),
   756 => (x"00",x"00",x"1a",x"58"),
   757 => (x"1c",x"16",x"27",x"4d"),
   758 => (x"27",x"4b",x"00",x"00"),
   759 => (x"00",x"00",x"1c",x"56"),
   760 => (x"72",x"4a",x"bf",x"9f"),
   761 => (x"1c",x"56",x"27",x"1e"),
   762 => (x"27",x"4a",x"00",x"00"),
   763 => (x"00",x"00",x"1a",x"58"),
   764 => (x"d0",x"1e",x"72",x"8a"),
   765 => (x"1e",x"c0",x"c8",x"1e"),
   766 => (x"00",x"18",x"6b",x"27"),
   767 => (x"17",x"27",x"1e",x"00"),
   768 => (x"0f",x"00",x"00",x"01"),
   769 => (x"4a",x"73",x"86",x"d4"),
   770 => (x"4c",x"6a",x"82",x"c8"),
   771 => (x"00",x"1c",x"56",x"27"),
   772 => (x"4a",x"bf",x"9f",x"00"),
   773 => (x"b7",x"ea",x"d6",x"c5"),
   774 => (x"d3",x"c0",x"05",x"aa"),
   775 => (x"c8",x"4a",x"73",x"87"),
   776 => (x"27",x"1e",x"6a",x"82"),
   777 => (x"00",x"00",x"12",x"8f"),
   778 => (x"70",x"86",x"c4",x"0f"),
   779 => (x"87",x"e4",x"c0",x"4c"),
   780 => (x"fe",x"c7",x"4a",x"75"),
   781 => (x"4a",x"6a",x"9f",x"82"),
   782 => (x"b7",x"d5",x"e9",x"ca"),
   783 => (x"d3",x"c0",x"02",x"aa"),
   784 => (x"18",x"4d",x"27",x"87"),
   785 => (x"27",x"1e",x"00",x"00"),
   786 => (x"00",x"00",x"00",x"5e"),
   787 => (x"c0",x"86",x"c4",x"0f"),
   788 => (x"87",x"d0",x"cb",x"48"),
   789 => (x"a8",x"27",x"1e",x"74"),
   790 => (x"1e",x"00",x"00",x"18"),
   791 => (x"00",x"01",x"17",x"27"),
   792 => (x"86",x"c8",x"0f",x"00"),
   793 => (x"00",x"1a",x"58",x"27"),
   794 => (x"1e",x"74",x"1e",x"00"),
   795 => (x"00",x"08",x"3a",x"27"),
   796 => (x"86",x"c8",x"0f",x"00"),
   797 => (x"9a",x"72",x"4a",x"70"),
   798 => (x"87",x"c5",x"c0",x"05"),
   799 => (x"e3",x"ca",x"48",x"c0"),
   800 => (x"18",x"c0",x"27",x"87"),
   801 => (x"27",x"1e",x"00",x"00"),
   802 => (x"00",x"00",x"00",x"5e"),
   803 => (x"27",x"86",x"c4",x"0f"),
   804 => (x"00",x"00",x"19",x"56"),
   805 => (x"01",x"17",x"27",x"1e"),
   806 => (x"c4",x"0f",x"00",x"00"),
   807 => (x"27",x"1e",x"c8",x"86"),
   808 => (x"00",x"00",x"19",x"6e"),
   809 => (x"1a",x"aa",x"27",x"1e"),
   810 => (x"27",x"1e",x"00",x"00"),
   811 => (x"00",x"00",x"0a",x"a7"),
   812 => (x"70",x"86",x"cc",x"0f"),
   813 => (x"05",x"9a",x"72",x"4a"),
   814 => (x"27",x"87",x"cb",x"c0"),
   815 => (x"00",x"00",x"1c",x"60"),
   816 => (x"c0",x"79",x"c1",x"49"),
   817 => (x"1e",x"c8",x"87",x"f1"),
   818 => (x"00",x"19",x"77",x"27"),
   819 => (x"8e",x"27",x"1e",x"00"),
   820 => (x"1e",x"00",x"00",x"1a"),
   821 => (x"00",x"0a",x"a7",x"27"),
   822 => (x"86",x"cc",x"0f",x"00"),
   823 => (x"9a",x"72",x"4a",x"70"),
   824 => (x"87",x"d3",x"c0",x"02"),
   825 => (x"00",x"18",x"e7",x"27"),
   826 => (x"17",x"27",x"1e",x"00"),
   827 => (x"0f",x"00",x"00",x"01"),
   828 => (x"48",x"c0",x"86",x"c4"),
   829 => (x"27",x"87",x"ed",x"c8"),
   830 => (x"00",x"00",x"1c",x"56"),
   831 => (x"c1",x"4a",x"bf",x"97"),
   832 => (x"05",x"aa",x"b7",x"d5"),
   833 => (x"27",x"87",x"d0",x"c0"),
   834 => (x"00",x"00",x"1c",x"57"),
   835 => (x"c2",x"4a",x"bf",x"97"),
   836 => (x"02",x"aa",x"b7",x"ea"),
   837 => (x"c0",x"87",x"c5",x"c0"),
   838 => (x"87",x"c8",x"c8",x"48"),
   839 => (x"00",x"1a",x"58",x"27"),
   840 => (x"4a",x"bf",x"97",x"00"),
   841 => (x"aa",x"b7",x"e9",x"c3"),
   842 => (x"87",x"d5",x"c0",x"02"),
   843 => (x"00",x"1a",x"58",x"27"),
   844 => (x"4a",x"bf",x"97",x"00"),
   845 => (x"aa",x"b7",x"eb",x"c3"),
   846 => (x"87",x"c5",x"c0",x"02"),
   847 => (x"e3",x"c7",x"48",x"c0"),
   848 => (x"1a",x"63",x"27",x"87"),
   849 => (x"bf",x"97",x"00",x"00"),
   850 => (x"05",x"9a",x"72",x"4a"),
   851 => (x"27",x"87",x"cf",x"c0"),
   852 => (x"00",x"00",x"1a",x"64"),
   853 => (x"c2",x"4a",x"bf",x"97"),
   854 => (x"c0",x"02",x"aa",x"b7"),
   855 => (x"48",x"c0",x"87",x"c5"),
   856 => (x"27",x"87",x"c1",x"c7"),
   857 => (x"00",x"00",x"1a",x"65"),
   858 => (x"27",x"48",x"bf",x"97"),
   859 => (x"00",x"00",x"1c",x"5c"),
   860 => (x"1c",x"58",x"27",x"58"),
   861 => (x"4a",x"bf",x"00",x"00"),
   862 => (x"8b",x"c1",x"4b",x"72"),
   863 => (x"00",x"1c",x"5c",x"27"),
   864 => (x"79",x"73",x"49",x"00"),
   865 => (x"1e",x"72",x"1e",x"73"),
   866 => (x"00",x"19",x"80",x"27"),
   867 => (x"17",x"27",x"1e",x"00"),
   868 => (x"0f",x"00",x"00",x"01"),
   869 => (x"66",x"27",x"86",x"cc"),
   870 => (x"97",x"00",x"00",x"1a"),
   871 => (x"82",x"74",x"4a",x"bf"),
   872 => (x"00",x"1a",x"67",x"27"),
   873 => (x"4b",x"bf",x"97",x"00"),
   874 => (x"48",x"73",x"33",x"c8"),
   875 => (x"70",x"27",x"80",x"72"),
   876 => (x"58",x"00",x"00",x"1c"),
   877 => (x"00",x"1a",x"68",x"27"),
   878 => (x"48",x"bf",x"97",x"00"),
   879 => (x"00",x"1c",x"84",x"27"),
   880 => (x"60",x"27",x"58",x"00"),
   881 => (x"bf",x"00",x"00",x"1c"),
   882 => (x"87",x"df",x"c3",x"02"),
   883 => (x"04",x"27",x"1e",x"c8"),
   884 => (x"1e",x"00",x"00",x"19"),
   885 => (x"00",x"1a",x"aa",x"27"),
   886 => (x"a7",x"27",x"1e",x"00"),
   887 => (x"0f",x"00",x"00",x"0a"),
   888 => (x"4a",x"70",x"86",x"cc"),
   889 => (x"c0",x"02",x"9a",x"72"),
   890 => (x"48",x"c0",x"87",x"c5"),
   891 => (x"27",x"87",x"f5",x"c4"),
   892 => (x"00",x"00",x"1c",x"58"),
   893 => (x"48",x"73",x"4b",x"bf"),
   894 => (x"88",x"27",x"30",x"c4"),
   895 => (x"58",x"00",x"00",x"1c"),
   896 => (x"00",x"1c",x"7c",x"27"),
   897 => (x"79",x"73",x"49",x"00"),
   898 => (x"00",x"1a",x"7d",x"27"),
   899 => (x"4a",x"bf",x"97",x"00"),
   900 => (x"7c",x"27",x"32",x"c8"),
   901 => (x"97",x"00",x"00",x"1a"),
   902 => (x"4a",x"72",x"4c",x"bf"),
   903 => (x"7e",x"27",x"82",x"74"),
   904 => (x"97",x"00",x"00",x"1a"),
   905 => (x"34",x"d0",x"4c",x"bf"),
   906 => (x"82",x"74",x"4a",x"72"),
   907 => (x"00",x"1a",x"7f",x"27"),
   908 => (x"4c",x"bf",x"97",x"00"),
   909 => (x"4a",x"72",x"34",x"d8"),
   910 => (x"88",x"27",x"82",x"74"),
   911 => (x"49",x"00",x"00",x"1c"),
   912 => (x"4a",x"72",x"79",x"72"),
   913 => (x"00",x"1c",x"80",x"27"),
   914 => (x"72",x"92",x"bf",x"00"),
   915 => (x"1c",x"6c",x"27",x"4a"),
   916 => (x"82",x"bf",x"00",x"00"),
   917 => (x"00",x"1c",x"70",x"27"),
   918 => (x"79",x"72",x"49",x"00"),
   919 => (x"00",x"1a",x"85",x"27"),
   920 => (x"4c",x"bf",x"97",x"00"),
   921 => (x"84",x"27",x"34",x"c8"),
   922 => (x"97",x"00",x"00",x"1a"),
   923 => (x"4c",x"74",x"4d",x"bf"),
   924 => (x"86",x"27",x"84",x"75"),
   925 => (x"97",x"00",x"00",x"1a"),
   926 => (x"35",x"d0",x"4d",x"bf"),
   927 => (x"84",x"75",x"4c",x"74"),
   928 => (x"00",x"1a",x"87",x"27"),
   929 => (x"4d",x"bf",x"97",x"00"),
   930 => (x"35",x"d8",x"9d",x"cf"),
   931 => (x"84",x"75",x"4c",x"74"),
   932 => (x"00",x"1c",x"74",x"27"),
   933 => (x"79",x"74",x"49",x"00"),
   934 => (x"4b",x"73",x"8c",x"c2"),
   935 => (x"48",x"73",x"93",x"74"),
   936 => (x"7c",x"27",x"80",x"72"),
   937 => (x"58",x"00",x"00",x"1c"),
   938 => (x"27",x"87",x"f7",x"c1"),
   939 => (x"00",x"00",x"1a",x"6a"),
   940 => (x"c8",x"4a",x"bf",x"97"),
   941 => (x"1a",x"69",x"27",x"32"),
   942 => (x"bf",x"97",x"00",x"00"),
   943 => (x"73",x"4a",x"72",x"4b"),
   944 => (x"1c",x"84",x"27",x"82"),
   945 => (x"72",x"49",x"00",x"00"),
   946 => (x"c7",x"32",x"c5",x"79"),
   947 => (x"2a",x"c9",x"82",x"ff"),
   948 => (x"00",x"1c",x"7c",x"27"),
   949 => (x"79",x"72",x"49",x"00"),
   950 => (x"00",x"1a",x"6f",x"27"),
   951 => (x"4b",x"bf",x"97",x"00"),
   952 => (x"6e",x"27",x"33",x"c8"),
   953 => (x"97",x"00",x"00",x"1a"),
   954 => (x"4b",x"73",x"4c",x"bf"),
   955 => (x"88",x"27",x"83",x"74"),
   956 => (x"49",x"00",x"00",x"1c"),
   957 => (x"4b",x"73",x"79",x"73"),
   958 => (x"00",x"1c",x"80",x"27"),
   959 => (x"73",x"93",x"bf",x"00"),
   960 => (x"1c",x"6c",x"27",x"4b"),
   961 => (x"83",x"bf",x"00",x"00"),
   962 => (x"00",x"1c",x"78",x"27"),
   963 => (x"79",x"73",x"49",x"00"),
   964 => (x"00",x"1c",x"74",x"27"),
   965 => (x"79",x"c0",x"49",x"00"),
   966 => (x"80",x"72",x"48",x"73"),
   967 => (x"00",x"1c",x"74",x"27"),
   968 => (x"48",x"c1",x"58",x"00"),
   969 => (x"4c",x"26",x"4d",x"26"),
   970 => (x"4a",x"26",x"4b",x"26"),
   971 => (x"5e",x"0e",x"4f",x"26"),
   972 => (x"5d",x"5c",x"5b",x"5a"),
   973 => (x"1c",x"60",x"27",x"0e"),
   974 => (x"02",x"bf",x"00",x"00"),
   975 => (x"d4",x"87",x"cf",x"c0"),
   976 => (x"b7",x"c7",x"4c",x"66"),
   977 => (x"4b",x"66",x"d4",x"2c"),
   978 => (x"c0",x"9b",x"ff",x"c1"),
   979 => (x"66",x"d4",x"87",x"cc"),
   980 => (x"2c",x"b7",x"c8",x"4c"),
   981 => (x"c3",x"4b",x"66",x"d4"),
   982 => (x"58",x"27",x"9b",x"ff"),
   983 => (x"1e",x"00",x"00",x"1a"),
   984 => (x"00",x"1c",x"6c",x"27"),
   985 => (x"74",x"4a",x"bf",x"00"),
   986 => (x"27",x"1e",x"72",x"82"),
   987 => (x"00",x"00",x"08",x"3a"),
   988 => (x"70",x"86",x"c8",x"0f"),
   989 => (x"05",x"9a",x"72",x"4a"),
   990 => (x"c0",x"87",x"c5",x"c0"),
   991 => (x"87",x"f2",x"c0",x"48"),
   992 => (x"00",x"1c",x"60",x"27"),
   993 => (x"c0",x"02",x"bf",x"00"),
   994 => (x"4a",x"73",x"87",x"d7"),
   995 => (x"4a",x"72",x"92",x"c4"),
   996 => (x"00",x"1a",x"58",x"27"),
   997 => (x"4d",x"6a",x"82",x"00"),
   998 => (x"ff",x"ff",x"ff",x"cf"),
   999 => (x"cf",x"c0",x"9d",x"ff"),
  1000 => (x"c2",x"4a",x"73",x"87"),
  1001 => (x"27",x"4a",x"72",x"92"),
  1002 => (x"00",x"00",x"1a",x"58"),
  1003 => (x"4d",x"6a",x"9f",x"82"),
  1004 => (x"4d",x"26",x"48",x"75"),
  1005 => (x"4b",x"26",x"4c",x"26"),
  1006 => (x"4f",x"26",x"4a",x"26"),
  1007 => (x"5b",x"5a",x"5e",x"0e"),
  1008 => (x"cc",x"0e",x"5d",x"5c"),
  1009 => (x"ff",x"ff",x"cf",x"8e"),
  1010 => (x"c0",x"4d",x"f8",x"ff"),
  1011 => (x"27",x"49",x"76",x"4c"),
  1012 => (x"00",x"00",x"1c",x"74"),
  1013 => (x"a6",x"c4",x"79",x"bf"),
  1014 => (x"1c",x"78",x"27",x"49"),
  1015 => (x"79",x"bf",x"00",x"00"),
  1016 => (x"00",x"1c",x"60",x"27"),
  1017 => (x"c0",x"02",x"bf",x"00"),
  1018 => (x"58",x"27",x"87",x"cc"),
  1019 => (x"bf",x"00",x"00",x"1c"),
  1020 => (x"c0",x"32",x"c4",x"4a"),
  1021 => (x"7c",x"27",x"87",x"c9"),
  1022 => (x"bf",x"00",x"00",x"1c"),
  1023 => (x"c8",x"32",x"c4",x"4a"),
  1024 => (x"79",x"72",x"49",x"a6"),
  1025 => (x"66",x"c8",x"4b",x"c0"),
  1026 => (x"06",x"a9",x"c0",x"49"),
  1027 => (x"73",x"87",x"d0",x"c3"),
  1028 => (x"72",x"9a",x"cf",x"4a"),
  1029 => (x"e4",x"c0",x"05",x"9a"),
  1030 => (x"1a",x"58",x"27",x"87"),
  1031 => (x"c8",x"1e",x"00",x"00"),
  1032 => (x"66",x"c8",x"4a",x"66"),
  1033 => (x"cc",x"80",x"c1",x"48"),
  1034 => (x"1e",x"72",x"58",x"a6"),
  1035 => (x"00",x"08",x"3a",x"27"),
  1036 => (x"86",x"c8",x"0f",x"00"),
  1037 => (x"00",x"1a",x"58",x"27"),
  1038 => (x"c3",x"c0",x"4c",x"00"),
  1039 => (x"84",x"e0",x"c0",x"87"),
  1040 => (x"72",x"4a",x"6c",x"97"),
  1041 => (x"cd",x"c2",x"02",x"9a"),
  1042 => (x"4a",x"6c",x"97",x"87"),
  1043 => (x"aa",x"b7",x"e5",x"c3"),
  1044 => (x"87",x"c2",x"c2",x"02"),
  1045 => (x"82",x"cb",x"4a",x"74"),
  1046 => (x"d8",x"4a",x"6a",x"97"),
  1047 => (x"05",x"9a",x"72",x"9a"),
  1048 => (x"74",x"87",x"f3",x"c1"),
  1049 => (x"00",x"5e",x"27",x"1e"),
  1050 => (x"c4",x"0f",x"00",x"00"),
  1051 => (x"c0",x"1e",x"cb",x"86"),
  1052 => (x"74",x"1e",x"66",x"e8"),
  1053 => (x"0a",x"a7",x"27",x"1e"),
  1054 => (x"cc",x"0f",x"00",x"00"),
  1055 => (x"72",x"4a",x"70",x"86"),
  1056 => (x"d1",x"c1",x"05",x"9a"),
  1057 => (x"dc",x"4b",x"74",x"87"),
  1058 => (x"66",x"e0",x"c0",x"83"),
  1059 => (x"6b",x"82",x"c4",x"4a"),
  1060 => (x"da",x"4b",x"74",x"7a"),
  1061 => (x"66",x"e0",x"c0",x"83"),
  1062 => (x"9f",x"82",x"c8",x"4a"),
  1063 => (x"7a",x"70",x"48",x"6b"),
  1064 => (x"60",x"27",x"4d",x"72"),
  1065 => (x"bf",x"00",x"00",x"1c"),
  1066 => (x"87",x"d5",x"c0",x"02"),
  1067 => (x"82",x"d4",x"4a",x"74"),
  1068 => (x"c0",x"4a",x"6a",x"9f"),
  1069 => (x"72",x"9a",x"ff",x"ff"),
  1070 => (x"c4",x"30",x"d0",x"48"),
  1071 => (x"c4",x"c0",x"58",x"a6"),
  1072 => (x"c0",x"49",x"76",x"87"),
  1073 => (x"6d",x"48",x"6e",x"79"),
  1074 => (x"c0",x"7d",x"70",x"80"),
  1075 => (x"c0",x"49",x"66",x"e0"),
  1076 => (x"c1",x"48",x"c1",x"79"),
  1077 => (x"83",x"c1",x"87",x"ce"),
  1078 => (x"04",x"ab",x"66",x"c8"),
  1079 => (x"cf",x"87",x"f0",x"fc"),
  1080 => (x"f8",x"ff",x"ff",x"ff"),
  1081 => (x"1c",x"60",x"27",x"4d"),
  1082 => (x"02",x"bf",x"00",x"00"),
  1083 => (x"6e",x"87",x"f3",x"c0"),
  1084 => (x"0f",x"2e",x"27",x"1e"),
  1085 => (x"c4",x"0f",x"00",x"00"),
  1086 => (x"58",x"a6",x"c4",x"86"),
  1087 => (x"9a",x"75",x"4a",x"6e"),
  1088 => (x"c0",x"02",x"aa",x"75"),
  1089 => (x"4a",x"6e",x"87",x"dc"),
  1090 => (x"4a",x"72",x"8a",x"c2"),
  1091 => (x"00",x"1c",x"58",x"27"),
  1092 => (x"27",x"92",x"bf",x"00"),
  1093 => (x"00",x"00",x"1c",x"70"),
  1094 => (x"80",x"72",x"48",x"bf"),
  1095 => (x"fb",x"58",x"a6",x"c8"),
  1096 => (x"48",x"c0",x"87",x"e2"),
  1097 => (x"ff",x"ff",x"ff",x"cf"),
  1098 => (x"86",x"cc",x"4d",x"f8"),
  1099 => (x"4c",x"26",x"4d",x"26"),
  1100 => (x"4a",x"26",x"4b",x"26"),
  1101 => (x"5e",x"0e",x"4f",x"26"),
  1102 => (x"cc",x"0e",x"5b",x"5a"),
  1103 => (x"c1",x"4a",x"bf",x"66"),
  1104 => (x"49",x"66",x"cc",x"82"),
  1105 => (x"4a",x"72",x"79",x"72"),
  1106 => (x"00",x"1c",x"5c",x"27"),
  1107 => (x"72",x"9a",x"bf",x"00"),
  1108 => (x"d3",x"c0",x"05",x"9a"),
  1109 => (x"4a",x"66",x"cc",x"87"),
  1110 => (x"1e",x"6a",x"82",x"c8"),
  1111 => (x"00",x"0f",x"2e",x"27"),
  1112 => (x"86",x"c4",x"0f",x"00"),
  1113 => (x"7a",x"73",x"4b",x"70"),
  1114 => (x"4b",x"26",x"48",x"c1"),
  1115 => (x"4f",x"26",x"4a",x"26"),
  1116 => (x"5b",x"5a",x"5e",x"0e"),
  1117 => (x"1c",x"70",x"27",x"0e"),
  1118 => (x"4a",x"bf",x"00",x"00"),
  1119 => (x"c8",x"4b",x"66",x"cc"),
  1120 => (x"c2",x"4b",x"6b",x"83"),
  1121 => (x"27",x"4b",x"73",x"8b"),
  1122 => (x"00",x"00",x"1c",x"58"),
  1123 => (x"4a",x"72",x"93",x"bf"),
  1124 => (x"5c",x"27",x"82",x"73"),
  1125 => (x"bf",x"00",x"00",x"1c"),
  1126 => (x"bf",x"66",x"cc",x"4b"),
  1127 => (x"73",x"4a",x"72",x"9b"),
  1128 => (x"1e",x"66",x"d0",x"82"),
  1129 => (x"3a",x"27",x"1e",x"72"),
  1130 => (x"0f",x"00",x"00",x"08"),
  1131 => (x"4a",x"70",x"86",x"c8"),
  1132 => (x"c0",x"05",x"9a",x"72"),
  1133 => (x"48",x"c0",x"87",x"c5"),
  1134 => (x"c1",x"87",x"c2",x"c0"),
  1135 => (x"26",x"4b",x"26",x"48"),
  1136 => (x"0e",x"4f",x"26",x"4a"),
  1137 => (x"5c",x"5b",x"5a",x"5e"),
  1138 => (x"66",x"d8",x"0e",x"5d"),
  1139 => (x"1e",x"66",x"d4",x"4c"),
  1140 => (x"00",x"1c",x"90",x"27"),
  1141 => (x"bc",x"27",x"1e",x"00"),
  1142 => (x"0f",x"00",x"00",x"0f"),
  1143 => (x"4a",x"70",x"86",x"c8"),
  1144 => (x"c1",x"02",x"9a",x"72"),
  1145 => (x"94",x"27",x"87",x"df"),
  1146 => (x"bf",x"00",x"00",x"1c"),
  1147 => (x"82",x"ff",x"c7",x"4a"),
  1148 => (x"4d",x"72",x"2a",x"c9"),
  1149 => (x"67",x"27",x"4b",x"c0"),
  1150 => (x"1e",x"00",x"00",x"12"),
  1151 => (x"00",x"00",x"5e",x"27"),
  1152 => (x"86",x"c4",x"0f",x"00"),
  1153 => (x"06",x"ad",x"b7",x"c0"),
  1154 => (x"74",x"87",x"d0",x"c1"),
  1155 => (x"1c",x"90",x"27",x"1e"),
  1156 => (x"27",x"1e",x"00",x"00"),
  1157 => (x"00",x"00",x"11",x"70"),
  1158 => (x"70",x"86",x"c8",x"0f"),
  1159 => (x"05",x"9a",x"72",x"4a"),
  1160 => (x"c0",x"87",x"c5",x"c0"),
  1161 => (x"87",x"f5",x"c0",x"48"),
  1162 => (x"00",x"1c",x"90",x"27"),
  1163 => (x"36",x"27",x"1e",x"00"),
  1164 => (x"0f",x"00",x"00",x"11"),
  1165 => (x"c0",x"c8",x"86",x"c4"),
  1166 => (x"75",x"83",x"c1",x"84"),
  1167 => (x"ff",x"04",x"ab",x"b7"),
  1168 => (x"d6",x"c0",x"87",x"c9"),
  1169 => (x"1e",x"66",x"d4",x"87"),
  1170 => (x"00",x"12",x"80",x"27"),
  1171 => (x"17",x"27",x"1e",x"00"),
  1172 => (x"0f",x"00",x"00",x"01"),
  1173 => (x"48",x"c0",x"86",x"c8"),
  1174 => (x"c1",x"87",x"c2",x"c0"),
  1175 => (x"26",x"4d",x"26",x"48"),
  1176 => (x"26",x"4b",x"26",x"4c"),
  1177 => (x"4f",x"4f",x"26",x"4a"),
  1178 => (x"65",x"6e",x"65",x"70"),
  1179 => (x"69",x"66",x"20",x"64"),
  1180 => (x"20",x"2c",x"65",x"6c"),
  1181 => (x"64",x"61",x"6f",x"6c"),
  1182 => (x"2e",x"67",x"6e",x"69"),
  1183 => (x"00",x"0a",x"2e",x"2e"),
  1184 => (x"27",x"6e",x"61",x"43"),
  1185 => (x"70",x"6f",x"20",x"74"),
  1186 => (x"25",x"20",x"6e",x"65"),
  1187 => (x"0e",x"00",x"0a",x"73"),
  1188 => (x"0e",x"5b",x"5a",x"5e"),
  1189 => (x"d8",x"4a",x"66",x"cc"),
  1190 => (x"9a",x"ff",x"c3",x"2a"),
  1191 => (x"c8",x"4b",x"66",x"cc"),
  1192 => (x"c0",x"fc",x"cf",x"2b"),
  1193 => (x"73",x"4a",x"72",x"9b"),
  1194 => (x"4b",x"66",x"cc",x"b2"),
  1195 => (x"ff",x"c0",x"33",x"c8"),
  1196 => (x"9b",x"c0",x"c0",x"f0"),
  1197 => (x"b2",x"73",x"4a",x"72"),
  1198 => (x"d8",x"4b",x"66",x"cc"),
  1199 => (x"c0",x"c0",x"ff",x"33"),
  1200 => (x"72",x"9b",x"c0",x"c0"),
  1201 => (x"72",x"b2",x"73",x"4a"),
  1202 => (x"26",x"4b",x"26",x"48"),
  1203 => (x"0e",x"4f",x"26",x"4a"),
  1204 => (x"0e",x"5b",x"5a",x"5e"),
  1205 => (x"c8",x"4b",x"66",x"cc"),
  1206 => (x"9b",x"ff",x"c3",x"2b"),
  1207 => (x"4a",x"66",x"cc",x"4b"),
  1208 => (x"fc",x"cf",x"32",x"c8"),
  1209 => (x"4a",x"72",x"9a",x"c0"),
  1210 => (x"72",x"4a",x"b2",x"73"),
  1211 => (x"26",x"4b",x"26",x"48"),
  1212 => (x"0e",x"4f",x"26",x"4a"),
  1213 => (x"0e",x"5b",x"5a",x"5e"),
  1214 => (x"d0",x"4a",x"66",x"cc"),
  1215 => (x"ff",x"ff",x"cf",x"2a"),
  1216 => (x"66",x"cc",x"4a",x"9a"),
  1217 => (x"f0",x"33",x"d0",x"4b"),
  1218 => (x"72",x"9b",x"c0",x"c0"),
  1219 => (x"72",x"b2",x"73",x"4a"),
  1220 => (x"26",x"4b",x"26",x"48"),
  1221 => (x"1e",x"4f",x"26",x"4a"),
  1222 => (x"26",x"87",x"fd",x"ff"),
  1223 => (x"1e",x"72",x"1e",x"4f"),
  1224 => (x"c3",x"4a",x"66",x"cc"),
  1225 => (x"f7",x"c0",x"9a",x"df"),
  1226 => (x"aa",x"b7",x"c0",x"8a"),
  1227 => (x"87",x"c3",x"c0",x"03"),
  1228 => (x"c8",x"82",x"e7",x"c0"),
  1229 => (x"30",x"c4",x"48",x"66"),
  1230 => (x"c8",x"58",x"a6",x"cc"),
  1231 => (x"b0",x"72",x"48",x"66"),
  1232 => (x"c8",x"58",x"a6",x"cc"),
  1233 => (x"4a",x"26",x"48",x"66"),
  1234 => (x"5e",x"0e",x"4f",x"26"),
  1235 => (x"0e",x"5c",x"5b",x"5a"),
  1236 => (x"00",x"1c",x"a0",x"27"),
  1237 => (x"c1",x"48",x"bf",x"00"),
  1238 => (x"1c",x"a4",x"27",x"80"),
  1239 => (x"97",x"58",x"00",x"00"),
  1240 => (x"c1",x"4a",x"66",x"d0"),
  1241 => (x"c0",x"c0",x"c0",x"c0"),
  1242 => (x"b7",x"c0",x"c4",x"92"),
  1243 => (x"d3",x"c1",x"4a",x"92"),
  1244 => (x"c0",x"05",x"aa",x"b7"),
  1245 => (x"a0",x"27",x"87",x"e9"),
  1246 => (x"49",x"00",x"00",x"1c"),
  1247 => (x"a4",x"27",x"79",x"c0"),
  1248 => (x"49",x"00",x"00",x"1c"),
  1249 => (x"ac",x"27",x"79",x"c0"),
  1250 => (x"49",x"00",x"00",x"1c"),
  1251 => (x"b0",x"27",x"79",x"c0"),
  1252 => (x"49",x"00",x"00",x"1c"),
  1253 => (x"c0",x"ff",x"79",x"c0"),
  1254 => (x"79",x"d3",x"c1",x"49"),
  1255 => (x"27",x"87",x"f6",x"c9"),
  1256 => (x"00",x"00",x"1c",x"a0"),
  1257 => (x"b7",x"c1",x"49",x"bf"),
  1258 => (x"db",x"c1",x"05",x"a9"),
  1259 => (x"49",x"c0",x"ff",x"87"),
  1260 => (x"97",x"79",x"f4",x"c1"),
  1261 => (x"c1",x"4a",x"66",x"d0"),
  1262 => (x"c0",x"c0",x"c0",x"c0"),
  1263 => (x"b7",x"c0",x"c4",x"92"),
  1264 => (x"1e",x"72",x"4a",x"92"),
  1265 => (x"00",x"1c",x"b0",x"27"),
  1266 => (x"27",x"1e",x"bf",x"00"),
  1267 => (x"00",x"00",x"13",x"1d"),
  1268 => (x"27",x"86",x"c8",x"0f"),
  1269 => (x"00",x"00",x"1c",x"b4"),
  1270 => (x"1c",x"b0",x"27",x"58"),
  1271 => (x"4c",x"bf",x"00",x"00"),
  1272 => (x"06",x"ac",x"b7",x"c3"),
  1273 => (x"ca",x"87",x"c6",x"c0"),
  1274 => (x"70",x"88",x"74",x"48"),
  1275 => (x"c1",x"4a",x"74",x"4c"),
  1276 => (x"c1",x"48",x"72",x"82"),
  1277 => (x"1c",x"ac",x"27",x"30"),
  1278 => (x"74",x"58",x"00",x"00"),
  1279 => (x"80",x"f0",x"c0",x"48"),
  1280 => (x"70",x"49",x"c0",x"ff"),
  1281 => (x"87",x"cd",x"c8",x"79"),
  1282 => (x"00",x"1c",x"b0",x"27"),
  1283 => (x"c9",x"49",x"bf",x"00"),
  1284 => (x"c7",x"01",x"a9",x"b7"),
  1285 => (x"b0",x"27",x"87",x"ff"),
  1286 => (x"bf",x"00",x"00",x"1c"),
  1287 => (x"a9",x"b7",x"c0",x"49"),
  1288 => (x"87",x"f1",x"c7",x"06"),
  1289 => (x"00",x"1c",x"b0",x"27"),
  1290 => (x"c0",x"48",x"bf",x"00"),
  1291 => (x"c0",x"ff",x"80",x"f0"),
  1292 => (x"27",x"79",x"70",x"49"),
  1293 => (x"00",x"00",x"1c",x"a0"),
  1294 => (x"b7",x"c3",x"49",x"bf"),
  1295 => (x"e9",x"c0",x"01",x"a9"),
  1296 => (x"66",x"d0",x"97",x"87"),
  1297 => (x"c0",x"c0",x"c1",x"4a"),
  1298 => (x"c4",x"92",x"c0",x"c0"),
  1299 => (x"4a",x"92",x"b7",x"c0"),
  1300 => (x"ac",x"27",x"1e",x"72"),
  1301 => (x"bf",x"00",x"00",x"1c"),
  1302 => (x"13",x"1d",x"27",x"1e"),
  1303 => (x"c8",x"0f",x"00",x"00"),
  1304 => (x"1c",x"b0",x"27",x"86"),
  1305 => (x"c6",x"58",x"00",x"00"),
  1306 => (x"a8",x"27",x"87",x"eb"),
  1307 => (x"bf",x"00",x"00",x"1c"),
  1308 => (x"27",x"82",x"c3",x"4a"),
  1309 => (x"00",x"00",x"1c",x"a0"),
  1310 => (x"b7",x"72",x"49",x"bf"),
  1311 => (x"f1",x"c0",x"01",x"a9"),
  1312 => (x"66",x"d0",x"97",x"87"),
  1313 => (x"c0",x"c0",x"c1",x"4a"),
  1314 => (x"c4",x"92",x"c0",x"c0"),
  1315 => (x"4a",x"92",x"b7",x"c0"),
  1316 => (x"a4",x"27",x"1e",x"72"),
  1317 => (x"bf",x"00",x"00",x"1c"),
  1318 => (x"13",x"1d",x"27",x"1e"),
  1319 => (x"c8",x"0f",x"00",x"00"),
  1320 => (x"1c",x"a8",x"27",x"86"),
  1321 => (x"27",x"58",x"00",x"00"),
  1322 => (x"00",x"00",x"1c",x"b4"),
  1323 => (x"c5",x"79",x"c1",x"49"),
  1324 => (x"b0",x"27",x"87",x"e3"),
  1325 => (x"bf",x"00",x"00",x"1c"),
  1326 => (x"a9",x"b7",x"c0",x"49"),
  1327 => (x"87",x"d0",x"c3",x"06"),
  1328 => (x"00",x"1c",x"b0",x"27"),
  1329 => (x"c3",x"49",x"bf",x"00"),
  1330 => (x"c3",x"01",x"a9",x"b7"),
  1331 => (x"ac",x"27",x"87",x"c2"),
  1332 => (x"bf",x"00",x"00",x"1c"),
  1333 => (x"c1",x"32",x"c1",x"4a"),
  1334 => (x"1c",x"a0",x"27",x"82"),
  1335 => (x"49",x"bf",x"00",x"00"),
  1336 => (x"01",x"a9",x"b7",x"72"),
  1337 => (x"97",x"87",x"c2",x"c2"),
  1338 => (x"c1",x"4a",x"66",x"d0"),
  1339 => (x"c0",x"c0",x"c0",x"c0"),
  1340 => (x"b7",x"c0",x"c4",x"92"),
  1341 => (x"1e",x"72",x"4a",x"92"),
  1342 => (x"00",x"1c",x"b8",x"27"),
  1343 => (x"27",x"1e",x"bf",x"00"),
  1344 => (x"00",x"00",x"13",x"1d"),
  1345 => (x"27",x"86",x"c8",x"0f"),
  1346 => (x"00",x"00",x"1c",x"bc"),
  1347 => (x"1c",x"b4",x"27",x"58"),
  1348 => (x"4a",x"bf",x"00",x"00"),
  1349 => (x"b4",x"27",x"8a",x"c1"),
  1350 => (x"49",x"00",x"00",x"1c"),
  1351 => (x"b7",x"c0",x"79",x"72"),
  1352 => (x"f0",x"c3",x"03",x"aa"),
  1353 => (x"1c",x"a4",x"27",x"87"),
  1354 => (x"4a",x"bf",x"00",x"00"),
  1355 => (x"00",x"1c",x"b8",x"27"),
  1356 => (x"52",x"bf",x"97",x"00"),
  1357 => (x"00",x"1c",x"a4",x"27"),
  1358 => (x"c1",x"4a",x"bf",x"00"),
  1359 => (x"1c",x"a4",x"27",x"82"),
  1360 => (x"72",x"49",x"00",x"00"),
  1361 => (x"1c",x"bc",x"27",x"79"),
  1362 => (x"b7",x"bf",x"00",x"00"),
  1363 => (x"cd",x"c0",x"06",x"aa"),
  1364 => (x"1c",x"bc",x"27",x"87"),
  1365 => (x"27",x"49",x"00",x"00"),
  1366 => (x"00",x"00",x"1c",x"a4"),
  1367 => (x"b4",x"27",x"79",x"bf"),
  1368 => (x"49",x"00",x"00",x"1c"),
  1369 => (x"ec",x"c2",x"79",x"c1"),
  1370 => (x"1c",x"b4",x"27",x"87"),
  1371 => (x"05",x"bf",x"00",x"00"),
  1372 => (x"27",x"87",x"e2",x"c2"),
  1373 => (x"00",x"00",x"1c",x"b8"),
  1374 => (x"33",x"c4",x"4b",x"bf"),
  1375 => (x"00",x"1c",x"b8",x"27"),
  1376 => (x"79",x"73",x"49",x"00"),
  1377 => (x"00",x"1c",x"a4",x"27"),
  1378 => (x"73",x"4a",x"bf",x"00"),
  1379 => (x"87",x"c5",x"c2",x"52"),
  1380 => (x"00",x"1c",x"b0",x"27"),
  1381 => (x"c7",x"49",x"bf",x"00"),
  1382 => (x"c1",x"04",x"a9",x"b7"),
  1383 => (x"4b",x"c0",x"87",x"e8"),
  1384 => (x"c1",x"49",x"f4",x"fe"),
  1385 => (x"1c",x"a4",x"27",x"79"),
  1386 => (x"c0",x"49",x"00",x"00"),
  1387 => (x"1c",x"bc",x"27",x"79"),
  1388 => (x"49",x"bf",x"00",x"00"),
  1389 => (x"06",x"a9",x"b7",x"c0"),
  1390 => (x"27",x"87",x"e5",x"c0"),
  1391 => (x"00",x"00",x"1c",x"a4"),
  1392 => (x"27",x"83",x"bf",x"bf"),
  1393 => (x"00",x"00",x"1c",x"a4"),
  1394 => (x"82",x"c4",x"4a",x"bf"),
  1395 => (x"00",x"1c",x"a4",x"27"),
  1396 => (x"79",x"72",x"49",x"00"),
  1397 => (x"00",x"1c",x"bc",x"27"),
  1398 => (x"aa",x"b7",x"bf",x"00"),
  1399 => (x"87",x"db",x"ff",x"04"),
  1400 => (x"bc",x"27",x"1e",x"73"),
  1401 => (x"bf",x"00",x"00",x"1c"),
  1402 => (x"19",x"a4",x"27",x"1e"),
  1403 => (x"27",x"1e",x"00",x"00"),
  1404 => (x"00",x"00",x"01",x"17"),
  1405 => (x"ff",x"86",x"cc",x"0f"),
  1406 => (x"c2",x"c1",x"49",x"c0"),
  1407 => (x"13",x"17",x"27",x"79"),
  1408 => (x"c0",x"0f",x"00",x"00"),
  1409 => (x"b0",x"27",x"87",x"cf"),
  1410 => (x"bf",x"00",x"00",x"1c"),
  1411 => (x"80",x"f0",x"c0",x"48"),
  1412 => (x"70",x"49",x"c0",x"ff"),
  1413 => (x"26",x"4c",x"26",x"79"),
  1414 => (x"26",x"4a",x"26",x"4b"),
  1415 => (x"fd",x"ff",x"1e",x"4f"),
  1416 => (x"0e",x"4f",x"26",x"87"),
  1417 => (x"5c",x"5b",x"5a",x"5e"),
  1418 => (x"0b",x"27",x"0e",x"5d"),
  1419 => (x"1e",x"00",x"00",x"18"),
  1420 => (x"00",x"00",x"5e",x"27"),
  1421 => (x"86",x"c4",x"0f",x"00"),
  1422 => (x"00",x"05",x"43",x"27"),
  1423 => (x"4a",x"70",x"0f",x"00"),
  1424 => (x"c4",x"02",x"9a",x"72"),
  1425 => (x"e8",x"27",x"87",x"ce"),
  1426 => (x"1e",x"00",x"00",x"17"),
  1427 => (x"00",x"00",x"5e",x"27"),
  1428 => (x"86",x"c4",x"0f",x"00"),
  1429 => (x"00",x"0b",x"04",x"27"),
  1430 => (x"c0",x"27",x"0f",x"00"),
  1431 => (x"1e",x"00",x"00",x"1c"),
  1432 => (x"00",x"17",x"ff",x"27"),
  1433 => (x"c3",x"27",x"1e",x"00"),
  1434 => (x"0f",x"00",x"00",x"11"),
  1435 => (x"4a",x"70",x"86",x"c8"),
  1436 => (x"c3",x"02",x"9a",x"72"),
  1437 => (x"c0",x"27",x"87",x"d0"),
  1438 => (x"4b",x"00",x"00",x"1c"),
  1439 => (x"00",x"17",x"bd",x"27"),
  1440 => (x"5e",x"27",x"1e",x"00"),
  1441 => (x"0f",x"00",x"00",x"00"),
  1442 => (x"4d",x"c0",x"86",x"c4"),
  1443 => (x"4a",x"74",x"4c",x"13"),
  1444 => (x"aa",x"b7",x"e0",x"c0"),
  1445 => (x"87",x"ed",x"c1",x"02"),
  1446 => (x"c0",x"ff",x"48",x"74"),
  1447 => (x"74",x"79",x"70",x"49"),
  1448 => (x"b7",x"e3",x"c0",x"4a"),
  1449 => (x"dc",x"c1",x"02",x"aa"),
  1450 => (x"c1",x"4a",x"74",x"87"),
  1451 => (x"05",x"aa",x"b7",x"c7"),
  1452 => (x"27",x"87",x"c6",x"c0"),
  1453 => (x"00",x"00",x"13",x"17"),
  1454 => (x"ca",x"4a",x"74",x"0f"),
  1455 => (x"c0",x"05",x"aa",x"b7"),
  1456 => (x"1d",x"27",x"87",x"c6"),
  1457 => (x"0f",x"00",x"00",x"16"),
  1458 => (x"cc",x"c1",x"4a",x"74"),
  1459 => (x"c0",x"05",x"aa",x"b7"),
  1460 => (x"c0",x"27",x"87",x"c6"),
  1461 => (x"4b",x"00",x"00",x"1c"),
  1462 => (x"df",x"ff",x"4a",x"74"),
  1463 => (x"72",x"8a",x"d0",x"9a"),
  1464 => (x"c0",x"4a",x"74",x"4c"),
  1465 => (x"04",x"aa",x"b7",x"f9"),
  1466 => (x"74",x"87",x"c6",x"c0"),
  1467 => (x"72",x"8a",x"d1",x"4a"),
  1468 => (x"74",x"35",x"c4",x"4c"),
  1469 => (x"72",x"4d",x"75",x"4a"),
  1470 => (x"74",x"4c",x"13",x"b5"),
  1471 => (x"b7",x"e0",x"c0",x"4a"),
  1472 => (x"d3",x"fe",x"05",x"aa"),
  1473 => (x"c0",x"4a",x"74",x"87"),
  1474 => (x"02",x"aa",x"b7",x"e3"),
  1475 => (x"13",x"87",x"e2",x"c0"),
  1476 => (x"b7",x"e0",x"c0",x"4a"),
  1477 => (x"ca",x"c0",x"05",x"aa"),
  1478 => (x"c0",x"4a",x"13",x"87"),
  1479 => (x"02",x"aa",x"b7",x"e0"),
  1480 => (x"c1",x"87",x"f6",x"ff"),
  1481 => (x"73",x"1e",x"75",x"8b"),
  1482 => (x"11",x"c3",x"27",x"1e"),
  1483 => (x"c8",x"0f",x"00",x"00"),
  1484 => (x"ca",x"4a",x"13",x"86"),
  1485 => (x"fd",x"02",x"aa",x"b7"),
  1486 => (x"4a",x"13",x"87",x"d0"),
  1487 => (x"05",x"aa",x"b7",x"ca"),
  1488 => (x"fd",x"87",x"f7",x"ff"),
  1489 => (x"cf",x"27",x"87",x"c4"),
  1490 => (x"1e",x"00",x"00",x"17"),
  1491 => (x"00",x"00",x"5e",x"27"),
  1492 => (x"86",x"c4",x"0f",x"00"),
  1493 => (x"00",x"18",x"21",x"27"),
  1494 => (x"5e",x"27",x"1e",x"00"),
  1495 => (x"0f",x"00",x"00",x"00"),
  1496 => (x"bc",x"27",x"86",x"c4"),
  1497 => (x"49",x"00",x"00",x"1c"),
  1498 => (x"f4",x"c3",x"79",x"c0"),
  1499 => (x"c0",x"4d",x"ff",x"c8"),
  1500 => (x"3f",x"27",x"1e",x"ee"),
  1501 => (x"0f",x"00",x"00",x"00"),
  1502 => (x"4b",x"75",x"86",x"c4"),
  1503 => (x"c0",x"c9",x"f4",x"c3"),
  1504 => (x"bf",x"c0",x"ff",x"4d"),
  1505 => (x"c8",x"4a",x"74",x"4c"),
  1506 => (x"9a",x"72",x"9a",x"c0"),
  1507 => (x"87",x"d1",x"c0",x"02"),
  1508 => (x"ff",x"c3",x"4a",x"74"),
  1509 => (x"27",x"1e",x"72",x"9a"),
  1510 => (x"00",x"00",x"13",x"4a"),
  1511 => (x"75",x"86",x"c4",x"0f"),
  1512 => (x"c1",x"4a",x"73",x"4b"),
  1513 => (x"05",x"9a",x"72",x"8b"),
  1514 => (x"c3",x"87",x"d6",x"ff"),
  1515 => (x"4d",x"ff",x"c8",x"f4"),
  1516 => (x"26",x"87",x"fc",x"fe"),
  1517 => (x"26",x"4c",x"26",x"4d"),
  1518 => (x"26",x"4a",x"26",x"4b"),
  1519 => (x"72",x"61",x"50",x"4f"),
  1520 => (x"67",x"6e",x"69",x"73"),
  1521 => (x"6e",x"61",x"6d",x"20"),
  1522 => (x"73",x"65",x"66",x"69"),
  1523 => (x"4c",x"00",x"0a",x"74"),
  1524 => (x"69",x"64",x"61",x"6f"),
  1525 => (x"6d",x"20",x"67",x"6e"),
  1526 => (x"66",x"69",x"6e",x"61"),
  1527 => (x"20",x"74",x"73",x"65"),
  1528 => (x"6c",x"69",x"61",x"66"),
  1529 => (x"00",x"0a",x"64",x"65"),
  1530 => (x"74",x"6e",x"75",x"48"),
  1531 => (x"20",x"67",x"6e",x"69"),
  1532 => (x"20",x"72",x"6f",x"66"),
  1533 => (x"74",x"72",x"61",x"70"),
  1534 => (x"6f",x"69",x"74",x"69"),
  1535 => (x"4d",x"00",x"0a",x"6e"),
  1536 => (x"46",x"49",x"4e",x"41"),
  1537 => (x"4d",x"54",x"53",x"45"),
  1538 => (x"49",x"00",x"54",x"53"),
  1539 => (x"69",x"74",x"69",x"6e"),
  1540 => (x"7a",x"69",x"6c",x"61"),
  1541 => (x"20",x"67",x"6e",x"69"),
  1542 => (x"63",x"20",x"44",x"53"),
  1543 => (x"0a",x"64",x"72",x"61"),
  1544 => (x"6f",x"6f",x"42",x"00"),
  1545 => (x"67",x"6e",x"69",x"74"),
  1546 => (x"6f",x"72",x"66",x"20"),
  1547 => (x"53",x"52",x"20",x"6d"),
  1548 => (x"2e",x"32",x"33",x"32"),
  1549 => (x"44",x"4d",x"43",x"00"),
  1550 => (x"61",x"65",x"52",x"00"),
  1551 => (x"66",x"6f",x"20",x"64"),
  1552 => (x"52",x"42",x"4d",x"20"),
  1553 => (x"69",x"61",x"66",x"20"),
  1554 => (x"0a",x"64",x"65",x"6c"),
  1555 => (x"20",x"6f",x"4e",x"00"),
  1556 => (x"74",x"72",x"61",x"70"),
  1557 => (x"6f",x"69",x"74",x"69"),
  1558 => (x"69",x"73",x"20",x"6e"),
  1559 => (x"74",x"61",x"6e",x"67"),
  1560 => (x"20",x"65",x"72",x"75"),
  1561 => (x"6e",x"75",x"6f",x"66"),
  1562 => (x"4d",x"00",x"0a",x"64"),
  1563 => (x"69",x"73",x"52",x"42"),
  1564 => (x"20",x"3a",x"65",x"7a"),
  1565 => (x"20",x"2c",x"64",x"25"),
  1566 => (x"74",x"72",x"61",x"70"),
  1567 => (x"6f",x"69",x"74",x"69"),
  1568 => (x"7a",x"69",x"73",x"6e"),
  1569 => (x"25",x"20",x"3a",x"65"),
  1570 => (x"6f",x"20",x"2c",x"64"),
  1571 => (x"65",x"73",x"66",x"66"),
  1572 => (x"66",x"6f",x"20",x"74"),
  1573 => (x"67",x"69",x"73",x"20"),
  1574 => (x"64",x"25",x"20",x"3a"),
  1575 => (x"69",x"73",x"20",x"2c"),
  1576 => (x"78",x"30",x"20",x"67"),
  1577 => (x"00",x"0a",x"78",x"25"),
  1578 => (x"64",x"61",x"65",x"52"),
  1579 => (x"20",x"67",x"6e",x"69"),
  1580 => (x"74",x"6f",x"6f",x"62"),
  1581 => (x"63",x"65",x"73",x"20"),
  1582 => (x"20",x"72",x"6f",x"74"),
  1583 => (x"00",x"0a",x"64",x"25"),
  1584 => (x"64",x"61",x"65",x"52"),
  1585 => (x"6f",x"6f",x"62",x"20"),
  1586 => (x"65",x"73",x"20",x"74"),
  1587 => (x"72",x"6f",x"74",x"63"),
  1588 => (x"6f",x"72",x"66",x"20"),
  1589 => (x"69",x"66",x"20",x"6d"),
  1590 => (x"20",x"74",x"73",x"72"),
  1591 => (x"74",x"72",x"61",x"70"),
  1592 => (x"6f",x"69",x"74",x"69"),
  1593 => (x"55",x"00",x"0a",x"6e"),
  1594 => (x"70",x"75",x"73",x"6e"),
  1595 => (x"74",x"72",x"6f",x"70"),
  1596 => (x"70",x"20",x"64",x"65"),
  1597 => (x"69",x"74",x"72",x"61"),
  1598 => (x"6e",x"6f",x"69",x"74"),
  1599 => (x"70",x"79",x"74",x"20"),
  1600 => (x"00",x"0d",x"21",x"65"),
  1601 => (x"33",x"54",x"41",x"46"),
  1602 => (x"20",x"20",x"20",x"32"),
  1603 => (x"61",x"65",x"52",x"00"),
  1604 => (x"67",x"6e",x"69",x"64"),
  1605 => (x"52",x"42",x"4d",x"20"),
  1606 => (x"42",x"4d",x"00",x"0a"),
  1607 => (x"75",x"73",x"20",x"52"),
  1608 => (x"73",x"65",x"63",x"63"),
  1609 => (x"6c",x"75",x"66",x"73"),
  1610 => (x"72",x"20",x"79",x"6c"),
  1611 => (x"0a",x"64",x"61",x"65"),
  1612 => (x"54",x"41",x"46",x"00"),
  1613 => (x"20",x"20",x"36",x"31"),
  1614 => (x"41",x"46",x"00",x"20"),
  1615 => (x"20",x"32",x"33",x"54"),
  1616 => (x"50",x"00",x"20",x"20"),
  1617 => (x"69",x"74",x"72",x"61"),
  1618 => (x"6e",x"6f",x"69",x"74"),
  1619 => (x"6e",x"75",x"6f",x"63"),
  1620 => (x"64",x"25",x"20",x"74"),
  1621 => (x"75",x"48",x"00",x"0a"),
  1622 => (x"6e",x"69",x"74",x"6e"),
  1623 => (x"6f",x"66",x"20",x"67"),
  1624 => (x"69",x"66",x"20",x"72"),
  1625 => (x"79",x"73",x"65",x"6c"),
  1626 => (x"6d",x"65",x"74",x"73"),
  1627 => (x"41",x"46",x"00",x"0a"),
  1628 => (x"20",x"32",x"33",x"54"),
  1629 => (x"46",x"00",x"20",x"20"),
  1630 => (x"36",x"31",x"54",x"41"),
  1631 => (x"00",x"20",x"20",x"20"),
  1632 => (x"73",x"75",x"6c",x"43"),
  1633 => (x"20",x"72",x"65",x"74"),
  1634 => (x"65",x"7a",x"69",x"73"),
  1635 => (x"64",x"25",x"20",x"3a"),
  1636 => (x"6c",x"43",x"20",x"2c"),
  1637 => (x"65",x"74",x"73",x"75"),
  1638 => (x"61",x"6d",x"20",x"72"),
  1639 => (x"20",x"2c",x"6b",x"73"),
  1640 => (x"00",x"0a",x"64",x"25"),
  1641 => (x"63",x"65",x"68",x"43"),
  1642 => (x"6d",x"75",x"73",x"6b"),
  1643 => (x"20",x"6f",x"74",x"20"),
  1644 => (x"20",x"3a",x"64",x"25"),
  1645 => (x"00",x"0a",x"64",x"25"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
