
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of OSDBoot_832_ROM is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"3b",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"38"),
    10 => (x"20",x"00",x"27",x"4f"),
    11 => (x"27",x"4e",x"00",x"00"),
    12 => (x"00",x"00",x"04",x"80"),
    13 => (x"87",x"fd",x"00",x"0f"),
    14 => (x"4f",x"87",x"fd",x"00"),
    15 => (x"5c",x"5b",x"5e",x"0e"),
    16 => (x"86",x"f0",x"0e",x"5d"),
    17 => (x"a6",x"c4",x"4c",x"c0"),
    18 => (x"c0",x"78",x"c0",x"48"),
    19 => (x"c0",x"4b",x"a6",x"e4"),
    20 => (x"48",x"49",x"66",x"e0"),
    21 => (x"e4",x"c0",x"80",x"c1"),
    22 => (x"4d",x"11",x"58",x"a6"),
    23 => (x"bd",x"85",x"c0",x"fe"),
    24 => (x"c4",x"02",x"9d",x"75"),
    25 => (x"66",x"c4",x"87",x"d3"),
    26 => (x"87",x"e1",x"c3",x"02"),
    27 => (x"c0",x"48",x"a6",x"c4"),
    28 => (x"c0",x"49",x"75",x"78"),
    29 => (x"c2",x"02",x"ad",x"f0"),
    30 => (x"e3",x"c1",x"87",x"ef"),
    31 => (x"f0",x"c2",x"02",x"a9"),
    32 => (x"a9",x"e4",x"c1",x"87"),
    33 => (x"87",x"e1",x"c0",x"02"),
    34 => (x"02",x"a9",x"ec",x"c1"),
    35 => (x"c1",x"87",x"da",x"c2"),
    36 => (x"d4",x"02",x"a9",x"f0"),
    37 => (x"a9",x"f3",x"c1",x"87"),
    38 => (x"87",x"f8",x"c1",x"02"),
    39 => (x"02",x"a9",x"f5",x"c1"),
    40 => (x"f8",x"c1",x"87",x"c7"),
    41 => (x"da",x"c2",x"05",x"a9"),
    42 => (x"73",x"83",x"c4",x"87"),
    43 => (x"76",x"89",x"c4",x"49"),
    44 => (x"6e",x"78",x"69",x"48"),
    45 => (x"87",x"ce",x"c1",x"02"),
    46 => (x"78",x"c0",x"80",x"c8"),
    47 => (x"c0",x"48",x"a6",x"cc"),
    48 => (x"4d",x"66",x"cc",x"78"),
    49 => (x"b7",x"dc",x"49",x"6e"),
    50 => (x"cf",x"4a",x"71",x"29"),
    51 => (x"c4",x"48",x"6e",x"9a"),
    52 => (x"58",x"a6",x"c4",x"30"),
    53 => (x"c5",x"02",x"9a",x"72"),
    54 => (x"48",x"a6",x"c8",x"87"),
    55 => (x"aa",x"c9",x"78",x"c1"),
    56 => (x"c0",x"87",x"c5",x"06"),
    57 => (x"87",x"c3",x"82",x"f7"),
    58 => (x"c8",x"82",x"f0",x"c0"),
    59 => (x"87",x"ca",x"02",x"66"),
    60 => (x"cf",x"c1",x"1e",x"72"),
    61 => (x"86",x"c4",x"87",x"ec"),
    62 => (x"85",x"c1",x"84",x"c1"),
    63 => (x"04",x"ad",x"b7",x"c8"),
    64 => (x"c1",x"87",x"c1",x"ff"),
    65 => (x"f0",x"c0",x"87",x"dc"),
    66 => (x"d5",x"cf",x"c1",x"1e"),
    67 => (x"c1",x"86",x"c4",x"87"),
    68 => (x"87",x"ce",x"c1",x"84"),
    69 => (x"49",x"73",x"83",x"c4"),
    70 => (x"1e",x"69",x"89",x"c4"),
    71 => (x"87",x"eb",x"cf",x"c1"),
    72 => (x"49",x"70",x"86",x"c4"),
    73 => (x"f9",x"c0",x"84",x"71"),
    74 => (x"48",x"a6",x"c4",x"87"),
    75 => (x"f1",x"c0",x"78",x"c1"),
    76 => (x"73",x"83",x"c4",x"87"),
    77 => (x"69",x"89",x"c4",x"49"),
    78 => (x"e5",x"ce",x"c1",x"1e"),
    79 => (x"c1",x"86",x"c4",x"87"),
    80 => (x"75",x"87",x"df",x"84"),
    81 => (x"d9",x"ce",x"c1",x"1e"),
    82 => (x"d5",x"86",x"c4",x"87"),
    83 => (x"ad",x"e5",x"c0",x"87"),
    84 => (x"c4",x"87",x"c7",x"05"),
    85 => (x"78",x"c1",x"48",x"a6"),
    86 => (x"1e",x"75",x"87",x"c8"),
    87 => (x"87",x"c2",x"ce",x"c1"),
    88 => (x"e0",x"c0",x"86",x"c4"),
    89 => (x"c1",x"48",x"49",x"66"),
    90 => (x"a6",x"e4",x"c0",x"80"),
    91 => (x"fe",x"4d",x"11",x"58"),
    92 => (x"75",x"bd",x"85",x"c0"),
    93 => (x"ed",x"fb",x"05",x"9d"),
    94 => (x"f0",x"48",x"74",x"87"),
    95 => (x"26",x"4d",x"26",x"8e"),
    96 => (x"26",x"4b",x"26",x"4c"),
    97 => (x"0e",x"5e",x"0e",x"4f"),
    98 => (x"d8",x"49",x"66",x"c4"),
    99 => (x"99",x"ff",x"c3",x"29"),
   100 => (x"c8",x"4a",x"66",x"c4"),
   101 => (x"c0",x"fc",x"cf",x"2a"),
   102 => (x"c4",x"b1",x"72",x"9a"),
   103 => (x"32",x"c8",x"4a",x"66"),
   104 => (x"c0",x"f0",x"ff",x"c0"),
   105 => (x"b1",x"72",x"9a",x"c0"),
   106 => (x"d8",x"4a",x"66",x"c4"),
   107 => (x"c0",x"fc",x"cf",x"32"),
   108 => (x"72",x"9a",x"c0",x"c0"),
   109 => (x"26",x"48",x"71",x"b1"),
   110 => (x"0e",x"5e",x"0e",x"4f"),
   111 => (x"c8",x"49",x"66",x"c4"),
   112 => (x"99",x"ff",x"c3",x"29"),
   113 => (x"c8",x"4a",x"66",x"c4"),
   114 => (x"c0",x"fc",x"cf",x"32"),
   115 => (x"71",x"b1",x"72",x"9a"),
   116 => (x"0e",x"4f",x"26",x"48"),
   117 => (x"66",x"c4",x"0e",x"5e"),
   118 => (x"cf",x"29",x"d0",x"49"),
   119 => (x"c4",x"99",x"ff",x"ff"),
   120 => (x"32",x"d0",x"4a",x"66"),
   121 => (x"9a",x"c0",x"c0",x"f0"),
   122 => (x"48",x"71",x"b1",x"72"),
   123 => (x"cf",x"1e",x"4f",x"26"),
   124 => (x"cb",x"f8",x"ff",x"ff"),
   125 => (x"26",x"87",x"fe",x"87"),
   126 => (x"66",x"c8",x"1e",x"4f"),
   127 => (x"99",x"df",x"c3",x"49"),
   128 => (x"c0",x"89",x"f7",x"c0"),
   129 => (x"c3",x"03",x"a9",x"b7"),
   130 => (x"81",x"e7",x"c0",x"87"),
   131 => (x"c4",x"48",x"66",x"c4"),
   132 => (x"58",x"a6",x"c8",x"30"),
   133 => (x"71",x"48",x"66",x"c4"),
   134 => (x"58",x"a6",x"c8",x"b0"),
   135 => (x"26",x"48",x"66",x"c4"),
   136 => (x"5b",x"5e",x"0e",x"4f"),
   137 => (x"f6",x"c0",x"0e",x"5c"),
   138 => (x"4b",x"c0",x"c0",x"e8"),
   139 => (x"bf",x"c8",x"d7",x"c1"),
   140 => (x"c1",x"80",x"c1",x"48"),
   141 => (x"97",x"58",x"cc",x"d7"),
   142 => (x"fe",x"49",x"66",x"cc"),
   143 => (x"c1",x"b9",x"81",x"c0"),
   144 => (x"de",x"05",x"a9",x"d3"),
   145 => (x"c8",x"d7",x"c1",x"87"),
   146 => (x"c1",x"78",x"c0",x"48"),
   147 => (x"c0",x"48",x"cc",x"d7"),
   148 => (x"d4",x"d7",x"c1",x"78"),
   149 => (x"c1",x"78",x"c0",x"48"),
   150 => (x"c0",x"48",x"d8",x"d7"),
   151 => (x"7b",x"d3",x"c1",x"78"),
   152 => (x"c1",x"87",x"d6",x"c7"),
   153 => (x"48",x"bf",x"c8",x"d7"),
   154 => (x"c1",x"05",x"a8",x"c1"),
   155 => (x"f4",x"c1",x"87",x"c2"),
   156 => (x"66",x"cc",x"97",x"7b"),
   157 => (x"81",x"c0",x"fe",x"49"),
   158 => (x"c1",x"1e",x"71",x"b9"),
   159 => (x"1e",x"bf",x"d8",x"d7"),
   160 => (x"c8",x"87",x"f6",x"fd"),
   161 => (x"dc",x"d7",x"c1",x"86"),
   162 => (x"d8",x"d7",x"c1",x"58"),
   163 => (x"b7",x"c3",x"4c",x"bf"),
   164 => (x"87",x"c6",x"06",x"ac"),
   165 => (x"88",x"74",x"48",x"ca"),
   166 => (x"49",x"74",x"4c",x"70"),
   167 => (x"48",x"71",x"81",x"c1"),
   168 => (x"d7",x"c1",x"30",x"c1"),
   169 => (x"48",x"74",x"58",x"d4"),
   170 => (x"70",x"80",x"f0",x"c0"),
   171 => (x"87",x"c9",x"c6",x"7b"),
   172 => (x"bf",x"d8",x"d7",x"c1"),
   173 => (x"a8",x"b7",x"c9",x"48"),
   174 => (x"87",x"fd",x"c5",x"01"),
   175 => (x"bf",x"d8",x"d7",x"c1"),
   176 => (x"a8",x"b7",x"c0",x"48"),
   177 => (x"87",x"f1",x"c5",x"06"),
   178 => (x"bf",x"d8",x"d7",x"c1"),
   179 => (x"80",x"f0",x"c0",x"48"),
   180 => (x"d7",x"c1",x"7b",x"70"),
   181 => (x"c3",x"48",x"bf",x"c8"),
   182 => (x"db",x"01",x"a8",x"b7"),
   183 => (x"66",x"cc",x"97",x"87"),
   184 => (x"81",x"c0",x"fe",x"49"),
   185 => (x"c1",x"1e",x"71",x"b9"),
   186 => (x"1e",x"bf",x"d4",x"d7"),
   187 => (x"c8",x"87",x"ca",x"fc"),
   188 => (x"d8",x"d7",x"c1",x"86"),
   189 => (x"87",x"c1",x"c5",x"58"),
   190 => (x"bf",x"d0",x"d7",x"c1"),
   191 => (x"c1",x"81",x"c3",x"49"),
   192 => (x"b7",x"bf",x"c8",x"d7"),
   193 => (x"e1",x"c0",x"04",x"a9"),
   194 => (x"66",x"cc",x"97",x"87"),
   195 => (x"81",x"c0",x"fe",x"49"),
   196 => (x"c1",x"1e",x"71",x"b9"),
   197 => (x"1e",x"bf",x"cc",x"d7"),
   198 => (x"c8",x"87",x"de",x"fb"),
   199 => (x"d0",x"d7",x"c1",x"86"),
   200 => (x"dc",x"d7",x"c1",x"58"),
   201 => (x"c4",x"78",x"c1",x"48"),
   202 => (x"d7",x"c1",x"87",x"cf"),
   203 => (x"c0",x"48",x"bf",x"d8"),
   204 => (x"c2",x"06",x"a8",x"b7"),
   205 => (x"d7",x"c1",x"87",x"db"),
   206 => (x"c3",x"48",x"bf",x"d8"),
   207 => (x"c2",x"01",x"a8",x"b7"),
   208 => (x"d7",x"c1",x"87",x"cf"),
   209 => (x"c1",x"49",x"bf",x"d4"),
   210 => (x"d7",x"c1",x"81",x"31"),
   211 => (x"a9",x"b7",x"bf",x"c8"),
   212 => (x"87",x"df",x"c1",x"04"),
   213 => (x"49",x"66",x"cc",x"97"),
   214 => (x"b9",x"81",x"c0",x"fe"),
   215 => (x"d7",x"c1",x"1e",x"71"),
   216 => (x"fa",x"1e",x"bf",x"e0"),
   217 => (x"86",x"c8",x"87",x"d3"),
   218 => (x"58",x"e4",x"d7",x"c1"),
   219 => (x"bf",x"dc",x"d7",x"c1"),
   220 => (x"c1",x"89",x"c1",x"49"),
   221 => (x"c0",x"59",x"e0",x"d7"),
   222 => (x"c2",x"03",x"a9",x"b7"),
   223 => (x"d7",x"c1",x"87",x"fb"),
   224 => (x"c1",x"49",x"bf",x"cc"),
   225 => (x"bf",x"97",x"e0",x"d7"),
   226 => (x"98",x"ff",x"c3",x"51"),
   227 => (x"bf",x"cc",x"d7",x"c1"),
   228 => (x"c1",x"81",x"c1",x"49"),
   229 => (x"c1",x"59",x"d0",x"d7"),
   230 => (x"b7",x"bf",x"e4",x"d7"),
   231 => (x"c9",x"c0",x"06",x"a9"),
   232 => (x"e4",x"d7",x"c1",x"87"),
   233 => (x"cc",x"d7",x"c1",x"48"),
   234 => (x"d7",x"c1",x"78",x"bf"),
   235 => (x"78",x"c1",x"48",x"dc"),
   236 => (x"c1",x"87",x"c6",x"c2"),
   237 => (x"05",x"bf",x"dc",x"d7"),
   238 => (x"c1",x"87",x"fe",x"c1"),
   239 => (x"49",x"bf",x"e0",x"d7"),
   240 => (x"d7",x"c1",x"31",x"c4"),
   241 => (x"d7",x"c1",x"59",x"e4"),
   242 => (x"97",x"09",x"bf",x"cc"),
   243 => (x"e8",x"c1",x"09",x"79"),
   244 => (x"d8",x"d7",x"c1",x"87"),
   245 => (x"b7",x"c7",x"48",x"bf"),
   246 => (x"d2",x"c1",x"04",x"a8"),
   247 => (x"fe",x"4a",x"c0",x"87"),
   248 => (x"78",x"c1",x"48",x"f4"),
   249 => (x"48",x"cc",x"d7",x"c1"),
   250 => (x"c0",x"c0",x"c0",x"d0"),
   251 => (x"c1",x"48",x"78",x"c0"),
   252 => (x"b7",x"bf",x"e4",x"d7"),
   253 => (x"db",x"c0",x"03",x"a8"),
   254 => (x"cc",x"d7",x"c1",x"87"),
   255 => (x"c1",x"82",x"bf",x"bf"),
   256 => (x"49",x"bf",x"cc",x"d7"),
   257 => (x"d7",x"c1",x"81",x"c4"),
   258 => (x"d7",x"c1",x"59",x"d0"),
   259 => (x"a9",x"b7",x"bf",x"e4"),
   260 => (x"87",x"e5",x"ff",x"04"),
   261 => (x"d7",x"c1",x"1e",x"72"),
   262 => (x"d9",x"1e",x"bf",x"e4"),
   263 => (x"db",x"f0",x"1e",x"e3"),
   264 => (x"c1",x"86",x"cc",x"87"),
   265 => (x"ff",x"cf",x"7b",x"c2"),
   266 => (x"87",x"d4",x"ef",x"ff"),
   267 => (x"c1",x"87",x"ca",x"c0"),
   268 => (x"48",x"bf",x"d8",x"d7"),
   269 => (x"70",x"80",x"f0",x"c0"),
   270 => (x"26",x"4c",x"26",x"7b"),
   271 => (x"0e",x"4f",x"26",x"4b"),
   272 => (x"5d",x"5c",x"5b",x"5e"),
   273 => (x"4d",x"66",x"d0",x"0e"),
   274 => (x"c0",x"4c",x"66",x"d4"),
   275 => (x"dc",x"49",x"75",x"4b"),
   276 => (x"4a",x"71",x"29",x"b7"),
   277 => (x"35",x"c4",x"9a",x"cf"),
   278 => (x"06",x"aa",x"b7",x"c9"),
   279 => (x"c0",x"87",x"c6",x"c0"),
   280 => (x"c3",x"c0",x"82",x"f7"),
   281 => (x"82",x"f0",x"c0",x"87"),
   282 => (x"c3",x"7c",x"97",x"72"),
   283 => (x"84",x"c1",x"98",x"ff"),
   284 => (x"ab",x"b7",x"c8",x"83"),
   285 => (x"87",x"d5",x"ff",x"04"),
   286 => (x"4c",x"26",x"4d",x"26"),
   287 => (x"4f",x"26",x"4b",x"26"),
   288 => (x"5c",x"5b",x"5e",x"0e"),
   289 => (x"86",x"f0",x"0e",x"5d"),
   290 => (x"c1",x"1e",x"f9",x"d8"),
   291 => (x"c4",x"87",x"fc",x"c1"),
   292 => (x"d0",x"fb",x"c0",x"86"),
   293 => (x"02",x"98",x"70",x"87"),
   294 => (x"d8",x"87",x"f2",x"c3"),
   295 => (x"c1",x"c1",x"1e",x"e2"),
   296 => (x"86",x"c4",x"87",x"e9"),
   297 => (x"70",x"87",x"d0",x"c8"),
   298 => (x"d7",x"c3",x"02",x"98"),
   299 => (x"c0",x"c0",x"d0",x"87"),
   300 => (x"d7",x"1e",x"c0",x"c0"),
   301 => (x"ff",x"dc",x"1e",x"fa"),
   302 => (x"70",x"86",x"c8",x"87"),
   303 => (x"02",x"9b",x"73",x"4b"),
   304 => (x"c8",x"87",x"ca",x"c3"),
   305 => (x"78",x"c0",x"48",x"a6"),
   306 => (x"c0",x"d0",x"80",x"fc"),
   307 => (x"78",x"c0",x"c0",x"c0"),
   308 => (x"83",x"c3",x"4d",x"c0"),
   309 => (x"c0",x"d0",x"9b",x"fc"),
   310 => (x"4c",x"c0",x"c0",x"c0"),
   311 => (x"1e",x"74",x"84",x"73"),
   312 => (x"dc",x"1e",x"ee",x"d7"),
   313 => (x"86",x"c8",x"87",x"d2"),
   314 => (x"c1",x"02",x"98",x"70"),
   315 => (x"ff",x"c7",x"87",x"ff"),
   316 => (x"c1",x"06",x"ab",x"b7"),
   317 => (x"c0",x"c8",x"87",x"f7"),
   318 => (x"49",x"66",x"c8",x"1e"),
   319 => (x"1e",x"71",x"81",x"75"),
   320 => (x"87",x"f0",x"c0",x"c1"),
   321 => (x"49",x"70",x"86",x"c8"),
   322 => (x"76",x"59",x"a6",x"d0"),
   323 => (x"c8",x"78",x"24",x"48"),
   324 => (x"cc",x"8b",x"85",x"c0"),
   325 => (x"a8",x"6e",x"48",x"66"),
   326 => (x"87",x"c9",x"c1",x"02"),
   327 => (x"c1",x"48",x"66",x"c8"),
   328 => (x"58",x"a6",x"cc",x"80"),
   329 => (x"1e",x"e8",x"d6",x"c1"),
   330 => (x"d2",x"fc",x"1e",x"75"),
   331 => (x"c1",x"86",x"c8",x"87"),
   332 => (x"c0",x"48",x"f0",x"d6"),
   333 => (x"80",x"c1",x"50",x"e0"),
   334 => (x"66",x"d0",x"1e",x"70"),
   335 => (x"87",x"ff",x"fb",x"1e"),
   336 => (x"d6",x"c1",x"86",x"c8"),
   337 => (x"e0",x"c0",x"48",x"f9"),
   338 => (x"70",x"80",x"c1",x"50"),
   339 => (x"1e",x"66",x"c4",x"1e"),
   340 => (x"c8",x"87",x"ec",x"fb"),
   341 => (x"c2",x"d7",x"c1",x"86"),
   342 => (x"e6",x"50",x"c0",x"48"),
   343 => (x"c0",x"1e",x"70",x"80"),
   344 => (x"c4",x"87",x"ea",x"e4"),
   345 => (x"b7",x"ff",x"c7",x"86"),
   346 => (x"c9",x"fe",x"01",x"ab"),
   347 => (x"05",x"66",x"c8",x"87"),
   348 => (x"d0",x"87",x"da",x"c0"),
   349 => (x"c0",x"c0",x"c0",x"c0"),
   350 => (x"fe",x"4b",x"bf",x"97"),
   351 => (x"73",x"bb",x"83",x"c0"),
   352 => (x"87",x"c9",x"c0",x"0f"),
   353 => (x"c0",x"1e",x"c6",x"d8"),
   354 => (x"c4",x"87",x"c0",x"fe"),
   355 => (x"1e",x"cf",x"d9",x"86"),
   356 => (x"87",x"f7",x"fd",x"c0"),
   357 => (x"d7",x"c1",x"86",x"c4"),
   358 => (x"78",x"c0",x"48",x"e4"),
   359 => (x"ff",x"c8",x"f4",x"c3"),
   360 => (x"e8",x"f6",x"c0",x"4d"),
   361 => (x"c0",x"4c",x"c0",x"c0"),
   362 => (x"fc",x"c0",x"1e",x"ee"),
   363 => (x"86",x"c4",x"87",x"f4"),
   364 => (x"f4",x"c3",x"4a",x"75"),
   365 => (x"6c",x"4d",x"c0",x"c9"),
   366 => (x"c8",x"49",x"73",x"4b"),
   367 => (x"99",x"71",x"99",x"c0"),
   368 => (x"87",x"ce",x"c0",x"02"),
   369 => (x"ff",x"c3",x"49",x"73"),
   370 => (x"f1",x"1e",x"71",x"99"),
   371 => (x"86",x"c4",x"87",x"d3"),
   372 => (x"49",x"72",x"4a",x"75"),
   373 => (x"99",x"71",x"8a",x"c1"),
   374 => (x"87",x"db",x"ff",x"05"),
   375 => (x"ff",x"c8",x"f4",x"c3"),
   376 => (x"87",x"c3",x"ff",x"4d"),
   377 => (x"4d",x"26",x"8e",x"f0"),
   378 => (x"4b",x"26",x"4c",x"26"),
   379 => (x"48",x"43",x"4f",x"26"),
   380 => (x"53",x"4b",x"43",x"45"),
   381 => (x"49",x"42",x"4d",x"55"),
   382 => (x"53",x"4f",x"00",x"4e"),
   383 => (x"32",x"33",x"38",x"44"),
   384 => (x"59",x"53",x"31",x"30"),
   385 => (x"6e",x"55",x"00",x"53"),
   386 => (x"65",x"6c",x"62",x"61"),
   387 => (x"20",x"6f",x"74",x"20"),
   388 => (x"61",x"63",x"6f",x"6c"),
   389 => (x"70",x"20",x"65",x"74"),
   390 => (x"69",x"74",x"72",x"61"),
   391 => (x"6e",x"6f",x"69",x"74"),
   392 => (x"75",x"48",x"00",x"0a"),
   393 => (x"6e",x"69",x"74",x"6e"),
   394 => (x"6f",x"66",x"20",x"67"),
   395 => (x"61",x"70",x"20",x"72"),
   396 => (x"74",x"69",x"74",x"72"),
   397 => (x"0a",x"6e",x"6f",x"69"),
   398 => (x"69",x"6e",x"49",x"00"),
   399 => (x"6c",x"61",x"69",x"74"),
   400 => (x"6e",x"69",x"7a",x"69"),
   401 => (x"44",x"53",x"20",x"67"),
   402 => (x"72",x"61",x"63",x"20"),
   403 => (x"42",x"00",x"0a",x"64"),
   404 => (x"69",x"74",x"6f",x"6f"),
   405 => (x"66",x"20",x"67",x"6e"),
   406 => (x"20",x"6d",x"6f",x"72"),
   407 => (x"33",x"32",x"53",x"52"),
   408 => (x"43",x"00",x"2e",x"32"),
   409 => (x"6b",x"63",x"65",x"68"),
   410 => (x"20",x"6d",x"75",x"73"),
   411 => (x"25",x"20",x"6f",x"74"),
   412 => (x"25",x"20",x"3a",x"64"),
   413 => (x"0e",x"00",x"0a",x"64"),
   414 => (x"5d",x"5c",x"5b",x"5e"),
   415 => (x"4d",x"66",x"d4",x"0e"),
   416 => (x"c0",x"4c",x"66",x"d0"),
   417 => (x"48",x"66",x"d8",x"4b"),
   418 => (x"06",x"a8",x"b7",x"c0"),
   419 => (x"4a",x"14",x"87",x"df"),
   420 => (x"ba",x"82",x"c0",x"fe"),
   421 => (x"c0",x"fe",x"49",x"15"),
   422 => (x"b7",x"71",x"b9",x"81"),
   423 => (x"87",x"c4",x"02",x"aa"),
   424 => (x"87",x"cb",x"48",x"c1"),
   425 => (x"66",x"d8",x"83",x"c1"),
   426 => (x"e1",x"04",x"ab",x"b7"),
   427 => (x"26",x"48",x"c0",x"87"),
   428 => (x"26",x"4c",x"26",x"4d"),
   429 => (x"0e",x"4f",x"26",x"4b"),
   430 => (x"5d",x"5c",x"5b",x"5e"),
   431 => (x"f0",x"df",x"c1",x"0e"),
   432 => (x"c0",x"78",x"c0",x"48"),
   433 => (x"c0",x"1e",x"f8",x"f5"),
   434 => (x"c4",x"87",x"c0",x"f9"),
   435 => (x"e8",x"d7",x"c1",x"86"),
   436 => (x"c0",x"1e",x"c0",x"1e"),
   437 => (x"c8",x"87",x"d6",x"f4"),
   438 => (x"05",x"98",x"70",x"86"),
   439 => (x"f2",x"c0",x"87",x"cf"),
   440 => (x"f8",x"c0",x"1e",x"e4"),
   441 => (x"86",x"c4",x"87",x"e5"),
   442 => (x"d2",x"cb",x"48",x"c0"),
   443 => (x"c5",x"f6",x"c0",x"87"),
   444 => (x"d6",x"f8",x"c0",x"1e"),
   445 => (x"c0",x"86",x"c4",x"87"),
   446 => (x"dc",x"e0",x"c1",x"4b"),
   447 => (x"c8",x"78",x"c1",x"48"),
   448 => (x"dc",x"f6",x"c0",x"1e"),
   449 => (x"de",x"d8",x"c1",x"1e"),
   450 => (x"87",x"eb",x"fd",x"1e"),
   451 => (x"98",x"70",x"86",x"cc"),
   452 => (x"c1",x"87",x"c6",x"05"),
   453 => (x"c0",x"48",x"dc",x"e0"),
   454 => (x"c0",x"1e",x"c8",x"78"),
   455 => (x"c1",x"1e",x"e5",x"f6"),
   456 => (x"fd",x"1e",x"fa",x"d8"),
   457 => (x"86",x"cc",x"87",x"d1"),
   458 => (x"c6",x"05",x"98",x"70"),
   459 => (x"dc",x"e0",x"c1",x"87"),
   460 => (x"c1",x"78",x"c0",x"48"),
   461 => (x"1e",x"bf",x"dc",x"e0"),
   462 => (x"1e",x"ee",x"f6",x"c0"),
   463 => (x"c8",x"87",x"fd",x"e3"),
   464 => (x"dc",x"e0",x"c1",x"86"),
   465 => (x"d7",x"c2",x"02",x"bf"),
   466 => (x"e8",x"d7",x"c1",x"87"),
   467 => (x"e6",x"de",x"c1",x"4d"),
   468 => (x"e6",x"df",x"c1",x"4c"),
   469 => (x"71",x"49",x"bf",x"9f"),
   470 => (x"e6",x"df",x"c1",x"1e"),
   471 => (x"e8",x"d7",x"c1",x"49"),
   472 => (x"d0",x"1e",x"71",x"89"),
   473 => (x"1e",x"c0",x"c8",x"1e"),
   474 => (x"1e",x"d6",x"f3",x"c0"),
   475 => (x"d4",x"87",x"cd",x"e3"),
   476 => (x"c8",x"49",x"74",x"86"),
   477 => (x"c1",x"4b",x"69",x"81"),
   478 => (x"bf",x"9f",x"e6",x"df"),
   479 => (x"ea",x"d6",x"c5",x"49"),
   480 => (x"d0",x"c0",x"05",x"a9"),
   481 => (x"c8",x"49",x"74",x"87"),
   482 => (x"e7",x"1e",x"69",x"81"),
   483 => (x"86",x"c4",x"87",x"f7"),
   484 => (x"df",x"c0",x"4b",x"70"),
   485 => (x"c7",x"49",x"75",x"87"),
   486 => (x"69",x"9f",x"81",x"fe"),
   487 => (x"d5",x"e9",x"ca",x"49"),
   488 => (x"cf",x"c0",x"02",x"a9"),
   489 => (x"f8",x"f2",x"c0",x"87"),
   490 => (x"de",x"f5",x"c0",x"1e"),
   491 => (x"c0",x"86",x"c4",x"87"),
   492 => (x"87",x"cb",x"c8",x"48"),
   493 => (x"f4",x"c0",x"1e",x"73"),
   494 => (x"ff",x"e1",x"1e",x"d3"),
   495 => (x"c1",x"86",x"c8",x"87"),
   496 => (x"73",x"1e",x"e8",x"d7"),
   497 => (x"e4",x"f0",x"c0",x"1e"),
   498 => (x"70",x"86",x"c8",x"87"),
   499 => (x"c5",x"c0",x"05",x"98"),
   500 => (x"c7",x"48",x"c0",x"87"),
   501 => (x"f4",x"c0",x"87",x"e9"),
   502 => (x"f4",x"c0",x"1e",x"eb"),
   503 => (x"86",x"c4",x"87",x"ed"),
   504 => (x"1e",x"c1",x"f7",x"c0"),
   505 => (x"c4",x"87",x"d5",x"e1"),
   506 => (x"c0",x"1e",x"c8",x"86"),
   507 => (x"c1",x"1e",x"d9",x"f7"),
   508 => (x"fa",x"1e",x"fa",x"d8"),
   509 => (x"86",x"cc",x"87",x"c1"),
   510 => (x"c0",x"05",x"98",x"70"),
   511 => (x"df",x"c1",x"87",x"c9"),
   512 => (x"78",x"c1",x"48",x"f0"),
   513 => (x"c8",x"87",x"e3",x"c0"),
   514 => (x"e2",x"f7",x"c0",x"1e"),
   515 => (x"de",x"d8",x"c1",x"1e"),
   516 => (x"87",x"e3",x"f9",x"1e"),
   517 => (x"98",x"70",x"86",x"cc"),
   518 => (x"87",x"ce",x"c0",x"02"),
   519 => (x"1e",x"d2",x"f5",x"c0"),
   520 => (x"c4",x"87",x"d9",x"e0"),
   521 => (x"c6",x"48",x"c0",x"86"),
   522 => (x"df",x"c1",x"87",x"d5"),
   523 => (x"49",x"bf",x"97",x"e6"),
   524 => (x"05",x"a9",x"d5",x"c1"),
   525 => (x"c1",x"87",x"cd",x"c0"),
   526 => (x"bf",x"97",x"e7",x"df"),
   527 => (x"a9",x"ea",x"c2",x"49"),
   528 => (x"87",x"c5",x"c0",x"02"),
   529 => (x"f6",x"c5",x"48",x"c0"),
   530 => (x"e8",x"d7",x"c1",x"87"),
   531 => (x"c3",x"49",x"bf",x"97"),
   532 => (x"c0",x"02",x"a9",x"e9"),
   533 => (x"d7",x"c1",x"87",x"d2"),
   534 => (x"49",x"bf",x"97",x"e8"),
   535 => (x"02",x"a9",x"eb",x"c3"),
   536 => (x"c0",x"87",x"c5",x"c0"),
   537 => (x"87",x"d7",x"c5",x"48"),
   538 => (x"97",x"f3",x"d7",x"c1"),
   539 => (x"99",x"71",x"49",x"bf"),
   540 => (x"87",x"cc",x"c0",x"05"),
   541 => (x"97",x"f4",x"d7",x"c1"),
   542 => (x"a9",x"c2",x"49",x"bf"),
   543 => (x"87",x"c5",x"c0",x"02"),
   544 => (x"fa",x"c4",x"48",x"c0"),
   545 => (x"f5",x"d7",x"c1",x"87"),
   546 => (x"c1",x"48",x"bf",x"97"),
   547 => (x"c1",x"58",x"ec",x"df"),
   548 => (x"49",x"bf",x"e8",x"df"),
   549 => (x"8a",x"c1",x"4a",x"71"),
   550 => (x"5a",x"f0",x"df",x"c1"),
   551 => (x"1e",x"71",x"1e",x"72"),
   552 => (x"1e",x"eb",x"f7",x"c0"),
   553 => (x"87",x"d4",x"de",x"ff"),
   554 => (x"d7",x"c1",x"86",x"cc"),
   555 => (x"49",x"bf",x"97",x"f6"),
   556 => (x"d7",x"c1",x"81",x"73"),
   557 => (x"4a",x"bf",x"97",x"f7"),
   558 => (x"48",x"72",x"32",x"c8"),
   559 => (x"e0",x"c1",x"80",x"71"),
   560 => (x"d7",x"c1",x"58",x"c0"),
   561 => (x"48",x"bf",x"97",x"f8"),
   562 => (x"58",x"d4",x"e0",x"c1"),
   563 => (x"bf",x"f0",x"df",x"c1"),
   564 => (x"87",x"da",x"c2",x"02"),
   565 => (x"f5",x"c0",x"1e",x"c8"),
   566 => (x"d8",x"c1",x"1e",x"ef"),
   567 => (x"d6",x"f6",x"1e",x"fa"),
   568 => (x"70",x"86",x"cc",x"87"),
   569 => (x"c5",x"c0",x"02",x"98"),
   570 => (x"c3",x"48",x"c0",x"87"),
   571 => (x"df",x"c1",x"87",x"d1"),
   572 => (x"72",x"4a",x"bf",x"e8"),
   573 => (x"c1",x"30",x"c4",x"48"),
   574 => (x"c1",x"58",x"d8",x"e0"),
   575 => (x"c1",x"5a",x"d0",x"e0"),
   576 => (x"bf",x"97",x"cd",x"d8"),
   577 => (x"c1",x"31",x"c8",x"49"),
   578 => (x"bf",x"97",x"cc",x"d8"),
   579 => (x"c1",x"81",x"73",x"4b"),
   580 => (x"bf",x"97",x"ce",x"d8"),
   581 => (x"73",x"33",x"d0",x"4b"),
   582 => (x"cf",x"d8",x"c1",x"81"),
   583 => (x"d8",x"4b",x"bf",x"97"),
   584 => (x"c1",x"81",x"73",x"33"),
   585 => (x"c1",x"59",x"dc",x"e0"),
   586 => (x"91",x"bf",x"d0",x"e0"),
   587 => (x"bf",x"fc",x"df",x"c1"),
   588 => (x"c4",x"e0",x"c1",x"81"),
   589 => (x"d5",x"d8",x"c1",x"59"),
   590 => (x"c8",x"4b",x"bf",x"97"),
   591 => (x"d4",x"d8",x"c1",x"33"),
   592 => (x"74",x"4c",x"bf",x"97"),
   593 => (x"d6",x"d8",x"c1",x"83"),
   594 => (x"d0",x"4c",x"bf",x"97"),
   595 => (x"c1",x"83",x"74",x"34"),
   596 => (x"bf",x"97",x"d7",x"d8"),
   597 => (x"d8",x"9c",x"cf",x"4c"),
   598 => (x"c1",x"83",x"74",x"34"),
   599 => (x"c2",x"5b",x"c8",x"e0"),
   600 => (x"72",x"92",x"73",x"8b"),
   601 => (x"c1",x"80",x"71",x"48"),
   602 => (x"c1",x"58",x"cc",x"e0"),
   603 => (x"d7",x"c1",x"87",x"cf"),
   604 => (x"49",x"bf",x"97",x"fa"),
   605 => (x"d7",x"c1",x"31",x"c8"),
   606 => (x"4a",x"bf",x"97",x"f9"),
   607 => (x"e0",x"c1",x"81",x"72"),
   608 => (x"31",x"c5",x"59",x"d8"),
   609 => (x"c9",x"81",x"ff",x"c7"),
   610 => (x"d0",x"e0",x"c1",x"29"),
   611 => (x"ff",x"d7",x"c1",x"59"),
   612 => (x"c8",x"4a",x"bf",x"97"),
   613 => (x"fe",x"d7",x"c1",x"32"),
   614 => (x"73",x"4b",x"bf",x"97"),
   615 => (x"dc",x"e0",x"c1",x"82"),
   616 => (x"d0",x"e0",x"c1",x"5a"),
   617 => (x"df",x"c1",x"92",x"bf"),
   618 => (x"c1",x"82",x"bf",x"fc"),
   619 => (x"c1",x"5a",x"cc",x"e0"),
   620 => (x"c0",x"48",x"c4",x"e0"),
   621 => (x"71",x"48",x"72",x"78"),
   622 => (x"c4",x"e0",x"c1",x"80"),
   623 => (x"26",x"48",x"c1",x"58"),
   624 => (x"26",x"4c",x"26",x"4d"),
   625 => (x"0e",x"4f",x"26",x"4b"),
   626 => (x"0e",x"5c",x"5b",x"5e"),
   627 => (x"bf",x"f0",x"df",x"c1"),
   628 => (x"87",x"cf",x"c0",x"02"),
   629 => (x"c7",x"4a",x"66",x"cc"),
   630 => (x"66",x"cc",x"2a",x"b7"),
   631 => (x"9b",x"ff",x"c1",x"4b"),
   632 => (x"cc",x"87",x"cc",x"c0"),
   633 => (x"b7",x"c8",x"4a",x"66"),
   634 => (x"4b",x"66",x"cc",x"2a"),
   635 => (x"c1",x"9b",x"ff",x"c3"),
   636 => (x"c1",x"1e",x"e8",x"d7"),
   637 => (x"49",x"bf",x"fc",x"df"),
   638 => (x"1e",x"71",x"81",x"72"),
   639 => (x"87",x"ed",x"e7",x"c0"),
   640 => (x"98",x"70",x"86",x"c8"),
   641 => (x"87",x"c5",x"c0",x"05"),
   642 => (x"ea",x"c0",x"48",x"c0"),
   643 => (x"f0",x"df",x"c1",x"87"),
   644 => (x"d4",x"c0",x"02",x"bf"),
   645 => (x"c4",x"49",x"73",x"87"),
   646 => (x"d7",x"c1",x"91",x"b7"),
   647 => (x"4c",x"69",x"81",x"e8"),
   648 => (x"ff",x"ff",x"ff",x"cf"),
   649 => (x"cc",x"c0",x"9c",x"ff"),
   650 => (x"c2",x"49",x"73",x"87"),
   651 => (x"d7",x"c1",x"91",x"b7"),
   652 => (x"69",x"9f",x"81",x"e8"),
   653 => (x"26",x"48",x"74",x"4c"),
   654 => (x"26",x"4b",x"26",x"4c"),
   655 => (x"5b",x"5e",x"0e",x"4f"),
   656 => (x"f0",x"0e",x"5d",x"5c"),
   657 => (x"ff",x"ff",x"cf",x"86"),
   658 => (x"c0",x"4c",x"f8",x"ff"),
   659 => (x"c1",x"48",x"76",x"4b"),
   660 => (x"78",x"bf",x"c4",x"e0"),
   661 => (x"e0",x"c1",x"80",x"c4"),
   662 => (x"c1",x"78",x"bf",x"c8"),
   663 => (x"02",x"bf",x"f0",x"df"),
   664 => (x"c1",x"87",x"ca",x"c0"),
   665 => (x"49",x"bf",x"e8",x"df"),
   666 => (x"c7",x"c0",x"31",x"c4"),
   667 => (x"cc",x"e0",x"c1",x"87"),
   668 => (x"31",x"c4",x"49",x"bf"),
   669 => (x"cc",x"59",x"a6",x"cc"),
   670 => (x"78",x"c0",x"48",x"a6"),
   671 => (x"c0",x"48",x"66",x"c8"),
   672 => (x"fc",x"c2",x"06",x"a8"),
   673 => (x"4d",x"66",x"cc",x"87"),
   674 => (x"99",x"cf",x"49",x"75"),
   675 => (x"c0",x"05",x"99",x"71"),
   676 => (x"d7",x"c1",x"87",x"dc"),
   677 => (x"66",x"c8",x"1e",x"e8"),
   678 => (x"80",x"c1",x"48",x"49"),
   679 => (x"71",x"58",x"a6",x"cc"),
   680 => (x"c8",x"e5",x"c0",x"1e"),
   681 => (x"c1",x"86",x"c8",x"87"),
   682 => (x"c0",x"4b",x"e8",x"d7"),
   683 => (x"e0",x"c0",x"87",x"c3"),
   684 => (x"49",x"6b",x"97",x"83"),
   685 => (x"c1",x"02",x"99",x"71"),
   686 => (x"6b",x"97",x"87",x"fe"),
   687 => (x"a9",x"e5",x"c3",x"49"),
   688 => (x"87",x"f4",x"c1",x"02"),
   689 => (x"81",x"cb",x"49",x"73"),
   690 => (x"d8",x"49",x"69",x"97"),
   691 => (x"05",x"99",x"71",x"99"),
   692 => (x"73",x"87",x"e5",x"c1"),
   693 => (x"f2",x"e8",x"c0",x"1e"),
   694 => (x"cb",x"86",x"c4",x"87"),
   695 => (x"66",x"e8",x"c0",x"1e"),
   696 => (x"ee",x"1e",x"73",x"1e"),
   697 => (x"86",x"cc",x"87",x"d1"),
   698 => (x"c1",x"05",x"98",x"70"),
   699 => (x"4a",x"73",x"87",x"ca"),
   700 => (x"e0",x"c0",x"82",x"dc"),
   701 => (x"81",x"c4",x"49",x"66"),
   702 => (x"4a",x"73",x"79",x"6a"),
   703 => (x"e0",x"c0",x"82",x"da"),
   704 => (x"81",x"c8",x"49",x"66"),
   705 => (x"70",x"48",x"6a",x"9f"),
   706 => (x"c1",x"4c",x"71",x"79"),
   707 => (x"02",x"bf",x"f0",x"df"),
   708 => (x"73",x"87",x"d2",x"c0"),
   709 => (x"9f",x"81",x"d4",x"49"),
   710 => (x"ff",x"c0",x"49",x"69"),
   711 => (x"4a",x"71",x"99",x"ff"),
   712 => (x"c2",x"c0",x"32",x"d0"),
   713 => (x"72",x"4a",x"c0",x"87"),
   714 => (x"70",x"80",x"6c",x"48"),
   715 => (x"66",x"e0",x"c0",x"7c"),
   716 => (x"c1",x"78",x"c0",x"48"),
   717 => (x"87",x"c3",x"c1",x"48"),
   718 => (x"66",x"c8",x"85",x"c1"),
   719 => (x"c7",x"fd",x"04",x"ad"),
   720 => (x"ff",x"ff",x"cf",x"87"),
   721 => (x"c1",x"4c",x"f8",x"ff"),
   722 => (x"02",x"bf",x"f0",x"df"),
   723 => (x"6e",x"87",x"ea",x"c0"),
   724 => (x"87",x"f3",x"f9",x"1e"),
   725 => (x"a6",x"c4",x"86",x"c4"),
   726 => (x"74",x"49",x"6e",x"58"),
   727 => (x"02",x"a9",x"74",x"99"),
   728 => (x"6e",x"87",x"d6",x"c0"),
   729 => (x"c1",x"89",x"c2",x"49"),
   730 => (x"91",x"bf",x"e8",x"df"),
   731 => (x"bf",x"c0",x"e0",x"c1"),
   732 => (x"c8",x"80",x"71",x"48"),
   733 => (x"fe",x"fb",x"58",x"a6"),
   734 => (x"cf",x"48",x"c0",x"87"),
   735 => (x"f8",x"ff",x"ff",x"ff"),
   736 => (x"26",x"8e",x"f0",x"4c"),
   737 => (x"26",x"4c",x"26",x"4d"),
   738 => (x"0e",x"4f",x"26",x"4b"),
   739 => (x"c8",x"0e",x"5b",x"5e"),
   740 => (x"c1",x"49",x"bf",x"66"),
   741 => (x"09",x"66",x"c8",x"81"),
   742 => (x"df",x"c1",x"09",x"79"),
   743 => (x"71",x"99",x"bf",x"ec"),
   744 => (x"d0",x"c0",x"05",x"99"),
   745 => (x"4b",x"66",x"c8",x"87"),
   746 => (x"1e",x"6b",x"83",x"c8"),
   747 => (x"c4",x"87",x"d8",x"f8"),
   748 => (x"71",x"49",x"70",x"86"),
   749 => (x"26",x"48",x"c1",x"7b"),
   750 => (x"0e",x"4f",x"26",x"4b"),
   751 => (x"e0",x"c1",x"0e",x"5e"),
   752 => (x"c4",x"49",x"bf",x"c0"),
   753 => (x"82",x"c8",x"4a",x"66"),
   754 => (x"8a",x"c2",x"4a",x"6a"),
   755 => (x"bf",x"e8",x"df",x"c1"),
   756 => (x"c1",x"81",x"72",x"92"),
   757 => (x"4a",x"bf",x"ec",x"df"),
   758 => (x"9a",x"bf",x"66",x"c4"),
   759 => (x"66",x"c8",x"81",x"72"),
   760 => (x"c0",x"1e",x"71",x"1e"),
   761 => (x"c8",x"87",x"c6",x"e0"),
   762 => (x"05",x"98",x"70",x"86"),
   763 => (x"c0",x"87",x"c5",x"c0"),
   764 => (x"87",x"c2",x"c0",x"48"),
   765 => (x"4f",x"26",x"48",x"c1"),
   766 => (x"5c",x"5b",x"5e",x"0e"),
   767 => (x"66",x"d4",x"0e",x"5d"),
   768 => (x"1e",x"66",x"d0",x"4c"),
   769 => (x"1e",x"e0",x"e0",x"c1"),
   770 => (x"c8",x"87",x"f2",x"f8"),
   771 => (x"02",x"98",x"70",x"86"),
   772 => (x"c1",x"87",x"cd",x"c1"),
   773 => (x"49",x"bf",x"e4",x"e0"),
   774 => (x"c9",x"81",x"ff",x"c7"),
   775 => (x"c0",x"4d",x"71",x"29"),
   776 => (x"fc",x"f1",x"c0",x"4b"),
   777 => (x"e2",x"e3",x"c0",x"1e"),
   778 => (x"c0",x"86",x"c4",x"87"),
   779 => (x"c1",x"06",x"ad",x"b7"),
   780 => (x"1e",x"74",x"87",x"c0"),
   781 => (x"1e",x"e0",x"e0",x"c1"),
   782 => (x"c8",x"87",x"c0",x"fe"),
   783 => (x"05",x"98",x"70",x"86"),
   784 => (x"c0",x"87",x"c5",x"c0"),
   785 => (x"87",x"ec",x"c0",x"48"),
   786 => (x"1e",x"e0",x"e0",x"c1"),
   787 => (x"c4",x"87",x"fc",x"fc"),
   788 => (x"84",x"c0",x"c8",x"86"),
   789 => (x"b7",x"75",x"83",x"c1"),
   790 => (x"d5",x"ff",x"04",x"ab"),
   791 => (x"87",x"d2",x"c0",x"87"),
   792 => (x"c0",x"1e",x"66",x"d0"),
   793 => (x"ff",x"1e",x"d5",x"f2"),
   794 => (x"c8",x"87",x"d1",x"cf"),
   795 => (x"c0",x"48",x"c0",x"86"),
   796 => (x"48",x"c1",x"87",x"c2"),
   797 => (x"4c",x"26",x"4d",x"26"),
   798 => (x"4f",x"26",x"4b",x"26"),
   799 => (x"6e",x"65",x"70",x"4f"),
   800 => (x"66",x"20",x"64",x"65"),
   801 => (x"2c",x"65",x"6c",x"69"),
   802 => (x"61",x"6f",x"6c",x"20"),
   803 => (x"67",x"6e",x"69",x"64"),
   804 => (x"0a",x"2e",x"2e",x"2e"),
   805 => (x"6e",x"61",x"43",x"00"),
   806 => (x"6f",x"20",x"74",x"27"),
   807 => (x"20",x"6e",x"65",x"70"),
   808 => (x"00",x"0a",x"73",x"25"),
   809 => (x"64",x"61",x"65",x"52"),
   810 => (x"20",x"66",x"6f",x"20"),
   811 => (x"20",x"52",x"42",x"4d"),
   812 => (x"6c",x"69",x"61",x"66"),
   813 => (x"00",x"0a",x"64",x"65"),
   814 => (x"70",x"20",x"6f",x"4e"),
   815 => (x"69",x"74",x"72",x"61"),
   816 => (x"6e",x"6f",x"69",x"74"),
   817 => (x"67",x"69",x"73",x"20"),
   818 => (x"75",x"74",x"61",x"6e"),
   819 => (x"66",x"20",x"65",x"72"),
   820 => (x"64",x"6e",x"75",x"6f"),
   821 => (x"42",x"4d",x"00",x"0a"),
   822 => (x"7a",x"69",x"73",x"52"),
   823 => (x"25",x"20",x"3a",x"65"),
   824 => (x"70",x"20",x"2c",x"64"),
   825 => (x"69",x"74",x"72",x"61"),
   826 => (x"6e",x"6f",x"69",x"74"),
   827 => (x"65",x"7a",x"69",x"73"),
   828 => (x"64",x"25",x"20",x"3a"),
   829 => (x"66",x"6f",x"20",x"2c"),
   830 => (x"74",x"65",x"73",x"66"),
   831 => (x"20",x"66",x"6f",x"20"),
   832 => (x"3a",x"67",x"69",x"73"),
   833 => (x"2c",x"64",x"25",x"20"),
   834 => (x"67",x"69",x"73",x"20"),
   835 => (x"25",x"78",x"30",x"20"),
   836 => (x"52",x"00",x"0a",x"78"),
   837 => (x"69",x"64",x"61",x"65"),
   838 => (x"62",x"20",x"67",x"6e"),
   839 => (x"20",x"74",x"6f",x"6f"),
   840 => (x"74",x"63",x"65",x"73"),
   841 => (x"25",x"20",x"72",x"6f"),
   842 => (x"52",x"00",x"0a",x"64"),
   843 => (x"20",x"64",x"61",x"65"),
   844 => (x"74",x"6f",x"6f",x"62"),
   845 => (x"63",x"65",x"73",x"20"),
   846 => (x"20",x"72",x"6f",x"74"),
   847 => (x"6d",x"6f",x"72",x"66"),
   848 => (x"72",x"69",x"66",x"20"),
   849 => (x"70",x"20",x"74",x"73"),
   850 => (x"69",x"74",x"72",x"61"),
   851 => (x"6e",x"6f",x"69",x"74"),
   852 => (x"6e",x"55",x"00",x"0a"),
   853 => (x"70",x"70",x"75",x"73"),
   854 => (x"65",x"74",x"72",x"6f"),
   855 => (x"61",x"70",x"20",x"64"),
   856 => (x"74",x"69",x"74",x"72"),
   857 => (x"20",x"6e",x"6f",x"69"),
   858 => (x"65",x"70",x"79",x"74"),
   859 => (x"46",x"00",x"0d",x"21"),
   860 => (x"32",x"33",x"54",x"41"),
   861 => (x"00",x"20",x"20",x"20"),
   862 => (x"64",x"61",x"65",x"52"),
   863 => (x"20",x"67",x"6e",x"69"),
   864 => (x"0a",x"52",x"42",x"4d"),
   865 => (x"52",x"42",x"4d",x"00"),
   866 => (x"63",x"75",x"73",x"20"),
   867 => (x"73",x"73",x"65",x"63"),
   868 => (x"6c",x"6c",x"75",x"66"),
   869 => (x"65",x"72",x"20",x"79"),
   870 => (x"00",x"0a",x"64",x"61"),
   871 => (x"31",x"54",x"41",x"46"),
   872 => (x"20",x"20",x"20",x"36"),
   873 => (x"54",x"41",x"46",x"00"),
   874 => (x"20",x"20",x"32",x"33"),
   875 => (x"61",x"50",x"00",x"20"),
   876 => (x"74",x"69",x"74",x"72"),
   877 => (x"63",x"6e",x"6f",x"69"),
   878 => (x"74",x"6e",x"75",x"6f"),
   879 => (x"0a",x"64",x"25",x"20"),
   880 => (x"6e",x"75",x"48",x"00"),
   881 => (x"67",x"6e",x"69",x"74"),
   882 => (x"72",x"6f",x"66",x"20"),
   883 => (x"6c",x"69",x"66",x"20"),
   884 => (x"73",x"79",x"73",x"65"),
   885 => (x"0a",x"6d",x"65",x"74"),
   886 => (x"54",x"41",x"46",x"00"),
   887 => (x"20",x"20",x"32",x"33"),
   888 => (x"41",x"46",x"00",x"20"),
   889 => (x"20",x"36",x"31",x"54"),
   890 => (x"43",x"00",x"20",x"20"),
   891 => (x"74",x"73",x"75",x"6c"),
   892 => (x"73",x"20",x"72",x"65"),
   893 => (x"3a",x"65",x"7a",x"69"),
   894 => (x"2c",x"64",x"25",x"20"),
   895 => (x"75",x"6c",x"43",x"20"),
   896 => (x"72",x"65",x"74",x"73"),
   897 => (x"73",x"61",x"6d",x"20"),
   898 => (x"25",x"20",x"2c",x"6b"),
   899 => (x"1e",x"00",x"0a",x"64"),
   900 => (x"cd",x"02",x"66",x"c4"),
   901 => (x"ec",x"e0",x"c1",x"87"),
   902 => (x"78",x"66",x"c4",x"48"),
   903 => (x"48",x"f4",x"e0",x"c1"),
   904 => (x"e0",x"c1",x"78",x"c0"),
   905 => (x"d5",x"05",x"bf",x"f4"),
   906 => (x"ec",x"e0",x"c1",x"87"),
   907 => (x"48",x"71",x"49",x"bf"),
   908 => (x"e0",x"c1",x"80",x"c4"),
   909 => (x"e0",x"c1",x"58",x"f0"),
   910 => (x"78",x"69",x"48",x"f0"),
   911 => (x"e0",x"c1",x"87",x"cb"),
   912 => (x"c8",x"48",x"bf",x"f0"),
   913 => (x"f4",x"e0",x"c1",x"30"),
   914 => (x"f4",x"e0",x"c1",x"58"),
   915 => (x"81",x"c1",x"49",x"bf"),
   916 => (x"98",x"c3",x"48",x"71"),
   917 => (x"58",x"f8",x"e0",x"c1"),
   918 => (x"bf",x"f0",x"e0",x"c1"),
   919 => (x"29",x"b7",x"d8",x"49"),
   920 => (x"4f",x"26",x"48",x"71"),
   921 => (x"0e",x"5b",x"5e",x"0e"),
   922 => (x"fe",x"1e",x"66",x"c8"),
   923 => (x"86",x"c4",x"87",x"e1"),
   924 => (x"4b",x"c0",x"49",x"70"),
   925 => (x"ce",x"02",x"99",x"71"),
   926 => (x"c0",x"83",x"c1",x"87"),
   927 => (x"87",x"cf",x"fe",x"1e"),
   928 => (x"49",x"70",x"86",x"c4"),
   929 => (x"73",x"87",x"ed",x"ff"),
   930 => (x"26",x"4b",x"26",x"48"),
   931 => (x"5b",x"5e",x"0e",x"4f"),
   932 => (x"f8",x"0e",x"5d",x"5c"),
   933 => (x"e4",x"f6",x"c0",x"86"),
   934 => (x"c0",x"4c",x"c4",x"c0"),
   935 => (x"c0",x"c0",x"e4",x"f6"),
   936 => (x"1e",x"66",x"d8",x"4b"),
   937 => (x"c4",x"87",x"fd",x"fe"),
   938 => (x"71",x"49",x"70",x"86"),
   939 => (x"76",x"85",x"c2",x"4d"),
   940 => (x"d0",x"78",x"c1",x"48"),
   941 => (x"c0",x"c1",x"7c",x"9f"),
   942 => (x"9f",x"7b",x"9f",x"c1"),
   943 => (x"9f",x"c0",x"49",x"6b"),
   944 => (x"9f",x"7b",x"9f",x"7b"),
   945 => (x"a6",x"c8",x"48",x"6b"),
   946 => (x"99",x"c0",x"c4",x"58"),
   947 => (x"c1",x"02",x"99",x"71"),
   948 => (x"02",x"6e",x"87",x"f5"),
   949 => (x"c4",x"87",x"e9",x"c0"),
   950 => (x"c0",x"c8",x"48",x"66"),
   951 => (x"c1",x"05",x"a8",x"c6"),
   952 => (x"48",x"76",x"87",x"e5"),
   953 => (x"eb",x"ca",x"78",x"c0"),
   954 => (x"c1",x"7b",x"9f",x"ca"),
   955 => (x"9f",x"c0",x"7b",x"9f"),
   956 => (x"7b",x"9f",x"75",x"7b"),
   957 => (x"98",x"ff",x"ff",x"cf"),
   958 => (x"9f",x"7b",x"9f",x"c0"),
   959 => (x"87",x"c7",x"c1",x"7b"),
   960 => (x"29",x"c1",x"49",x"75"),
   961 => (x"b1",x"c0",x"c0",x"c8"),
   962 => (x"05",x"a9",x"66",x"c4"),
   963 => (x"d8",x"87",x"f8",x"c0"),
   964 => (x"fa",x"fb",x"1e",x"66"),
   965 => (x"70",x"86",x"c4",x"87"),
   966 => (x"c1",x"49",x"75",x"4a"),
   967 => (x"02",x"99",x"71",x"8d"),
   968 => (x"97",x"72",x"87",x"de"),
   969 => (x"98",x"ff",x"c3",x"7b"),
   970 => (x"c9",x"02",x"9a",x"72"),
   971 => (x"fb",x"1e",x"c0",x"87"),
   972 => (x"86",x"c4",x"87",x"dd"),
   973 => (x"49",x"75",x"4a",x"70"),
   974 => (x"99",x"71",x"8d",x"c1"),
   975 => (x"87",x"e2",x"ff",x"05"),
   976 => (x"c1",x"7c",x"9f",x"d1"),
   977 => (x"d1",x"87",x"c6",x"48"),
   978 => (x"e6",x"fd",x"7c",x"9f"),
   979 => (x"26",x"8e",x"f8",x"87"),
   980 => (x"26",x"4c",x"26",x"4d"),
   981 => (x"0e",x"4f",x"26",x"4b"),
   982 => (x"ff",x"0e",x"5b",x"5e"),
   983 => (x"ff",x"c3",x"86",x"dc"),
   984 => (x"e4",x"f6",x"c0",x"4b"),
   985 => (x"73",x"4a",x"c0",x"c0"),
   986 => (x"73",x"49",x"6a",x"7a"),
   987 => (x"6a",x"7a",x"73",x"99"),
   988 => (x"c4",x"98",x"73",x"48"),
   989 => (x"48",x"6e",x"58",x"a6"),
   990 => (x"a6",x"c8",x"30",x"c8"),
   991 => (x"59",x"a6",x"cc",x"58"),
   992 => (x"73",x"b1",x"66",x"c4"),
   993 => (x"73",x"48",x"6a",x"7a"),
   994 => (x"58",x"a6",x"d0",x"98"),
   995 => (x"d0",x"48",x"66",x"cc"),
   996 => (x"58",x"a6",x"d4",x"30"),
   997 => (x"d0",x"59",x"a6",x"d8"),
   998 => (x"7a",x"73",x"b1",x"66"),
   999 => (x"98",x"73",x"48",x"6a"),
  1000 => (x"d8",x"58",x"a6",x"dc"),
  1001 => (x"30",x"d8",x"48",x"66"),
  1002 => (x"58",x"a6",x"e0",x"c0"),
  1003 => (x"59",x"a6",x"e4",x"c0"),
  1004 => (x"71",x"b1",x"66",x"dc"),
  1005 => (x"8e",x"dc",x"ff",x"48"),
  1006 => (x"4f",x"26",x"4b",x"26"),
  1007 => (x"0e",x"5b",x"5e",x"0e"),
  1008 => (x"ff",x"c3",x"86",x"e8"),
  1009 => (x"e4",x"f6",x"c0",x"4b"),
  1010 => (x"73",x"4a",x"c0",x"c0"),
  1011 => (x"73",x"49",x"6a",x"7a"),
  1012 => (x"c8",x"7a",x"73",x"99"),
  1013 => (x"73",x"48",x"6a",x"31"),
  1014 => (x"58",x"a6",x"c4",x"98"),
  1015 => (x"6e",x"59",x"a6",x"c8"),
  1016 => (x"c8",x"7a",x"73",x"b1"),
  1017 => (x"73",x"48",x"6a",x"31"),
  1018 => (x"58",x"a6",x"cc",x"98"),
  1019 => (x"c8",x"59",x"a6",x"d0"),
  1020 => (x"7a",x"73",x"b1",x"66"),
  1021 => (x"48",x"6a",x"31",x"c8"),
  1022 => (x"a6",x"d4",x"98",x"73"),
  1023 => (x"59",x"a6",x"d8",x"58"),
  1024 => (x"71",x"b1",x"66",x"d0"),
  1025 => (x"26",x"8e",x"e8",x"48"),
  1026 => (x"0e",x"4f",x"26",x"4b"),
  1027 => (x"5d",x"5c",x"5b",x"5e"),
  1028 => (x"4d",x"ff",x"c3",x"0e"),
  1029 => (x"c0",x"e4",x"f6",x"c0"),
  1030 => (x"66",x"d0",x"4b",x"c0"),
  1031 => (x"98",x"ff",x"c3",x"48"),
  1032 => (x"e0",x"c1",x"7b",x"70"),
  1033 => (x"c8",x"05",x"bf",x"f8"),
  1034 => (x"48",x"66",x"d4",x"87"),
  1035 => (x"a6",x"d8",x"30",x"c9"),
  1036 => (x"49",x"66",x"d4",x"58"),
  1037 => (x"48",x"71",x"29",x"d8"),
  1038 => (x"70",x"98",x"ff",x"c3"),
  1039 => (x"49",x"66",x"d4",x"7b"),
  1040 => (x"48",x"71",x"29",x"d0"),
  1041 => (x"70",x"98",x"ff",x"c3"),
  1042 => (x"49",x"66",x"d4",x"7b"),
  1043 => (x"48",x"71",x"29",x"c8"),
  1044 => (x"70",x"98",x"ff",x"c3"),
  1045 => (x"48",x"66",x"d4",x"7b"),
  1046 => (x"70",x"98",x"ff",x"c3"),
  1047 => (x"49",x"66",x"d0",x"7b"),
  1048 => (x"48",x"71",x"29",x"d0"),
  1049 => (x"70",x"98",x"ff",x"c3"),
  1050 => (x"75",x"4c",x"6b",x"7b"),
  1051 => (x"ff",x"f0",x"c9",x"9c"),
  1052 => (x"05",x"ac",x"75",x"4a"),
  1053 => (x"7b",x"75",x"87",x"d2"),
  1054 => (x"9c",x"75",x"4c",x"6b"),
  1055 => (x"9a",x"72",x"8a",x"c1"),
  1056 => (x"75",x"87",x"c5",x"02"),
  1057 => (x"87",x"ee",x"02",x"ac"),
  1058 => (x"d3",x"c1",x"1e",x"74"),
  1059 => (x"fe",x"fe",x"1e",x"d2"),
  1060 => (x"86",x"c8",x"87",x"ea"),
  1061 => (x"4d",x"26",x"48",x"74"),
  1062 => (x"4b",x"26",x"4c",x"26"),
  1063 => (x"5e",x"0e",x"4f",x"26"),
  1064 => (x"e4",x"f6",x"c0",x"0e"),
  1065 => (x"c0",x"4a",x"c0",x"c0"),
  1066 => (x"7a",x"ff",x"c3",x"49"),
  1067 => (x"c8",x"c3",x"81",x"c1"),
  1068 => (x"f4",x"04",x"a9",x"b7"),
  1069 => (x"0e",x"4f",x"26",x"87"),
  1070 => (x"5d",x"5c",x"5b",x"5e"),
  1071 => (x"c0",x"c0",x"c1",x"0e"),
  1072 => (x"4c",x"c0",x"c0",x"c0"),
  1073 => (x"c0",x"e4",x"f6",x"c0"),
  1074 => (x"d1",x"ff",x"4b",x"c0"),
  1075 => (x"df",x"f8",x"c4",x"87"),
  1076 => (x"c0",x"1e",x"c0",x"4d"),
  1077 => (x"f7",x"c1",x"f0",x"ff"),
  1078 => (x"87",x"ef",x"fc",x"1e"),
  1079 => (x"49",x"70",x"86",x"c8"),
  1080 => (x"c1",x"05",x"a9",x"c1"),
  1081 => (x"1e",x"71",x"87",x"c8"),
  1082 => (x"1e",x"d6",x"c5",x"c1"),
  1083 => (x"87",x"cc",x"fd",x"fe"),
  1084 => (x"ff",x"c3",x"86",x"c8"),
  1085 => (x"c0",x"1e",x"74",x"7b"),
  1086 => (x"e9",x"c1",x"f0",x"e1"),
  1087 => (x"87",x"cb",x"fc",x"1e"),
  1088 => (x"49",x"70",x"86",x"c8"),
  1089 => (x"d4",x"05",x"99",x"71"),
  1090 => (x"c1",x"1e",x"71",x"87"),
  1091 => (x"fe",x"1e",x"cc",x"c5"),
  1092 => (x"c8",x"87",x"e9",x"fc"),
  1093 => (x"7b",x"ff",x"c3",x"86"),
  1094 => (x"e7",x"c0",x"48",x"c1"),
  1095 => (x"c1",x"1e",x"71",x"87"),
  1096 => (x"fe",x"1e",x"e0",x"c5"),
  1097 => (x"c8",x"87",x"d5",x"fc"),
  1098 => (x"87",x"f2",x"fd",x"86"),
  1099 => (x"1e",x"71",x"87",x"cc"),
  1100 => (x"1e",x"ea",x"c5",x"c1"),
  1101 => (x"87",x"c4",x"fc",x"fe"),
  1102 => (x"8d",x"c1",x"86",x"c8"),
  1103 => (x"fe",x"05",x"9d",x"75"),
  1104 => (x"48",x"c0",x"87",x"cf"),
  1105 => (x"4c",x"26",x"4d",x"26"),
  1106 => (x"4f",x"26",x"4b",x"26"),
  1107 => (x"34",x"44",x"4d",x"43"),
  1108 => (x"64",x"25",x"20",x"31"),
  1109 => (x"4d",x"43",x"00",x"0a"),
  1110 => (x"20",x"35",x"35",x"44"),
  1111 => (x"00",x"0a",x"64",x"25"),
  1112 => (x"34",x"44",x"4d",x"43"),
  1113 => (x"64",x"25",x"20",x"31"),
  1114 => (x"4d",x"43",x"00",x"0a"),
  1115 => (x"20",x"35",x"35",x"44"),
  1116 => (x"00",x"0a",x"64",x"25"),
  1117 => (x"5c",x"5b",x"5e",x"0e"),
  1118 => (x"ff",x"c0",x"0e",x"5d"),
  1119 => (x"4d",x"c1",x"c1",x"f0"),
  1120 => (x"c0",x"e4",x"f6",x"c0"),
  1121 => (x"ff",x"c3",x"4b",x"c0"),
  1122 => (x"ee",x"c7",x"c1",x"7b"),
  1123 => (x"87",x"fb",x"cd",x"1e"),
  1124 => (x"4c",x"d3",x"86",x"c4"),
  1125 => (x"1e",x"75",x"1e",x"c0"),
  1126 => (x"c8",x"87",x"f0",x"f9"),
  1127 => (x"71",x"49",x"70",x"86"),
  1128 => (x"87",x"d3",x"05",x"99"),
  1129 => (x"c7",x"c1",x"1e",x"71"),
  1130 => (x"fa",x"fe",x"1e",x"d8"),
  1131 => (x"86",x"c8",x"87",x"ce"),
  1132 => (x"c1",x"7b",x"ff",x"c3"),
  1133 => (x"71",x"87",x"d9",x"48"),
  1134 => (x"e3",x"c7",x"c1",x"1e"),
  1135 => (x"fb",x"f9",x"fe",x"1e"),
  1136 => (x"fb",x"86",x"c8",x"87"),
  1137 => (x"8c",x"c1",x"87",x"d8"),
  1138 => (x"ff",x"05",x"9c",x"74"),
  1139 => (x"48",x"c0",x"87",x"c6"),
  1140 => (x"4c",x"26",x"4d",x"26"),
  1141 => (x"4f",x"26",x"4b",x"26"),
  1142 => (x"74",x"69",x"6e",x"69"),
  1143 => (x"0a",x"64",x"25",x"20"),
  1144 => (x"69",x"00",x"20",x"20"),
  1145 => (x"20",x"74",x"69",x"6e"),
  1146 => (x"20",x"0a",x"64",x"25"),
  1147 => (x"6d",x"43",x"00",x"20"),
  1148 => (x"6e",x"69",x"5f",x"64"),
  1149 => (x"00",x"0a",x"74",x"69"),
  1150 => (x"5c",x"5b",x"5e",x"0e"),
  1151 => (x"86",x"fc",x"0e",x"5d"),
  1152 => (x"c0",x"4d",x"ff",x"c3"),
  1153 => (x"c0",x"c0",x"e4",x"f6"),
  1154 => (x"87",x"d2",x"fa",x"4c"),
  1155 => (x"c0",x"1e",x"ea",x"c6"),
  1156 => (x"c8",x"c1",x"f0",x"e1"),
  1157 => (x"87",x"f3",x"f7",x"1e"),
  1158 => (x"4b",x"70",x"86",x"c8"),
  1159 => (x"cd",x"c1",x"1e",x"73"),
  1160 => (x"f8",x"fe",x"1e",x"ce"),
  1161 => (x"86",x"c8",x"87",x"d6"),
  1162 => (x"c0",x"02",x"ab",x"c1"),
  1163 => (x"c3",x"fd",x"87",x"c8"),
  1164 => (x"c2",x"48",x"c0",x"87"),
  1165 => (x"c3",x"f6",x"87",x"f7"),
  1166 => (x"73",x"4b",x"70",x"87"),
  1167 => (x"ff",x"ff",x"cf",x"49"),
  1168 => (x"a9",x"ea",x"c6",x"99"),
  1169 => (x"87",x"d4",x"c0",x"02"),
  1170 => (x"cb",x"c1",x"1e",x"73"),
  1171 => (x"f7",x"fe",x"1e",x"f7"),
  1172 => (x"86",x"c8",x"87",x"ea"),
  1173 => (x"c0",x"87",x"dd",x"fc"),
  1174 => (x"87",x"d1",x"c2",x"48"),
  1175 => (x"48",x"76",x"7c",x"75"),
  1176 => (x"f9",x"78",x"f1",x"c0"),
  1177 => (x"98",x"70",x"87",x"d1"),
  1178 => (x"87",x"dc",x"c1",x"02"),
  1179 => (x"ff",x"c0",x"1e",x"c0"),
  1180 => (x"1e",x"fa",x"c1",x"f0"),
  1181 => (x"c8",x"87",x"d4",x"f6"),
  1182 => (x"73",x"4b",x"70",x"86"),
  1183 => (x"fb",x"c0",x"05",x"9b"),
  1184 => (x"c1",x"1e",x"73",x"87"),
  1185 => (x"fe",x"1e",x"cc",x"cc"),
  1186 => (x"c8",x"87",x"f1",x"f6"),
  1187 => (x"6c",x"7c",x"75",x"86"),
  1188 => (x"73",x"9b",x"75",x"4b"),
  1189 => (x"d8",x"cc",x"c1",x"1e"),
  1190 => (x"df",x"f6",x"fe",x"1e"),
  1191 => (x"75",x"86",x"c8",x"87"),
  1192 => (x"75",x"7c",x"75",x"7c"),
  1193 => (x"73",x"7c",x"75",x"7c"),
  1194 => (x"99",x"c0",x"c1",x"49"),
  1195 => (x"c0",x"02",x"99",x"71"),
  1196 => (x"48",x"c1",x"87",x"c5"),
  1197 => (x"c0",x"87",x"f6",x"c0"),
  1198 => (x"87",x"f1",x"c0",x"48"),
  1199 => (x"cc",x"c1",x"1e",x"73"),
  1200 => (x"f5",x"fe",x"1e",x"e6"),
  1201 => (x"86",x"c8",x"87",x"f6"),
  1202 => (x"a8",x"c2",x"48",x"6e"),
  1203 => (x"87",x"cf",x"c0",x"05"),
  1204 => (x"1e",x"f2",x"cc",x"c1"),
  1205 => (x"87",x"e4",x"f5",x"fe"),
  1206 => (x"48",x"c0",x"86",x"c4"),
  1207 => (x"6e",x"87",x"ce",x"c0"),
  1208 => (x"c4",x"88",x"c1",x"48"),
  1209 => (x"05",x"6e",x"58",x"a6"),
  1210 => (x"c0",x"87",x"f8",x"fd"),
  1211 => (x"26",x"8e",x"fc",x"48"),
  1212 => (x"26",x"4c",x"26",x"4d"),
  1213 => (x"43",x"4f",x"26",x"4b"),
  1214 => (x"5f",x"38",x"44",x"4d"),
  1215 => (x"65",x"72",x"20",x"34"),
  1216 => (x"6e",x"6f",x"70",x"73"),
  1217 => (x"20",x"3a",x"65",x"73"),
  1218 => (x"00",x"0a",x"64",x"25"),
  1219 => (x"35",x"44",x"4d",x"43"),
  1220 => (x"64",x"25",x"20",x"38"),
  1221 => (x"00",x"20",x"20",x"0a"),
  1222 => (x"35",x"44",x"4d",x"43"),
  1223 => (x"20",x"32",x"5f",x"38"),
  1224 => (x"20",x"0a",x"64",x"25"),
  1225 => (x"4d",x"43",x"00",x"20"),
  1226 => (x"20",x"38",x"35",x"44"),
  1227 => (x"20",x"0a",x"64",x"25"),
  1228 => (x"44",x"53",x"00",x"20"),
  1229 => (x"49",x"20",x"43",x"48"),
  1230 => (x"69",x"74",x"69",x"6e"),
  1231 => (x"7a",x"69",x"6c",x"61"),
  1232 => (x"6f",x"69",x"74",x"61"),
  1233 => (x"72",x"65",x"20",x"6e"),
  1234 => (x"21",x"72",x"6f",x"72"),
  1235 => (x"6d",x"63",x"00",x"0a"),
  1236 => (x"4d",x"43",x"5f",x"64"),
  1237 => (x"72",x"20",x"38",x"44"),
  1238 => (x"6f",x"70",x"73",x"65"),
  1239 => (x"3a",x"65",x"73",x"6e"),
  1240 => (x"0a",x"64",x"25",x"20"),
  1241 => (x"5b",x"5e",x"0e",x"00"),
  1242 => (x"c0",x"0e",x"5d",x"5c"),
  1243 => (x"c0",x"c0",x"e4",x"f6"),
  1244 => (x"e4",x"f6",x"c0",x"4d"),
  1245 => (x"c1",x"4b",x"c4",x"c0"),
  1246 => (x"c1",x"48",x"f8",x"e0"),
  1247 => (x"e4",x"f6",x"c0",x"78"),
  1248 => (x"c0",x"48",x"c8",x"c0"),
  1249 => (x"4c",x"c7",x"78",x"e0"),
  1250 => (x"d1",x"f4",x"7b",x"c3"),
  1251 => (x"c3",x"7b",x"c2",x"87"),
  1252 => (x"1e",x"c0",x"7d",x"ff"),
  1253 => (x"c1",x"d0",x"e5",x"c0"),
  1254 => (x"ee",x"f1",x"1e",x"c0"),
  1255 => (x"c1",x"86",x"c8",x"87"),
  1256 => (x"c2",x"c0",x"05",x"a8"),
  1257 => (x"c2",x"4c",x"c1",x"87"),
  1258 => (x"c5",x"c0",x"05",x"ac"),
  1259 => (x"c0",x"48",x"c0",x"87"),
  1260 => (x"8c",x"c1",x"87",x"ee"),
  1261 => (x"ff",x"05",x"9c",x"74"),
  1262 => (x"fb",x"f8",x"87",x"ce"),
  1263 => (x"fc",x"e0",x"c1",x"87"),
  1264 => (x"f8",x"e0",x"c1",x"58"),
  1265 => (x"cd",x"c0",x"05",x"bf"),
  1266 => (x"c0",x"1e",x"c1",x"87"),
  1267 => (x"d0",x"c1",x"f0",x"ff"),
  1268 => (x"87",x"f7",x"f0",x"1e"),
  1269 => (x"ff",x"c3",x"86",x"c8"),
  1270 => (x"c3",x"7b",x"c3",x"7d"),
  1271 => (x"48",x"c1",x"7d",x"ff"),
  1272 => (x"4c",x"26",x"4d",x"26"),
  1273 => (x"4f",x"26",x"4b",x"26"),
  1274 => (x"26",x"48",x"c0",x"1e"),
  1275 => (x"5b",x"5e",x"0e",x"4f"),
  1276 => (x"fc",x"0e",x"5d",x"5c"),
  1277 => (x"4d",x"66",x"d8",x"86"),
  1278 => (x"c0",x"e4",x"f6",x"c0"),
  1279 => (x"48",x"76",x"4b",x"c0"),
  1280 => (x"1e",x"75",x"78",x"c0"),
  1281 => (x"c1",x"1e",x"66",x"d8"),
  1282 => (x"fe",x"1e",x"fb",x"d2"),
  1283 => (x"cc",x"87",x"ed",x"f0"),
  1284 => (x"7b",x"ff",x"c3",x"86"),
  1285 => (x"c0",x"e4",x"f6",x"c0"),
  1286 => (x"78",x"c2",x"48",x"c4"),
  1287 => (x"c0",x"e4",x"f6",x"c0"),
  1288 => (x"78",x"c1",x"48",x"c8"),
  1289 => (x"d4",x"7b",x"ff",x"c3"),
  1290 => (x"ff",x"c0",x"1e",x"66"),
  1291 => (x"1e",x"d1",x"c1",x"f0"),
  1292 => (x"c8",x"87",x"d8",x"ef"),
  1293 => (x"71",x"49",x"70",x"86"),
  1294 => (x"d2",x"c0",x"02",x"99"),
  1295 => (x"d8",x"1e",x"71",x"87"),
  1296 => (x"d2",x"c1",x"1e",x"66"),
  1297 => (x"ef",x"fe",x"1e",x"db"),
  1298 => (x"86",x"cc",x"87",x"f2"),
  1299 => (x"c5",x"87",x"c0",x"c1"),
  1300 => (x"4a",x"df",x"cd",x"ee"),
  1301 => (x"6b",x"7b",x"ff",x"c3"),
  1302 => (x"99",x"ff",x"c3",x"49"),
  1303 => (x"05",x"a9",x"fe",x"c3"),
  1304 => (x"c0",x"87",x"d9",x"c0"),
  1305 => (x"87",x"ef",x"eb",x"4c"),
  1306 => (x"85",x"c4",x"7d",x"70"),
  1307 => (x"c0",x"c2",x"84",x"c1"),
  1308 => (x"ff",x"04",x"ac",x"b7"),
  1309 => (x"4a",x"c1",x"87",x"ef"),
  1310 => (x"78",x"c1",x"48",x"76"),
  1311 => (x"9a",x"72",x"8a",x"c1"),
  1312 => (x"87",x"d0",x"ff",x"05"),
  1313 => (x"c0",x"7b",x"ff",x"c3"),
  1314 => (x"c4",x"c0",x"e4",x"f6"),
  1315 => (x"6e",x"78",x"c3",x"48"),
  1316 => (x"26",x"8e",x"fc",x"48"),
  1317 => (x"26",x"4c",x"26",x"4d"),
  1318 => (x"52",x"4f",x"26",x"4b"),
  1319 => (x"20",x"64",x"61",x"65"),
  1320 => (x"6d",x"6d",x"6f",x"63"),
  1321 => (x"20",x"64",x"6e",x"61"),
  1322 => (x"6c",x"69",x"61",x"66"),
  1323 => (x"61",x"20",x"64",x"65"),
  1324 => (x"64",x"25",x"20",x"74"),
  1325 => (x"64",x"25",x"28",x"20"),
  1326 => (x"73",x"00",x"0a",x"29"),
  1327 => (x"65",x"72",x"5f",x"64"),
  1328 => (x"73",x"5f",x"64",x"61"),
  1329 => (x"6f",x"74",x"63",x"65"),
  1330 => (x"64",x"25",x"20",x"72"),
  1331 => (x"64",x"25",x"20",x"2c"),
  1332 => (x"6f",x"47",x"00",x"0a"),
  1333 => (x"65",x"72",x"20",x"74"),
  1334 => (x"74",x"6c",x"75",x"73"),
  1335 => (x"20",x"64",x"25",x"20"),
  1336 => (x"fc",x"1e",x"00",x"0a"),
  1337 => (x"e8",x"f6",x"c0",x"86"),
  1338 => (x"69",x"49",x"c0",x"c0"),
  1339 => (x"98",x"c0",x"c4",x"48"),
  1340 => (x"6e",x"58",x"a6",x"c4"),
  1341 => (x"69",x"87",x"cc",x"05"),
  1342 => (x"98",x"c0",x"c4",x"48"),
  1343 => (x"6e",x"58",x"a6",x"c4"),
  1344 => (x"c8",x"87",x"f4",x"02"),
  1345 => (x"fc",x"48",x"79",x"66"),
  1346 => (x"0e",x"4f",x"26",x"8e"),
  1347 => (x"5d",x"5c",x"5b",x"5e"),
  1348 => (x"4c",x"66",x"d0",x"0e"),
  1349 => (x"4b",x"14",x"4d",x"c0"),
  1350 => (x"bb",x"83",x"c0",x"fe"),
  1351 => (x"c1",x"ff",x"1e",x"73"),
  1352 => (x"c1",x"86",x"c4",x"87"),
  1353 => (x"05",x"9b",x"73",x"85"),
  1354 => (x"48",x"75",x"87",x"ec"),
  1355 => (x"4c",x"26",x"4d",x"26"),
  1356 => (x"4f",x"26",x"4b",x"26"),
  1357 => (x"5c",x"5b",x"5e",x"0e"),
  1358 => (x"86",x"f8",x"0e",x"5d"),
  1359 => (x"d8",x"4b",x"66",x"dc"),
  1360 => (x"48",x"76",x"49",x"66"),
  1361 => (x"ab",x"b7",x"78",x"c0"),
  1362 => (x"87",x"cf",x"c1",x"06"),
  1363 => (x"32",x"c8",x"4a",x"11"),
  1364 => (x"b7",x"c0",x"8b",x"c1"),
  1365 => (x"87",x"c7",x"06",x"ab"),
  1366 => (x"a6",x"c8",x"48",x"11"),
  1367 => (x"c4",x"87",x"c5",x"58"),
  1368 => (x"78",x"c0",x"48",x"a6"),
  1369 => (x"c8",x"b2",x"66",x"c4"),
  1370 => (x"c0",x"8b",x"c1",x"32"),
  1371 => (x"c4",x"06",x"ab",x"b7"),
  1372 => (x"c2",x"4c",x"11",x"87"),
  1373 => (x"74",x"4c",x"c0",x"87"),
  1374 => (x"c1",x"32",x"c8",x"b2"),
  1375 => (x"ab",x"b7",x"c0",x"8b"),
  1376 => (x"11",x"87",x"c4",x"06"),
  1377 => (x"c0",x"87",x"c2",x"4d"),
  1378 => (x"72",x"b2",x"75",x"4d"),
  1379 => (x"c4",x"80",x"6e",x"48"),
  1380 => (x"8b",x"c1",x"58",x"a6"),
  1381 => (x"01",x"ab",x"b7",x"c0"),
  1382 => (x"6e",x"87",x"f1",x"fe"),
  1383 => (x"26",x"8e",x"f8",x"48"),
  1384 => (x"26",x"4c",x"26",x"4d"),
  1385 => (x"26",x"4f",x"26",x"4b"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
