
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"3b",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"38"),
    10 => (x"20",x"00",x"27",x"4f"),
    11 => (x"27",x"4e",x"00",x"00"),
    12 => (x"00",x"00",x"04",x"0e"),
    13 => (x"87",x"fd",x"00",x"0f"),
    14 => (x"4f",x"87",x"fd",x"00"),
    15 => (x"ff",x"86",x"fc",x"1e"),
    16 => (x"48",x"69",x"49",x"c0"),
    17 => (x"c4",x"98",x"c0",x"c4"),
    18 => (x"02",x"6e",x"58",x"a6"),
    19 => (x"66",x"c8",x"87",x"f4"),
    20 => (x"8e",x"fc",x"48",x"79"),
    21 => (x"5e",x"0e",x"4f",x"26"),
    22 => (x"0e",x"5d",x"5c",x"5b"),
    23 => (x"c0",x"4b",x"66",x"d0"),
    24 => (x"c3",x"49",x"13",x"4c"),
    25 => (x"99",x"71",x"99",x"ff"),
    26 => (x"71",x"87",x"dd",x"02"),
    27 => (x"4a",x"c0",x"ff",x"4d"),
    28 => (x"c0",x"c4",x"49",x"6a"),
    29 => (x"02",x"99",x"71",x"99"),
    30 => (x"7a",x"75",x"87",x"f6"),
    31 => (x"49",x"13",x"84",x"c1"),
    32 => (x"71",x"99",x"ff",x"c3"),
    33 => (x"87",x"e3",x"05",x"99"),
    34 => (x"4d",x"26",x"48",x"74"),
    35 => (x"4b",x"26",x"4c",x"26"),
    36 => (x"5e",x"0e",x"4f",x"26"),
    37 => (x"0e",x"5d",x"5c",x"5b"),
    38 => (x"f4",x"c0",x"86",x"e4"),
    39 => (x"a6",x"c4",x"4d",x"66"),
    40 => (x"c4",x"78",x"c0",x"48"),
    41 => (x"c0",x"78",x"c0",x"80"),
    42 => (x"bf",x"97",x"66",x"ec"),
    43 => (x"83",x"c0",x"fe",x"4b"),
    44 => (x"66",x"ec",x"c0",x"bb"),
    45 => (x"c0",x"80",x"c1",x"48"),
    46 => (x"73",x"58",x"a6",x"f0"),
    47 => (x"f7",x"c7",x"02",x"9b"),
    48 => (x"02",x"66",x"c8",x"87"),
    49 => (x"d0",x"87",x"c0",x"c7"),
    50 => (x"78",x"c0",x"48",x"a6"),
    51 => (x"78",x"c0",x"80",x"f8"),
    52 => (x"02",x"ab",x"f0",x"c0"),
    53 => (x"c1",x"87",x"ea",x"c2"),
    54 => (x"c2",x"02",x"ab",x"e3"),
    55 => (x"e4",x"c1",x"87",x"eb"),
    56 => (x"e2",x"c0",x"02",x"ab"),
    57 => (x"ab",x"ec",x"c1",x"87"),
    58 => (x"87",x"d5",x"c2",x"02"),
    59 => (x"02",x"ab",x"f0",x"c1"),
    60 => (x"f3",x"c1",x"87",x"dd"),
    61 => (x"87",x"df",x"02",x"ab"),
    62 => (x"02",x"ab",x"f5",x"c1"),
    63 => (x"f8",x"c1",x"87",x"c9"),
    64 => (x"87",x"cb",x"02",x"ab"),
    65 => (x"d0",x"87",x"e7",x"c2"),
    66 => (x"78",x"ca",x"48",x"a6"),
    67 => (x"d0",x"87",x"c2",x"c3"),
    68 => (x"78",x"d0",x"48",x"a6"),
    69 => (x"c0",x"87",x"fa",x"c2"),
    70 => (x"c4",x"48",x"66",x"f0"),
    71 => (x"a6",x"f4",x"c0",x"80"),
    72 => (x"66",x"f0",x"c0",x"58"),
    73 => (x"76",x"89",x"c4",x"49"),
    74 => (x"d4",x"78",x"69",x"48"),
    75 => (x"6e",x"78",x"ff",x"80"),
    76 => (x"fe",x"48",x"bf",x"97"),
    77 => (x"dc",x"b8",x"80",x"c0"),
    78 => (x"48",x"6e",x"58",x"a6"),
    79 => (x"a6",x"c4",x"80",x"c1"),
    80 => (x"5b",x"a6",x"d0",x"58"),
    81 => (x"c0",x"02",x"66",x"d8"),
    82 => (x"66",x"d8",x"87",x"e8"),
    83 => (x"d4",x"4b",x"6e",x"4c"),
    84 => (x"80",x"c1",x"48",x"66"),
    85 => (x"c0",x"58",x"a6",x"d8"),
    86 => (x"74",x"1e",x"66",x"f8"),
    87 => (x"c8",x"0f",x"75",x"1e"),
    88 => (x"05",x"a8",x"74",x"86"),
    89 => (x"4c",x"13",x"87",x"cc"),
    90 => (x"bc",x"84",x"c0",x"fe"),
    91 => (x"ff",x"05",x"9c",x"74"),
    92 => (x"66",x"cc",x"87",x"dd"),
    93 => (x"48",x"66",x"d4",x"4b"),
    94 => (x"c8",x"80",x"66",x"c4"),
    95 => (x"d0",x"c1",x"58",x"a6"),
    96 => (x"48",x"a6",x"c8",x"87"),
    97 => (x"c8",x"c1",x"78",x"c1"),
    98 => (x"66",x"f8",x"c0",x"87"),
    99 => (x"66",x"f4",x"c0",x"1e"),
   100 => (x"c0",x"80",x"c4",x"48"),
   101 => (x"c0",x"58",x"a6",x"f8"),
   102 => (x"c4",x"49",x"66",x"f4"),
   103 => (x"75",x"1e",x"69",x"89"),
   104 => (x"c4",x"86",x"c8",x"0f"),
   105 => (x"80",x"c1",x"48",x"66"),
   106 => (x"c0",x"58",x"a6",x"c8"),
   107 => (x"e5",x"c0",x"87",x"e3"),
   108 => (x"87",x"cb",x"02",x"ab"),
   109 => (x"1e",x"66",x"f8",x"c0"),
   110 => (x"75",x"1e",x"e5",x"c0"),
   111 => (x"c0",x"86",x"c8",x"0f"),
   112 => (x"73",x"1e",x"66",x"f8"),
   113 => (x"c8",x"0f",x"75",x"1e"),
   114 => (x"48",x"66",x"c4",x"86"),
   115 => (x"a6",x"c8",x"80",x"c1"),
   116 => (x"02",x"66",x"d0",x"58"),
   117 => (x"c0",x"87",x"c7",x"c3"),
   118 => (x"c4",x"48",x"66",x"f0"),
   119 => (x"a6",x"f4",x"c0",x"80"),
   120 => (x"66",x"f0",x"c0",x"58"),
   121 => (x"76",x"89",x"c4",x"49"),
   122 => (x"c1",x"78",x"69",x"48"),
   123 => (x"d8",x"05",x"ab",x"e4"),
   124 => (x"c0",x"48",x"6e",x"87"),
   125 => (x"d0",x"03",x"a8",x"b7"),
   126 => (x"1e",x"ed",x"c0",x"87"),
   127 => (x"c4",x"87",x"fd",x"f8"),
   128 => (x"c0",x"48",x"6e",x"86"),
   129 => (x"a6",x"c4",x"88",x"08"),
   130 => (x"c1",x"4a",x"6e",x"58"),
   131 => (x"cc",x"4c",x"e8",x"d8"),
   132 => (x"78",x"c0",x"48",x"a6"),
   133 => (x"87",x"ce",x"05",x"6e"),
   134 => (x"4c",x"e9",x"d8",x"c1"),
   135 => (x"48",x"e8",x"d8",x"c1"),
   136 => (x"c0",x"50",x"f0",x"c0"),
   137 => (x"02",x"6e",x"87",x"eb"),
   138 => (x"d0",x"87",x"e6",x"c0"),
   139 => (x"1e",x"72",x"4b",x"66"),
   140 => (x"4a",x"73",x"49",x"72"),
   141 => (x"26",x"87",x"da",x"c5"),
   142 => (x"81",x"c0",x"ce",x"4a"),
   143 => (x"1e",x"71",x"54",x"11"),
   144 => (x"4a",x"73",x"49",x"72"),
   145 => (x"70",x"87",x"ca",x"c5"),
   146 => (x"72",x"49",x"26",x"4a"),
   147 => (x"dd",x"ff",x"05",x"9a"),
   148 => (x"e8",x"d8",x"c1",x"87"),
   149 => (x"e3",x"c0",x"02",x"ac"),
   150 => (x"66",x"f8",x"c0",x"87"),
   151 => (x"97",x"8c",x"c1",x"1e"),
   152 => (x"c0",x"fe",x"49",x"6c"),
   153 => (x"1e",x"71",x"b9",x"81"),
   154 => (x"86",x"c8",x"0f",x"75"),
   155 => (x"c1",x"48",x"66",x"cc"),
   156 => (x"58",x"a6",x"d0",x"80"),
   157 => (x"ac",x"e8",x"d8",x"c1"),
   158 => (x"87",x"dd",x"ff",x"05"),
   159 => (x"c4",x"48",x"66",x"cc"),
   160 => (x"a6",x"c8",x"80",x"66"),
   161 => (x"c0",x"87",x"d7",x"58"),
   162 => (x"c7",x"05",x"ab",x"e5"),
   163 => (x"48",x"a6",x"c8",x"87"),
   164 => (x"87",x"ca",x"78",x"c1"),
   165 => (x"1e",x"66",x"f8",x"c0"),
   166 => (x"0f",x"75",x"1e",x"73"),
   167 => (x"ec",x"c0",x"86",x"c8"),
   168 => (x"4b",x"bf",x"97",x"66"),
   169 => (x"bb",x"83",x"c0",x"fe"),
   170 => (x"48",x"66",x"ec",x"c0"),
   171 => (x"f0",x"c0",x"80",x"c1"),
   172 => (x"9b",x"73",x"58",x"a6"),
   173 => (x"87",x"c9",x"f8",x"05"),
   174 => (x"e4",x"48",x"66",x"c4"),
   175 => (x"26",x"4d",x"26",x"8e"),
   176 => (x"26",x"4b",x"26",x"4c"),
   177 => (x"1e",x"c0",x"1e",x"4f"),
   178 => (x"d0",x"1e",x"fc",x"c0"),
   179 => (x"66",x"d0",x"1e",x"66"),
   180 => (x"87",x"fe",x"f6",x"1e"),
   181 => (x"4f",x"26",x"86",x"d0"),
   182 => (x"c0",x"1e",x"c0",x"1e"),
   183 => (x"a6",x"d0",x"1e",x"fc"),
   184 => (x"1e",x"66",x"d0",x"1e"),
   185 => (x"d0",x"87",x"eb",x"f6"),
   186 => (x"1e",x"4f",x"26",x"86"),
   187 => (x"48",x"76",x"86",x"f8"),
   188 => (x"c4",x"78",x"66",x"cc"),
   189 => (x"76",x"78",x"ff",x"80"),
   190 => (x"1e",x"ce",x"cd",x"1e"),
   191 => (x"dc",x"1e",x"a6",x"dc"),
   192 => (x"cd",x"f6",x"1e",x"66"),
   193 => (x"f8",x"86",x"d0",x"87"),
   194 => (x"1e",x"4f",x"26",x"8e"),
   195 => (x"48",x"76",x"86",x"f8"),
   196 => (x"c4",x"78",x"66",x"cc"),
   197 => (x"78",x"66",x"d0",x"80"),
   198 => (x"ce",x"cd",x"1e",x"76"),
   199 => (x"a6",x"e0",x"c0",x"1e"),
   200 => (x"66",x"e0",x"c0",x"1e"),
   201 => (x"87",x"ea",x"f5",x"1e"),
   202 => (x"8e",x"f8",x"86",x"d0"),
   203 => (x"f8",x"1e",x"4f",x"26"),
   204 => (x"cc",x"48",x"76",x"86"),
   205 => (x"80",x"c4",x"78",x"66"),
   206 => (x"1e",x"76",x"78",x"ff"),
   207 => (x"dc",x"1e",x"ce",x"cd"),
   208 => (x"66",x"dc",x"1e",x"66"),
   209 => (x"87",x"ca",x"f5",x"1e"),
   210 => (x"8e",x"f8",x"86",x"d0"),
   211 => (x"c8",x"1e",x"4f",x"26"),
   212 => (x"82",x"c4",x"4a",x"66"),
   213 => (x"e0",x"c0",x"02",x"6a"),
   214 => (x"c1",x"48",x"6a",x"87"),
   215 => (x"c8",x"7a",x"70",x"88"),
   216 => (x"71",x"49",x"bf",x"66"),
   217 => (x"c8",x"80",x"c1",x"48"),
   218 => (x"08",x"78",x"08",x"66"),
   219 => (x"51",x"66",x"c4",x"97"),
   220 => (x"c4",x"98",x"ff",x"c3"),
   221 => (x"c2",x"c0",x"48",x"66"),
   222 => (x"26",x"48",x"c0",x"87"),
   223 => (x"00",x"00",x"00",x"4f"),
   224 => (x"33",x"32",x"31",x"30"),
   225 => (x"37",x"36",x"35",x"34"),
   226 => (x"42",x"41",x"39",x"38"),
   227 => (x"46",x"45",x"44",x"43"),
   228 => (x"1e",x"73",x"1e",x"00"),
   229 => (x"c0",x"02",x"9a",x"72"),
   230 => (x"48",x"c0",x"87",x"e7"),
   231 => (x"a9",x"72",x"4b",x"c1"),
   232 => (x"72",x"87",x"d1",x"06"),
   233 => (x"87",x"c9",x"06",x"82"),
   234 => (x"a9",x"72",x"83",x"73"),
   235 => (x"c3",x"87",x"f4",x"01"),
   236 => (x"3a",x"b2",x"c1",x"87"),
   237 => (x"89",x"03",x"a9",x"72"),
   238 => (x"c1",x"07",x"80",x"73"),
   239 => (x"f3",x"05",x"2b",x"2a"),
   240 => (x"26",x"4b",x"26",x"87"),
   241 => (x"1e",x"75",x"1e",x"4f"),
   242 => (x"b7",x"71",x"4d",x"c4"),
   243 => (x"b9",x"ff",x"04",x"a1"),
   244 => (x"bd",x"c3",x"81",x"c1"),
   245 => (x"a2",x"b7",x"72",x"07"),
   246 => (x"c1",x"ba",x"ff",x"04"),
   247 => (x"07",x"bd",x"c1",x"82"),
   248 => (x"c1",x"87",x"ee",x"fe"),
   249 => (x"b8",x"ff",x"04",x"2d"),
   250 => (x"2d",x"07",x"80",x"c1"),
   251 => (x"c1",x"b9",x"ff",x"04"),
   252 => (x"4d",x"26",x"07",x"81"),
   253 => (x"72",x"1e",x"4f",x"26"),
   254 => (x"11",x"48",x"12",x"1e"),
   255 => (x"88",x"87",x"c4",x"02"),
   256 => (x"26",x"87",x"f6",x"02"),
   257 => (x"1e",x"4f",x"26",x"4a"),
   258 => (x"48",x"bf",x"c8",x"ff"),
   259 => (x"5e",x"0e",x"4f",x"26"),
   260 => (x"0e",x"5d",x"5c",x"5b"),
   261 => (x"c1",x"86",x"dc",x"ff"),
   262 => (x"c3",x"48",x"fc",x"d8"),
   263 => (x"c1",x"78",x"c0",x"f9"),
   264 => (x"c3",x"48",x"f8",x"d8"),
   265 => (x"48",x"78",x"f0",x"f9"),
   266 => (x"78",x"c0",x"f9",x"c3"),
   267 => (x"48",x"f4",x"f9",x"c3"),
   268 => (x"80",x"c4",x"78",x"c0"),
   269 => (x"f9",x"c3",x"78",x"c2"),
   270 => (x"e8",x"c0",x"48",x"fc"),
   271 => (x"c3",x"1e",x"71",x"78"),
   272 => (x"c0",x"49",x"c0",x"fa"),
   273 => (x"20",x"48",x"d4",x"f6"),
   274 => (x"20",x"41",x"20",x"41"),
   275 => (x"20",x"41",x"20",x"41"),
   276 => (x"20",x"41",x"20",x"41"),
   277 => (x"10",x"51",x"10",x"41"),
   278 => (x"26",x"51",x"10",x"51"),
   279 => (x"c3",x"1e",x"71",x"49"),
   280 => (x"c0",x"49",x"e0",x"fa"),
   281 => (x"20",x"48",x"f4",x"f6"),
   282 => (x"20",x"41",x"20",x"41"),
   283 => (x"20",x"41",x"20",x"41"),
   284 => (x"20",x"41",x"20",x"41"),
   285 => (x"10",x"51",x"10",x"41"),
   286 => (x"26",x"51",x"10",x"51"),
   287 => (x"f4",x"f5",x"c1",x"49"),
   288 => (x"c0",x"78",x"ca",x"48"),
   289 => (x"f9",x"1e",x"d4",x"f7"),
   290 => (x"86",x"c4",x"87",x"ce"),
   291 => (x"1e",x"d8",x"f7",x"c0"),
   292 => (x"c4",x"87",x"c5",x"f9"),
   293 => (x"c8",x"f8",x"c0",x"86"),
   294 => (x"87",x"fc",x"f8",x"1e"),
   295 => (x"ef",x"c0",x"86",x"c4"),
   296 => (x"d4",x"02",x"bf",x"f8"),
   297 => (x"c0",x"f0",x"c0",x"87"),
   298 => (x"87",x"ec",x"f8",x"1e"),
   299 => (x"f0",x"c0",x"86",x"c4"),
   300 => (x"e3",x"f8",x"1e",x"ec"),
   301 => (x"d2",x"86",x"c4",x"87"),
   302 => (x"f0",x"f0",x"c0",x"87"),
   303 => (x"87",x"d8",x"f8",x"1e"),
   304 => (x"f1",x"c0",x"86",x"c4"),
   305 => (x"cf",x"f8",x"1e",x"e0"),
   306 => (x"c0",x"86",x"c4",x"87"),
   307 => (x"1e",x"bf",x"fc",x"ef"),
   308 => (x"1e",x"cc",x"f8",x"c0"),
   309 => (x"c8",x"87",x"c1",x"f8"),
   310 => (x"e8",x"f8",x"c3",x"86"),
   311 => (x"bf",x"c8",x"ff",x"48"),
   312 => (x"48",x"a6",x"c8",x"78"),
   313 => (x"ef",x"c0",x"78",x"c1"),
   314 => (x"c0",x"48",x"bf",x"fc"),
   315 => (x"c9",x"06",x"a8",x"b7"),
   316 => (x"a6",x"cc",x"87",x"dd"),
   317 => (x"58",x"a6",x"d4",x"48"),
   318 => (x"a6",x"dc",x"80",x"c8"),
   319 => (x"48",x"a6",x"dc",x"58"),
   320 => (x"c1",x"58",x"a6",x"c8"),
   321 => (x"c1",x"48",x"c8",x"d9"),
   322 => (x"d9",x"c1",x"50",x"c1"),
   323 => (x"78",x"c0",x"48",x"c4"),
   324 => (x"97",x"c8",x"d9",x"c1"),
   325 => (x"c0",x"fe",x"49",x"bf"),
   326 => (x"c1",x"c1",x"b9",x"81"),
   327 => (x"c7",x"c0",x"02",x"a9"),
   328 => (x"c0",x"48",x"76",x"87"),
   329 => (x"87",x"c4",x"c0",x"78"),
   330 => (x"78",x"c1",x"48",x"76"),
   331 => (x"bf",x"c4",x"d9",x"c1"),
   332 => (x"c1",x"b0",x"6e",x"48"),
   333 => (x"c1",x"58",x"c8",x"d9"),
   334 => (x"c1",x"48",x"cc",x"d9"),
   335 => (x"a6",x"dc",x"50",x"c2"),
   336 => (x"c4",x"78",x"c2",x"48"),
   337 => (x"c3",x"78",x"c3",x"80"),
   338 => (x"c0",x"49",x"c0",x"fb"),
   339 => (x"20",x"48",x"c4",x"f2"),
   340 => (x"20",x"41",x"20",x"41"),
   341 => (x"20",x"41",x"20",x"41"),
   342 => (x"20",x"41",x"20",x"41"),
   343 => (x"10",x"51",x"10",x"41"),
   344 => (x"d4",x"51",x"10",x"51"),
   345 => (x"78",x"c1",x"48",x"a6"),
   346 => (x"1e",x"c0",x"fb",x"c3"),
   347 => (x"1e",x"e0",x"fa",x"c3"),
   348 => (x"87",x"ed",x"c0",x"c1"),
   349 => (x"98",x"70",x"86",x"c8"),
   350 => (x"87",x"c5",x"c0",x"05"),
   351 => (x"c2",x"c0",x"49",x"c1"),
   352 => (x"c1",x"49",x"c0",x"87"),
   353 => (x"dc",x"59",x"c8",x"d9"),
   354 => (x"b7",x"c3",x"48",x"66"),
   355 => (x"ef",x"c0",x"03",x"a8"),
   356 => (x"49",x"66",x"dc",x"87"),
   357 => (x"71",x"91",x"b7",x"c5"),
   358 => (x"d0",x"88",x"c3",x"48"),
   359 => (x"66",x"d0",x"58",x"a6"),
   360 => (x"c0",x"1e",x"c3",x"1e"),
   361 => (x"c0",x"1e",x"66",x"e4"),
   362 => (x"cc",x"87",x"ce",x"fc"),
   363 => (x"48",x"66",x"dc",x"86"),
   364 => (x"e0",x"c0",x"80",x"c1"),
   365 => (x"66",x"dc",x"58",x"a6"),
   366 => (x"a8",x"b7",x"c3",x"48"),
   367 => (x"87",x"d1",x"ff",x"04"),
   368 => (x"c0",x"1e",x"66",x"cc"),
   369 => (x"c1",x"1e",x"66",x"e0"),
   370 => (x"c1",x"1e",x"d8",x"dc"),
   371 => (x"c0",x"1e",x"d0",x"d9"),
   372 => (x"d0",x"87",x"f8",x"fb"),
   373 => (x"f8",x"d8",x"c1",x"86"),
   374 => (x"d8",x"c1",x"4c",x"bf"),
   375 => (x"4b",x"bf",x"bf",x"f8"),
   376 => (x"49",x"73",x"1e",x"72"),
   377 => (x"bf",x"f8",x"d8",x"c1"),
   378 => (x"a1",x"f0",x"c0",x"48"),
   379 => (x"71",x"41",x"20",x"4a"),
   380 => (x"f8",x"ff",x"05",x"aa"),
   381 => (x"74",x"4a",x"26",x"87"),
   382 => (x"c4",x"80",x"c8",x"48"),
   383 => (x"49",x"74",x"58",x"a6"),
   384 => (x"79",x"c5",x"81",x"cc"),
   385 => (x"85",x"cc",x"4d",x"73"),
   386 => (x"7b",x"6c",x"7d",x"69"),
   387 => (x"fa",x"d6",x"1e",x"73"),
   388 => (x"73",x"86",x"c4",x"87"),
   389 => (x"69",x"81",x"c4",x"49"),
   390 => (x"87",x"e7",x"c0",x"05"),
   391 => (x"81",x"c8",x"49",x"73"),
   392 => (x"1e",x"71",x"7d",x"c6"),
   393 => (x"1e",x"bf",x"66",x"c4"),
   394 => (x"87",x"df",x"f8",x"c0"),
   395 => (x"d8",x"c1",x"86",x"c8"),
   396 => (x"7b",x"bf",x"bf",x"f8"),
   397 => (x"1e",x"ca",x"1e",x"75"),
   398 => (x"f9",x"c0",x"1e",x"6d"),
   399 => (x"86",x"cc",x"87",x"fb"),
   400 => (x"6c",x"87",x"d9",x"c0"),
   401 => (x"72",x"1e",x"71",x"49"),
   402 => (x"48",x"49",x"74",x"1e"),
   403 => (x"4a",x"a1",x"f0",x"c0"),
   404 => (x"aa",x"71",x"41",x"20"),
   405 => (x"87",x"f8",x"ff",x"05"),
   406 => (x"49",x"26",x"4a",x"26"),
   407 => (x"c1",x"c1",x"48",x"76"),
   408 => (x"cc",x"d9",x"c1",x"50"),
   409 => (x"fe",x"49",x"bf",x"97"),
   410 => (x"c1",x"b9",x"81",x"c0"),
   411 => (x"04",x"a9",x"b7",x"c1"),
   412 => (x"97",x"87",x"ed",x"c1"),
   413 => (x"c3",x"c1",x"4b",x"6e"),
   414 => (x"fe",x"49",x"73",x"1e"),
   415 => (x"71",x"b9",x"81",x"c0"),
   416 => (x"f1",x"fb",x"c0",x"1e"),
   417 => (x"d4",x"86",x"c8",x"87"),
   418 => (x"c0",x"05",x"a8",x"66"),
   419 => (x"66",x"d8",x"87",x"f9"),
   420 => (x"c0",x"1e",x"c0",x"1e"),
   421 => (x"c8",x"87",x"f4",x"f6"),
   422 => (x"c3",x"1e",x"71",x"86"),
   423 => (x"c0",x"49",x"c0",x"fb"),
   424 => (x"20",x"48",x"e4",x"f1"),
   425 => (x"20",x"41",x"20",x"41"),
   426 => (x"20",x"41",x"20",x"41"),
   427 => (x"20",x"41",x"20",x"41"),
   428 => (x"10",x"51",x"10",x"41"),
   429 => (x"26",x"51",x"10",x"51"),
   430 => (x"a6",x"e0",x"c0",x"49"),
   431 => (x"78",x"66",x"c8",x"48"),
   432 => (x"48",x"c0",x"d9",x"c1"),
   433 => (x"c1",x"78",x"66",x"c8"),
   434 => (x"fe",x"4a",x"73",x"83"),
   435 => (x"c1",x"ba",x"82",x"c0"),
   436 => (x"bf",x"97",x"cc",x"d9"),
   437 => (x"81",x"c0",x"fe",x"49"),
   438 => (x"aa",x"b7",x"71",x"b9"),
   439 => (x"87",x"d6",x"fe",x"06"),
   440 => (x"48",x"66",x"e0",x"c0"),
   441 => (x"90",x"b7",x"66",x"dc"),
   442 => (x"58",x"a6",x"e4",x"c0"),
   443 => (x"1e",x"72",x"1e",x"71"),
   444 => (x"49",x"66",x"e8",x"c0"),
   445 => (x"f3",x"4a",x"66",x"d4"),
   446 => (x"4a",x"26",x"87",x"cb"),
   447 => (x"e0",x"c0",x"49",x"26"),
   448 => (x"e0",x"c0",x"58",x"a6"),
   449 => (x"66",x"cc",x"49",x"66"),
   450 => (x"91",x"b7",x"c7",x"89"),
   451 => (x"66",x"dc",x"48",x"71"),
   452 => (x"a6",x"e4",x"c0",x"88"),
   453 => (x"bf",x"66",x"c4",x"58"),
   454 => (x"c1",x"82",x"ca",x"4a"),
   455 => (x"bf",x"97",x"c8",x"d9"),
   456 => (x"81",x"c0",x"fe",x"49"),
   457 => (x"a9",x"c1",x"c1",x"b9"),
   458 => (x"87",x"ce",x"c0",x"05"),
   459 => (x"48",x"72",x"8a",x"c1"),
   460 => (x"bf",x"c0",x"d9",x"c1"),
   461 => (x"08",x"66",x"c4",x"88"),
   462 => (x"66",x"c8",x"08",x"78"),
   463 => (x"cc",x"80",x"c1",x"48"),
   464 => (x"66",x"c8",x"58",x"a6"),
   465 => (x"fc",x"ef",x"c0",x"48"),
   466 => (x"06",x"a8",x"b7",x"bf"),
   467 => (x"c3",x"87",x"f4",x"f6"),
   468 => (x"ff",x"48",x"ec",x"f8"),
   469 => (x"c0",x"78",x"bf",x"c8"),
   470 => (x"ed",x"1e",x"fc",x"f8"),
   471 => (x"86",x"c4",x"87",x"fa"),
   472 => (x"1e",x"cc",x"f9",x"c0"),
   473 => (x"c4",x"87",x"f1",x"ed"),
   474 => (x"d0",x"f9",x"c0",x"86"),
   475 => (x"87",x"e8",x"ed",x"1e"),
   476 => (x"fa",x"c0",x"86",x"c4"),
   477 => (x"df",x"ed",x"1e",x"c8"),
   478 => (x"c1",x"86",x"c4",x"87"),
   479 => (x"1e",x"bf",x"c0",x"d9"),
   480 => (x"1e",x"cc",x"fa",x"c0"),
   481 => (x"c8",x"87",x"d1",x"ed"),
   482 => (x"c0",x"1e",x"c5",x"86"),
   483 => (x"ed",x"1e",x"e8",x"fa"),
   484 => (x"86",x"c8",x"87",x"c6"),
   485 => (x"bf",x"c4",x"d9",x"c1"),
   486 => (x"c4",x"fb",x"c0",x"1e"),
   487 => (x"87",x"f8",x"ec",x"1e"),
   488 => (x"1e",x"c1",x"86",x"c8"),
   489 => (x"1e",x"e0",x"fb",x"c0"),
   490 => (x"c8",x"87",x"ed",x"ec"),
   491 => (x"c8",x"d9",x"c1",x"86"),
   492 => (x"fe",x"49",x"bf",x"97"),
   493 => (x"71",x"b9",x"81",x"c0"),
   494 => (x"fc",x"fb",x"c0",x"1e"),
   495 => (x"87",x"d8",x"ec",x"1e"),
   496 => (x"c1",x"c1",x"86",x"c8"),
   497 => (x"d8",x"fc",x"c0",x"1e"),
   498 => (x"87",x"cc",x"ec",x"1e"),
   499 => (x"d9",x"c1",x"86",x"c8"),
   500 => (x"49",x"bf",x"97",x"cc"),
   501 => (x"b9",x"81",x"c0",x"fe"),
   502 => (x"fc",x"c0",x"1e",x"71"),
   503 => (x"f7",x"eb",x"1e",x"f4"),
   504 => (x"c1",x"86",x"c8",x"87"),
   505 => (x"fd",x"c0",x"1e",x"c2"),
   506 => (x"eb",x"eb",x"1e",x"d0"),
   507 => (x"c1",x"86",x"c8",x"87"),
   508 => (x"1e",x"bf",x"f0",x"d9"),
   509 => (x"1e",x"ec",x"fd",x"c0"),
   510 => (x"c8",x"87",x"dd",x"eb"),
   511 => (x"c0",x"1e",x"c7",x"86"),
   512 => (x"eb",x"1e",x"c8",x"fe"),
   513 => (x"86",x"c8",x"87",x"d2"),
   514 => (x"bf",x"f4",x"f5",x"c1"),
   515 => (x"e4",x"fe",x"c0",x"1e"),
   516 => (x"87",x"c4",x"eb",x"1e"),
   517 => (x"ff",x"c0",x"86",x"c8"),
   518 => (x"fb",x"ea",x"1e",x"c0"),
   519 => (x"c0",x"86",x"c4",x"87"),
   520 => (x"ea",x"1e",x"ec",x"ff"),
   521 => (x"86",x"c4",x"87",x"f2"),
   522 => (x"bf",x"f8",x"d8",x"c1"),
   523 => (x"ff",x"c0",x"1e",x"bf"),
   524 => (x"e3",x"ea",x"1e",x"f8"),
   525 => (x"c1",x"86",x"c8",x"87"),
   526 => (x"ea",x"1e",x"d4",x"c0"),
   527 => (x"86",x"c4",x"87",x"da"),
   528 => (x"bf",x"f8",x"d8",x"c1"),
   529 => (x"69",x"81",x"c4",x"49"),
   530 => (x"c8",x"c1",x"c1",x"1e"),
   531 => (x"87",x"c8",x"ea",x"1e"),
   532 => (x"1e",x"c0",x"86",x"c8"),
   533 => (x"1e",x"e4",x"c1",x"c1"),
   534 => (x"c8",x"87",x"fd",x"e9"),
   535 => (x"f8",x"d8",x"c1",x"86"),
   536 => (x"81",x"c8",x"49",x"bf"),
   537 => (x"c2",x"c1",x"1e",x"69"),
   538 => (x"eb",x"e9",x"1e",x"c0"),
   539 => (x"c2",x"86",x"c8",x"87"),
   540 => (x"dc",x"c2",x"c1",x"1e"),
   541 => (x"87",x"e0",x"e9",x"1e"),
   542 => (x"d8",x"c1",x"86",x"c8"),
   543 => (x"cc",x"49",x"bf",x"f8"),
   544 => (x"c1",x"1e",x"69",x"81"),
   545 => (x"e9",x"1e",x"f8",x"c2"),
   546 => (x"86",x"c8",x"87",x"ce"),
   547 => (x"c3",x"c1",x"1e",x"d1"),
   548 => (x"c3",x"e9",x"1e",x"d4"),
   549 => (x"c1",x"86",x"c8",x"87"),
   550 => (x"49",x"bf",x"f8",x"d8"),
   551 => (x"1e",x"71",x"81",x"d0"),
   552 => (x"1e",x"f0",x"c3",x"c1"),
   553 => (x"c8",x"87",x"f1",x"e8"),
   554 => (x"cc",x"c4",x"c1",x"86"),
   555 => (x"87",x"e8",x"e8",x"1e"),
   556 => (x"c5",x"c1",x"86",x"c4"),
   557 => (x"df",x"e8",x"1e",x"c4"),
   558 => (x"c1",x"86",x"c4",x"87"),
   559 => (x"bf",x"bf",x"fc",x"d8"),
   560 => (x"d8",x"c5",x"c1",x"1e"),
   561 => (x"87",x"d0",x"e8",x"1e"),
   562 => (x"c5",x"c1",x"86",x"c8"),
   563 => (x"c7",x"e8",x"1e",x"f4"),
   564 => (x"c1",x"86",x"c4",x"87"),
   565 => (x"49",x"bf",x"fc",x"d8"),
   566 => (x"1e",x"69",x"81",x"c4"),
   567 => (x"1e",x"f4",x"c6",x"c1"),
   568 => (x"c8",x"87",x"f5",x"e7"),
   569 => (x"c1",x"1e",x"c0",x"86"),
   570 => (x"e7",x"1e",x"d0",x"c7"),
   571 => (x"86",x"c8",x"87",x"ea"),
   572 => (x"bf",x"fc",x"d8",x"c1"),
   573 => (x"69",x"81",x"c8",x"49"),
   574 => (x"ec",x"c7",x"c1",x"1e"),
   575 => (x"87",x"d8",x"e7",x"1e"),
   576 => (x"1e",x"c1",x"86",x"c8"),
   577 => (x"1e",x"c8",x"c8",x"c1"),
   578 => (x"c8",x"87",x"cd",x"e7"),
   579 => (x"fc",x"d8",x"c1",x"86"),
   580 => (x"81",x"cc",x"49",x"bf"),
   581 => (x"c8",x"c1",x"1e",x"69"),
   582 => (x"fb",x"e6",x"1e",x"e4"),
   583 => (x"d2",x"86",x"c8",x"87"),
   584 => (x"c0",x"c9",x"c1",x"1e"),
   585 => (x"87",x"f0",x"e6",x"1e"),
   586 => (x"d8",x"c1",x"86",x"c8"),
   587 => (x"d0",x"49",x"bf",x"fc"),
   588 => (x"c1",x"1e",x"71",x"81"),
   589 => (x"e6",x"1e",x"dc",x"c9"),
   590 => (x"86",x"c8",x"87",x"de"),
   591 => (x"1e",x"f8",x"c9",x"c1"),
   592 => (x"c4",x"87",x"d5",x"e6"),
   593 => (x"1e",x"66",x"dc",x"86"),
   594 => (x"1e",x"f0",x"ca",x"c1"),
   595 => (x"c8",x"87",x"c9",x"e6"),
   596 => (x"c1",x"1e",x"c5",x"86"),
   597 => (x"e5",x"1e",x"cc",x"cb"),
   598 => (x"86",x"c8",x"87",x"fe"),
   599 => (x"1e",x"66",x"e0",x"c0"),
   600 => (x"1e",x"e8",x"cb",x"c1"),
   601 => (x"c8",x"87",x"f1",x"e5"),
   602 => (x"c1",x"1e",x"cd",x"86"),
   603 => (x"e5",x"1e",x"c4",x"cc"),
   604 => (x"86",x"c8",x"87",x"e6"),
   605 => (x"c1",x"1e",x"66",x"cc"),
   606 => (x"e5",x"1e",x"e0",x"cc"),
   607 => (x"86",x"c8",x"87",x"da"),
   608 => (x"cc",x"c1",x"1e",x"c7"),
   609 => (x"cf",x"e5",x"1e",x"fc"),
   610 => (x"d4",x"86",x"c8",x"87"),
   611 => (x"cd",x"c1",x"1e",x"66"),
   612 => (x"c3",x"e5",x"1e",x"d8"),
   613 => (x"c1",x"86",x"c8",x"87"),
   614 => (x"f4",x"cd",x"c1",x"1e"),
   615 => (x"87",x"f8",x"e4",x"1e"),
   616 => (x"fa",x"c3",x"86",x"c8"),
   617 => (x"ce",x"c1",x"1e",x"e0"),
   618 => (x"eb",x"e4",x"1e",x"d0"),
   619 => (x"c1",x"86",x"c8",x"87"),
   620 => (x"e4",x"1e",x"ec",x"ce"),
   621 => (x"86",x"c4",x"87",x"e2"),
   622 => (x"1e",x"c0",x"fb",x"c3"),
   623 => (x"1e",x"e4",x"cf",x"c1"),
   624 => (x"c8",x"87",x"d5",x"e4"),
   625 => (x"c0",x"d0",x"c1",x"86"),
   626 => (x"87",x"cc",x"e4",x"1e"),
   627 => (x"d0",x"c1",x"86",x"c4"),
   628 => (x"c3",x"e4",x"1e",x"f8"),
   629 => (x"c3",x"86",x"c4",x"87"),
   630 => (x"49",x"bf",x"ec",x"f8"),
   631 => (x"bf",x"e8",x"f8",x"c3"),
   632 => (x"f4",x"f8",x"c3",x"89"),
   633 => (x"c1",x"1e",x"71",x"59"),
   634 => (x"e3",x"1e",x"fc",x"d0"),
   635 => (x"86",x"c8",x"87",x"ea"),
   636 => (x"bf",x"f0",x"f8",x"c3"),
   637 => (x"b7",x"f8",x"c1",x"48"),
   638 => (x"db",x"c0",x"03",x"a8"),
   639 => (x"e4",x"f2",x"c0",x"87"),
   640 => (x"87",x"d4",x"e3",x"1e"),
   641 => (x"f3",x"c0",x"86",x"c4"),
   642 => (x"cb",x"e3",x"1e",x"dc"),
   643 => (x"c0",x"86",x"c4",x"87"),
   644 => (x"e3",x"1e",x"fc",x"f3"),
   645 => (x"86",x"c4",x"87",x"c2"),
   646 => (x"bf",x"f0",x"f8",x"c3"),
   647 => (x"cf",x"4a",x"71",x"49"),
   648 => (x"71",x"92",x"b7",x"e8"),
   649 => (x"72",x"1e",x"72",x"1e"),
   650 => (x"fc",x"ef",x"c0",x"49"),
   651 => (x"d4",x"e6",x"4a",x"bf"),
   652 => (x"26",x"4a",x"26",x"87"),
   653 => (x"f8",x"f8",x"c3",x"49"),
   654 => (x"fc",x"ef",x"c0",x"58"),
   655 => (x"4b",x"72",x"4a",x"bf"),
   656 => (x"93",x"b7",x"e8",x"cf"),
   657 => (x"1e",x"72",x"1e",x"71"),
   658 => (x"e5",x"4a",x"09",x"73"),
   659 => (x"4a",x"26",x"87",x"f7"),
   660 => (x"f8",x"c3",x"49",x"26"),
   661 => (x"f9",x"c8",x"58",x"fc"),
   662 => (x"1e",x"71",x"92",x"b7"),
   663 => (x"09",x"72",x"1e",x"72"),
   664 => (x"87",x"e1",x"e5",x"4a"),
   665 => (x"49",x"26",x"4a",x"26"),
   666 => (x"58",x"c0",x"f9",x"c3"),
   667 => (x"1e",x"c0",x"f4",x"c0"),
   668 => (x"c4",x"87",x"e5",x"e1"),
   669 => (x"f4",x"f8",x"c3",x"86"),
   670 => (x"f4",x"c0",x"1e",x"bf"),
   671 => (x"d7",x"e1",x"1e",x"f0"),
   672 => (x"c0",x"86",x"c8",x"87"),
   673 => (x"e1",x"1e",x"f8",x"f4"),
   674 => (x"86",x"c4",x"87",x"ce"),
   675 => (x"bf",x"f8",x"f8",x"c3"),
   676 => (x"e8",x"f5",x"c0",x"1e"),
   677 => (x"87",x"c0",x"e1",x"1e"),
   678 => (x"f8",x"c3",x"86",x"c8"),
   679 => (x"c0",x"1e",x"bf",x"fc"),
   680 => (x"e0",x"1e",x"f0",x"f5"),
   681 => (x"86",x"c8",x"87",x"f2"),
   682 => (x"1e",x"d0",x"f6",x"c0"),
   683 => (x"c4",x"87",x"e9",x"e0"),
   684 => (x"ff",x"48",x"c0",x"86"),
   685 => (x"4d",x"26",x"8e",x"dc"),
   686 => (x"4b",x"26",x"4c",x"26"),
   687 => (x"c1",x"1e",x"4f",x"26"),
   688 => (x"c1",x"48",x"c8",x"d9"),
   689 => (x"d9",x"c1",x"50",x"c1"),
   690 => (x"78",x"c0",x"48",x"c4"),
   691 => (x"c1",x"1e",x"4f",x"26"),
   692 => (x"bf",x"97",x"c8",x"d9"),
   693 => (x"81",x"c0",x"fe",x"49"),
   694 => (x"a9",x"c1",x"c1",x"b9"),
   695 => (x"87",x"c5",x"c0",x"02"),
   696 => (x"c2",x"c0",x"49",x"c0"),
   697 => (x"c1",x"49",x"c1",x"87"),
   698 => (x"48",x"bf",x"c4",x"d9"),
   699 => (x"d9",x"c1",x"b0",x"71"),
   700 => (x"d9",x"c1",x"58",x"c8"),
   701 => (x"c2",x"c1",x"48",x"cc"),
   702 => (x"0e",x"4f",x"26",x"50"),
   703 => (x"5d",x"5c",x"5b",x"5e"),
   704 => (x"d4",x"86",x"fc",x"0e"),
   705 => (x"4b",x"6d",x"4d",x"66"),
   706 => (x"d8",x"c1",x"49",x"73"),
   707 => (x"c0",x"48",x"bf",x"f8"),
   708 => (x"20",x"4a",x"a1",x"f0"),
   709 => (x"05",x"aa",x"71",x"41"),
   710 => (x"75",x"87",x"f8",x"ff"),
   711 => (x"c4",x"80",x"c8",x"48"),
   712 => (x"49",x"75",x"58",x"a6"),
   713 => (x"79",x"c5",x"81",x"cc"),
   714 => (x"84",x"cc",x"4c",x"73"),
   715 => (x"7b",x"6d",x"7c",x"c5"),
   716 => (x"bf",x"f8",x"d8",x"c1"),
   717 => (x"87",x"c6",x"c0",x"02"),
   718 => (x"bf",x"f8",x"d8",x"c1"),
   719 => (x"d8",x"c1",x"7b",x"bf"),
   720 => (x"cc",x"49",x"bf",x"f8"),
   721 => (x"c1",x"1e",x"71",x"81"),
   722 => (x"1e",x"bf",x"c0",x"d9"),
   723 => (x"e5",x"c0",x"1e",x"ca"),
   724 => (x"86",x"cc",x"87",x"e7"),
   725 => (x"81",x"c4",x"49",x"73"),
   726 => (x"e7",x"c0",x"05",x"69"),
   727 => (x"c8",x"49",x"73",x"87"),
   728 => (x"71",x"7c",x"c6",x"81"),
   729 => (x"bf",x"66",x"c4",x"1e"),
   730 => (x"de",x"e3",x"c0",x"1e"),
   731 => (x"c1",x"86",x"c8",x"87"),
   732 => (x"bf",x"bf",x"f8",x"d8"),
   733 => (x"ca",x"1e",x"74",x"7b"),
   734 => (x"c0",x"1e",x"6c",x"1e"),
   735 => (x"cc",x"87",x"fa",x"e4"),
   736 => (x"87",x"d5",x"c0",x"86"),
   737 => (x"1e",x"71",x"49",x"6d"),
   738 => (x"c0",x"48",x"49",x"75"),
   739 => (x"20",x"4a",x"a1",x"f0"),
   740 => (x"05",x"aa",x"71",x"41"),
   741 => (x"26",x"87",x"f8",x"ff"),
   742 => (x"26",x"8e",x"fc",x"49"),
   743 => (x"26",x"4c",x"26",x"4d"),
   744 => (x"1e",x"4f",x"26",x"4b"),
   745 => (x"4a",x"bf",x"66",x"c4"),
   746 => (x"d9",x"c1",x"82",x"ca"),
   747 => (x"49",x"bf",x"97",x"c8"),
   748 => (x"b9",x"81",x"c0",x"fe"),
   749 => (x"05",x"a9",x"c1",x"c1"),
   750 => (x"c1",x"87",x"ce",x"c0"),
   751 => (x"c1",x"48",x"72",x"8a"),
   752 => (x"88",x"bf",x"c0",x"d9"),
   753 => (x"78",x"08",x"66",x"c4"),
   754 => (x"1e",x"4f",x"26",x"08"),
   755 => (x"bf",x"f8",x"d8",x"c1"),
   756 => (x"87",x"c9",x"c0",x"02"),
   757 => (x"c1",x"48",x"66",x"c4"),
   758 => (x"bf",x"bf",x"f8",x"d8"),
   759 => (x"f8",x"d8",x"c1",x"78"),
   760 => (x"81",x"cc",x"49",x"bf"),
   761 => (x"d9",x"c1",x"1e",x"71"),
   762 => (x"ca",x"1e",x"bf",x"c0"),
   763 => (x"c8",x"e3",x"c0",x"1e"),
   764 => (x"26",x"86",x"cc",x"87"),
   765 => (x"00",x"00",x"00",x"4f"),
   766 => (x"00",x"00",x"00",x"00"),
   767 => (x"00",x"00",x"61",x"a8"),
   768 => (x"67",x"6f",x"72",x"50"),
   769 => (x"20",x"6d",x"61",x"72"),
   770 => (x"70",x"6d",x"6f",x"63"),
   771 => (x"64",x"65",x"6c",x"69"),
   772 => (x"74",x"69",x"77",x"20"),
   773 => (x"72",x"27",x"20",x"68"),
   774 => (x"73",x"69",x"67",x"65"),
   775 => (x"27",x"72",x"65",x"74"),
   776 => (x"74",x"74",x"61",x"20"),
   777 => (x"75",x"62",x"69",x"72"),
   778 => (x"00",x"0a",x"65",x"74"),
   779 => (x"00",x"00",x"00",x"0a"),
   780 => (x"67",x"6f",x"72",x"50"),
   781 => (x"20",x"6d",x"61",x"72"),
   782 => (x"70",x"6d",x"6f",x"63"),
   783 => (x"64",x"65",x"6c",x"69"),
   784 => (x"74",x"69",x"77",x"20"),
   785 => (x"74",x"75",x"6f",x"68"),
   786 => (x"65",x"72",x"27",x"20"),
   787 => (x"74",x"73",x"69",x"67"),
   788 => (x"20",x"27",x"72",x"65"),
   789 => (x"72",x"74",x"74",x"61"),
   790 => (x"74",x"75",x"62",x"69"),
   791 => (x"00",x"00",x"0a",x"65"),
   792 => (x"00",x"00",x"00",x"0a"),
   793 => (x"59",x"52",x"48",x"44"),
   794 => (x"4e",x"4f",x"54",x"53"),
   795 => (x"52",x"50",x"20",x"45"),
   796 => (x"41",x"52",x"47",x"4f"),
   797 => (x"33",x"20",x"2c",x"4d"),
   798 => (x"20",x"44",x"52",x"27"),
   799 => (x"49",x"52",x"54",x"53"),
   800 => (x"00",x"00",x"47",x"4e"),
   801 => (x"59",x"52",x"48",x"44"),
   802 => (x"4e",x"4f",x"54",x"53"),
   803 => (x"52",x"50",x"20",x"45"),
   804 => (x"41",x"52",x"47",x"4f"),
   805 => (x"32",x"20",x"2c",x"4d"),
   806 => (x"20",x"44",x"4e",x"27"),
   807 => (x"49",x"52",x"54",x"53"),
   808 => (x"00",x"00",x"47",x"4e"),
   809 => (x"73",x"61",x"65",x"4d"),
   810 => (x"64",x"65",x"72",x"75"),
   811 => (x"6d",x"69",x"74",x"20"),
   812 => (x"6f",x"74",x"20",x"65"),
   813 => (x"6d",x"73",x"20",x"6f"),
   814 => (x"20",x"6c",x"6c",x"61"),
   815 => (x"6f",x"20",x"6f",x"74"),
   816 => (x"69",x"61",x"74",x"62"),
   817 => (x"65",x"6d",x"20",x"6e"),
   818 => (x"6e",x"69",x"6e",x"61"),
   819 => (x"6c",x"75",x"66",x"67"),
   820 => (x"73",x"65",x"72",x"20"),
   821 => (x"73",x"74",x"6c",x"75"),
   822 => (x"00",x"00",x"00",x"0a"),
   823 => (x"61",x"65",x"6c",x"50"),
   824 => (x"69",x"20",x"65",x"73"),
   825 => (x"65",x"72",x"63",x"6e"),
   826 => (x"20",x"65",x"73",x"61"),
   827 => (x"62",x"6d",x"75",x"6e"),
   828 => (x"6f",x"20",x"72",x"65"),
   829 => (x"75",x"72",x"20",x"66"),
   830 => (x"00",x"0a",x"73",x"6e"),
   831 => (x"00",x"00",x"00",x"0a"),
   832 => (x"72",x"63",x"69",x"4d"),
   833 => (x"63",x"65",x"73",x"6f"),
   834 => (x"73",x"64",x"6e",x"6f"),
   835 => (x"72",x"6f",x"66",x"20"),
   836 => (x"65",x"6e",x"6f",x"20"),
   837 => (x"6e",x"75",x"72",x"20"),
   838 => (x"72",x"68",x"74",x"20"),
   839 => (x"68",x"67",x"75",x"6f"),
   840 => (x"72",x"68",x"44",x"20"),
   841 => (x"6f",x"74",x"73",x"79"),
   842 => (x"20",x"3a",x"65",x"6e"),
   843 => (x"00",x"00",x"00",x"00"),
   844 => (x"0a",x"20",x"64",x"25"),
   845 => (x"00",x"00",x"00",x"00"),
   846 => (x"79",x"72",x"68",x"44"),
   847 => (x"6e",x"6f",x"74",x"73"),
   848 => (x"70",x"20",x"73",x"65"),
   849 => (x"53",x"20",x"72",x"65"),
   850 => (x"6e",x"6f",x"63",x"65"),
   851 => (x"20",x"20",x"3a",x"64"),
   852 => (x"20",x"20",x"20",x"20"),
   853 => (x"20",x"20",x"20",x"20"),
   854 => (x"20",x"20",x"20",x"20"),
   855 => (x"20",x"20",x"20",x"20"),
   856 => (x"20",x"20",x"20",x"20"),
   857 => (x"00",x"00",x"00",x"00"),
   858 => (x"0a",x"20",x"64",x"25"),
   859 => (x"00",x"00",x"00",x"00"),
   860 => (x"20",x"58",x"41",x"56"),
   861 => (x"53",x"50",x"49",x"4d"),
   862 => (x"74",x"61",x"72",x"20"),
   863 => (x"20",x"67",x"6e",x"69"),
   864 => (x"30",x"31",x"20",x"2a"),
   865 => (x"3d",x"20",x"30",x"30"),
   866 => (x"20",x"64",x"25",x"20"),
   867 => (x"00",x"00",x"00",x"0a"),
   868 => (x"00",x"00",x"00",x"0a"),
   869 => (x"59",x"52",x"48",x"44"),
   870 => (x"4e",x"4f",x"54",x"53"),
   871 => (x"52",x"50",x"20",x"45"),
   872 => (x"41",x"52",x"47",x"4f"),
   873 => (x"53",x"20",x"2c",x"4d"),
   874 => (x"20",x"45",x"4d",x"4f"),
   875 => (x"49",x"52",x"54",x"53"),
   876 => (x"00",x"00",x"47",x"4e"),
   877 => (x"59",x"52",x"48",x"44"),
   878 => (x"4e",x"4f",x"54",x"53"),
   879 => (x"52",x"50",x"20",x"45"),
   880 => (x"41",x"52",x"47",x"4f"),
   881 => (x"31",x"20",x"2c",x"4d"),
   882 => (x"20",x"54",x"53",x"27"),
   883 => (x"49",x"52",x"54",x"53"),
   884 => (x"00",x"00",x"47",x"4e"),
   885 => (x"00",x"00",x"00",x"0a"),
   886 => (x"79",x"72",x"68",x"44"),
   887 => (x"6e",x"6f",x"74",x"73"),
   888 => (x"65",x"42",x"20",x"65"),
   889 => (x"6d",x"68",x"63",x"6e"),
   890 => (x"2c",x"6b",x"72",x"61"),
   891 => (x"72",x"65",x"56",x"20"),
   892 => (x"6e",x"6f",x"69",x"73"),
   893 => (x"31",x"2e",x"32",x"20"),
   894 => (x"61",x"4c",x"28",x"20"),
   895 => (x"61",x"75",x"67",x"6e"),
   896 => (x"20",x"3a",x"65",x"67"),
   897 => (x"00",x"0a",x"29",x"43"),
   898 => (x"00",x"00",x"00",x"0a"),
   899 => (x"63",x"65",x"78",x"45"),
   900 => (x"6f",x"69",x"74",x"75"),
   901 => (x"74",x"73",x"20",x"6e"),
   902 => (x"73",x"74",x"72",x"61"),
   903 => (x"64",x"25",x"20",x"2c"),
   904 => (x"6e",x"75",x"72",x"20"),
   905 => (x"68",x"74",x"20",x"73"),
   906 => (x"67",x"75",x"6f",x"72"),
   907 => (x"68",x"44",x"20",x"68"),
   908 => (x"74",x"73",x"79",x"72"),
   909 => (x"0a",x"65",x"6e",x"6f"),
   910 => (x"00",x"00",x"00",x"00"),
   911 => (x"63",x"65",x"78",x"45"),
   912 => (x"6f",x"69",x"74",x"75"),
   913 => (x"6e",x"65",x"20",x"6e"),
   914 => (x"00",x"0a",x"73",x"64"),
   915 => (x"00",x"00",x"00",x"0a"),
   916 => (x"61",x"6e",x"69",x"46"),
   917 => (x"61",x"76",x"20",x"6c"),
   918 => (x"73",x"65",x"75",x"6c"),
   919 => (x"20",x"66",x"6f",x"20"),
   920 => (x"20",x"65",x"68",x"74"),
   921 => (x"69",x"72",x"61",x"76"),
   922 => (x"65",x"6c",x"62",x"61"),
   923 => (x"73",x"75",x"20",x"73"),
   924 => (x"69",x"20",x"64",x"65"),
   925 => (x"68",x"74",x"20",x"6e"),
   926 => (x"65",x"62",x"20",x"65"),
   927 => (x"6d",x"68",x"63",x"6e"),
   928 => (x"3a",x"6b",x"72",x"61"),
   929 => (x"00",x"00",x"00",x"0a"),
   930 => (x"00",x"00",x"00",x"0a"),
   931 => (x"5f",x"74",x"6e",x"49"),
   932 => (x"62",x"6f",x"6c",x"47"),
   933 => (x"20",x"20",x"20",x"3a"),
   934 => (x"20",x"20",x"20",x"20"),
   935 => (x"20",x"20",x"20",x"20"),
   936 => (x"0a",x"64",x"25",x"20"),
   937 => (x"00",x"00",x"00",x"00"),
   938 => (x"20",x"20",x"20",x"20"),
   939 => (x"20",x"20",x"20",x"20"),
   940 => (x"75",x"6f",x"68",x"73"),
   941 => (x"62",x"20",x"64",x"6c"),
   942 => (x"20",x"20",x"3a",x"65"),
   943 => (x"0a",x"64",x"25",x"20"),
   944 => (x"00",x"00",x"00",x"00"),
   945 => (x"6c",x"6f",x"6f",x"42"),
   946 => (x"6f",x"6c",x"47",x"5f"),
   947 => (x"20",x"20",x"3a",x"62"),
   948 => (x"20",x"20",x"20",x"20"),
   949 => (x"20",x"20",x"20",x"20"),
   950 => (x"0a",x"64",x"25",x"20"),
   951 => (x"00",x"00",x"00",x"00"),
   952 => (x"20",x"20",x"20",x"20"),
   953 => (x"20",x"20",x"20",x"20"),
   954 => (x"75",x"6f",x"68",x"73"),
   955 => (x"62",x"20",x"64",x"6c"),
   956 => (x"20",x"20",x"3a",x"65"),
   957 => (x"0a",x"64",x"25",x"20"),
   958 => (x"00",x"00",x"00",x"00"),
   959 => (x"31",x"5f",x"68",x"43"),
   960 => (x"6f",x"6c",x"47",x"5f"),
   961 => (x"20",x"20",x"3a",x"62"),
   962 => (x"20",x"20",x"20",x"20"),
   963 => (x"20",x"20",x"20",x"20"),
   964 => (x"0a",x"63",x"25",x"20"),
   965 => (x"00",x"00",x"00",x"00"),
   966 => (x"20",x"20",x"20",x"20"),
   967 => (x"20",x"20",x"20",x"20"),
   968 => (x"75",x"6f",x"68",x"73"),
   969 => (x"62",x"20",x"64",x"6c"),
   970 => (x"20",x"20",x"3a",x"65"),
   971 => (x"0a",x"63",x"25",x"20"),
   972 => (x"00",x"00",x"00",x"00"),
   973 => (x"32",x"5f",x"68",x"43"),
   974 => (x"6f",x"6c",x"47",x"5f"),
   975 => (x"20",x"20",x"3a",x"62"),
   976 => (x"20",x"20",x"20",x"20"),
   977 => (x"20",x"20",x"20",x"20"),
   978 => (x"0a",x"63",x"25",x"20"),
   979 => (x"00",x"00",x"00",x"00"),
   980 => (x"20",x"20",x"20",x"20"),
   981 => (x"20",x"20",x"20",x"20"),
   982 => (x"75",x"6f",x"68",x"73"),
   983 => (x"62",x"20",x"64",x"6c"),
   984 => (x"20",x"20",x"3a",x"65"),
   985 => (x"0a",x"63",x"25",x"20"),
   986 => (x"00",x"00",x"00",x"00"),
   987 => (x"5f",x"72",x"72",x"41"),
   988 => (x"6c",x"47",x"5f",x"31"),
   989 => (x"38",x"5b",x"62",x"6f"),
   990 => (x"20",x"20",x"3a",x"5d"),
   991 => (x"20",x"20",x"20",x"20"),
   992 => (x"0a",x"64",x"25",x"20"),
   993 => (x"00",x"00",x"00",x"00"),
   994 => (x"20",x"20",x"20",x"20"),
   995 => (x"20",x"20",x"20",x"20"),
   996 => (x"75",x"6f",x"68",x"73"),
   997 => (x"62",x"20",x"64",x"6c"),
   998 => (x"20",x"20",x"3a",x"65"),
   999 => (x"0a",x"64",x"25",x"20"),
  1000 => (x"00",x"00",x"00",x"00"),
  1001 => (x"5f",x"72",x"72",x"41"),
  1002 => (x"6c",x"47",x"5f",x"32"),
  1003 => (x"38",x"5b",x"62",x"6f"),
  1004 => (x"5d",x"37",x"5b",x"5d"),
  1005 => (x"20",x"20",x"20",x"3a"),
  1006 => (x"0a",x"64",x"25",x"20"),
  1007 => (x"00",x"00",x"00",x"00"),
  1008 => (x"20",x"20",x"20",x"20"),
  1009 => (x"20",x"20",x"20",x"20"),
  1010 => (x"75",x"6f",x"68",x"73"),
  1011 => (x"62",x"20",x"64",x"6c"),
  1012 => (x"20",x"20",x"3a",x"65"),
  1013 => (x"6d",x"75",x"4e",x"20"),
  1014 => (x"5f",x"72",x"65",x"62"),
  1015 => (x"52",x"5f",x"66",x"4f"),
  1016 => (x"20",x"73",x"6e",x"75"),
  1017 => (x"30",x"31",x"20",x"2b"),
  1018 => (x"00",x"00",x"00",x"0a"),
  1019 => (x"5f",x"72",x"74",x"50"),
  1020 => (x"62",x"6f",x"6c",x"47"),
  1021 => (x"00",x"0a",x"3e",x"2d"),
  1022 => (x"74",x"50",x"20",x"20"),
  1023 => (x"6f",x"43",x"5f",x"72"),
  1024 => (x"20",x"3a",x"70",x"6d"),
  1025 => (x"20",x"20",x"20",x"20"),
  1026 => (x"20",x"20",x"20",x"20"),
  1027 => (x"0a",x"64",x"25",x"20"),
  1028 => (x"00",x"00",x"00",x"00"),
  1029 => (x"20",x"20",x"20",x"20"),
  1030 => (x"20",x"20",x"20",x"20"),
  1031 => (x"75",x"6f",x"68",x"73"),
  1032 => (x"62",x"20",x"64",x"6c"),
  1033 => (x"20",x"20",x"3a",x"65"),
  1034 => (x"6d",x"69",x"28",x"20"),
  1035 => (x"6d",x"65",x"6c",x"70"),
  1036 => (x"61",x"74",x"6e",x"65"),
  1037 => (x"6e",x"6f",x"69",x"74"),
  1038 => (x"70",x"65",x"64",x"2d"),
  1039 => (x"65",x"64",x"6e",x"65"),
  1040 => (x"0a",x"29",x"74",x"6e"),
  1041 => (x"00",x"00",x"00",x"00"),
  1042 => (x"69",x"44",x"20",x"20"),
  1043 => (x"3a",x"72",x"63",x"73"),
  1044 => (x"20",x"20",x"20",x"20"),
  1045 => (x"20",x"20",x"20",x"20"),
  1046 => (x"20",x"20",x"20",x"20"),
  1047 => (x"0a",x"64",x"25",x"20"),
  1048 => (x"00",x"00",x"00",x"00"),
  1049 => (x"20",x"20",x"20",x"20"),
  1050 => (x"20",x"20",x"20",x"20"),
  1051 => (x"75",x"6f",x"68",x"73"),
  1052 => (x"62",x"20",x"64",x"6c"),
  1053 => (x"20",x"20",x"3a",x"65"),
  1054 => (x"0a",x"64",x"25",x"20"),
  1055 => (x"00",x"00",x"00",x"00"),
  1056 => (x"6e",x"45",x"20",x"20"),
  1057 => (x"43",x"5f",x"6d",x"75"),
  1058 => (x"3a",x"70",x"6d",x"6f"),
  1059 => (x"20",x"20",x"20",x"20"),
  1060 => (x"20",x"20",x"20",x"20"),
  1061 => (x"0a",x"64",x"25",x"20"),
  1062 => (x"00",x"00",x"00",x"00"),
  1063 => (x"20",x"20",x"20",x"20"),
  1064 => (x"20",x"20",x"20",x"20"),
  1065 => (x"75",x"6f",x"68",x"73"),
  1066 => (x"62",x"20",x"64",x"6c"),
  1067 => (x"20",x"20",x"3a",x"65"),
  1068 => (x"0a",x"64",x"25",x"20"),
  1069 => (x"00",x"00",x"00",x"00"),
  1070 => (x"6e",x"49",x"20",x"20"),
  1071 => (x"6f",x"43",x"5f",x"74"),
  1072 => (x"20",x"3a",x"70",x"6d"),
  1073 => (x"20",x"20",x"20",x"20"),
  1074 => (x"20",x"20",x"20",x"20"),
  1075 => (x"0a",x"64",x"25",x"20"),
  1076 => (x"00",x"00",x"00",x"00"),
  1077 => (x"20",x"20",x"20",x"20"),
  1078 => (x"20",x"20",x"20",x"20"),
  1079 => (x"75",x"6f",x"68",x"73"),
  1080 => (x"62",x"20",x"64",x"6c"),
  1081 => (x"20",x"20",x"3a",x"65"),
  1082 => (x"0a",x"64",x"25",x"20"),
  1083 => (x"00",x"00",x"00",x"00"),
  1084 => (x"74",x"53",x"20",x"20"),
  1085 => (x"6f",x"43",x"5f",x"72"),
  1086 => (x"20",x"3a",x"70",x"6d"),
  1087 => (x"20",x"20",x"20",x"20"),
  1088 => (x"20",x"20",x"20",x"20"),
  1089 => (x"0a",x"73",x"25",x"20"),
  1090 => (x"00",x"00",x"00",x"00"),
  1091 => (x"20",x"20",x"20",x"20"),
  1092 => (x"20",x"20",x"20",x"20"),
  1093 => (x"75",x"6f",x"68",x"73"),
  1094 => (x"62",x"20",x"64",x"6c"),
  1095 => (x"20",x"20",x"3a",x"65"),
  1096 => (x"52",x"48",x"44",x"20"),
  1097 => (x"4f",x"54",x"53",x"59"),
  1098 => (x"50",x"20",x"45",x"4e"),
  1099 => (x"52",x"47",x"4f",x"52"),
  1100 => (x"20",x"2c",x"4d",x"41"),
  1101 => (x"45",x"4d",x"4f",x"53"),
  1102 => (x"52",x"54",x"53",x"20"),
  1103 => (x"0a",x"47",x"4e",x"49"),
  1104 => (x"00",x"00",x"00",x"00"),
  1105 => (x"74",x"78",x"65",x"4e"),
  1106 => (x"72",x"74",x"50",x"5f"),
  1107 => (x"6f",x"6c",x"47",x"5f"),
  1108 => (x"0a",x"3e",x"2d",x"62"),
  1109 => (x"00",x"00",x"00",x"00"),
  1110 => (x"74",x"50",x"20",x"20"),
  1111 => (x"6f",x"43",x"5f",x"72"),
  1112 => (x"20",x"3a",x"70",x"6d"),
  1113 => (x"20",x"20",x"20",x"20"),
  1114 => (x"20",x"20",x"20",x"20"),
  1115 => (x"0a",x"64",x"25",x"20"),
  1116 => (x"00",x"00",x"00",x"00"),
  1117 => (x"20",x"20",x"20",x"20"),
  1118 => (x"20",x"20",x"20",x"20"),
  1119 => (x"75",x"6f",x"68",x"73"),
  1120 => (x"62",x"20",x"64",x"6c"),
  1121 => (x"20",x"20",x"3a",x"65"),
  1122 => (x"6d",x"69",x"28",x"20"),
  1123 => (x"6d",x"65",x"6c",x"70"),
  1124 => (x"61",x"74",x"6e",x"65"),
  1125 => (x"6e",x"6f",x"69",x"74"),
  1126 => (x"70",x"65",x"64",x"2d"),
  1127 => (x"65",x"64",x"6e",x"65"),
  1128 => (x"2c",x"29",x"74",x"6e"),
  1129 => (x"6d",x"61",x"73",x"20"),
  1130 => (x"73",x"61",x"20",x"65"),
  1131 => (x"6f",x"62",x"61",x"20"),
  1132 => (x"00",x"0a",x"65",x"76"),
  1133 => (x"69",x"44",x"20",x"20"),
  1134 => (x"3a",x"72",x"63",x"73"),
  1135 => (x"20",x"20",x"20",x"20"),
  1136 => (x"20",x"20",x"20",x"20"),
  1137 => (x"20",x"20",x"20",x"20"),
  1138 => (x"0a",x"64",x"25",x"20"),
  1139 => (x"00",x"00",x"00",x"00"),
  1140 => (x"20",x"20",x"20",x"20"),
  1141 => (x"20",x"20",x"20",x"20"),
  1142 => (x"75",x"6f",x"68",x"73"),
  1143 => (x"62",x"20",x"64",x"6c"),
  1144 => (x"20",x"20",x"3a",x"65"),
  1145 => (x"0a",x"64",x"25",x"20"),
  1146 => (x"00",x"00",x"00",x"00"),
  1147 => (x"6e",x"45",x"20",x"20"),
  1148 => (x"43",x"5f",x"6d",x"75"),
  1149 => (x"3a",x"70",x"6d",x"6f"),
  1150 => (x"20",x"20",x"20",x"20"),
  1151 => (x"20",x"20",x"20",x"20"),
  1152 => (x"0a",x"64",x"25",x"20"),
  1153 => (x"00",x"00",x"00",x"00"),
  1154 => (x"20",x"20",x"20",x"20"),
  1155 => (x"20",x"20",x"20",x"20"),
  1156 => (x"75",x"6f",x"68",x"73"),
  1157 => (x"62",x"20",x"64",x"6c"),
  1158 => (x"20",x"20",x"3a",x"65"),
  1159 => (x"0a",x"64",x"25",x"20"),
  1160 => (x"00",x"00",x"00",x"00"),
  1161 => (x"6e",x"49",x"20",x"20"),
  1162 => (x"6f",x"43",x"5f",x"74"),
  1163 => (x"20",x"3a",x"70",x"6d"),
  1164 => (x"20",x"20",x"20",x"20"),
  1165 => (x"20",x"20",x"20",x"20"),
  1166 => (x"0a",x"64",x"25",x"20"),
  1167 => (x"00",x"00",x"00",x"00"),
  1168 => (x"20",x"20",x"20",x"20"),
  1169 => (x"20",x"20",x"20",x"20"),
  1170 => (x"75",x"6f",x"68",x"73"),
  1171 => (x"62",x"20",x"64",x"6c"),
  1172 => (x"20",x"20",x"3a",x"65"),
  1173 => (x"0a",x"64",x"25",x"20"),
  1174 => (x"00",x"00",x"00",x"00"),
  1175 => (x"74",x"53",x"20",x"20"),
  1176 => (x"6f",x"43",x"5f",x"72"),
  1177 => (x"20",x"3a",x"70",x"6d"),
  1178 => (x"20",x"20",x"20",x"20"),
  1179 => (x"20",x"20",x"20",x"20"),
  1180 => (x"0a",x"73",x"25",x"20"),
  1181 => (x"00",x"00",x"00",x"00"),
  1182 => (x"20",x"20",x"20",x"20"),
  1183 => (x"20",x"20",x"20",x"20"),
  1184 => (x"75",x"6f",x"68",x"73"),
  1185 => (x"62",x"20",x"64",x"6c"),
  1186 => (x"20",x"20",x"3a",x"65"),
  1187 => (x"52",x"48",x"44",x"20"),
  1188 => (x"4f",x"54",x"53",x"59"),
  1189 => (x"50",x"20",x"45",x"4e"),
  1190 => (x"52",x"47",x"4f",x"52"),
  1191 => (x"20",x"2c",x"4d",x"41"),
  1192 => (x"45",x"4d",x"4f",x"53"),
  1193 => (x"52",x"54",x"53",x"20"),
  1194 => (x"0a",x"47",x"4e",x"49"),
  1195 => (x"00",x"00",x"00",x"00"),
  1196 => (x"5f",x"74",x"6e",x"49"),
  1197 => (x"6f",x"4c",x"5f",x"31"),
  1198 => (x"20",x"20",x"3a",x"63"),
  1199 => (x"20",x"20",x"20",x"20"),
  1200 => (x"20",x"20",x"20",x"20"),
  1201 => (x"0a",x"64",x"25",x"20"),
  1202 => (x"00",x"00",x"00",x"00"),
  1203 => (x"20",x"20",x"20",x"20"),
  1204 => (x"20",x"20",x"20",x"20"),
  1205 => (x"75",x"6f",x"68",x"73"),
  1206 => (x"62",x"20",x"64",x"6c"),
  1207 => (x"20",x"20",x"3a",x"65"),
  1208 => (x"0a",x"64",x"25",x"20"),
  1209 => (x"00",x"00",x"00",x"00"),
  1210 => (x"5f",x"74",x"6e",x"49"),
  1211 => (x"6f",x"4c",x"5f",x"32"),
  1212 => (x"20",x"20",x"3a",x"63"),
  1213 => (x"20",x"20",x"20",x"20"),
  1214 => (x"20",x"20",x"20",x"20"),
  1215 => (x"0a",x"64",x"25",x"20"),
  1216 => (x"00",x"00",x"00",x"00"),
  1217 => (x"20",x"20",x"20",x"20"),
  1218 => (x"20",x"20",x"20",x"20"),
  1219 => (x"75",x"6f",x"68",x"73"),
  1220 => (x"62",x"20",x"64",x"6c"),
  1221 => (x"20",x"20",x"3a",x"65"),
  1222 => (x"0a",x"64",x"25",x"20"),
  1223 => (x"00",x"00",x"00",x"00"),
  1224 => (x"5f",x"74",x"6e",x"49"),
  1225 => (x"6f",x"4c",x"5f",x"33"),
  1226 => (x"20",x"20",x"3a",x"63"),
  1227 => (x"20",x"20",x"20",x"20"),
  1228 => (x"20",x"20",x"20",x"20"),
  1229 => (x"0a",x"64",x"25",x"20"),
  1230 => (x"00",x"00",x"00",x"00"),
  1231 => (x"20",x"20",x"20",x"20"),
  1232 => (x"20",x"20",x"20",x"20"),
  1233 => (x"75",x"6f",x"68",x"73"),
  1234 => (x"62",x"20",x"64",x"6c"),
  1235 => (x"20",x"20",x"3a",x"65"),
  1236 => (x"0a",x"64",x"25",x"20"),
  1237 => (x"00",x"00",x"00",x"00"),
  1238 => (x"6d",x"75",x"6e",x"45"),
  1239 => (x"63",x"6f",x"4c",x"5f"),
  1240 => (x"20",x"20",x"20",x"3a"),
  1241 => (x"20",x"20",x"20",x"20"),
  1242 => (x"20",x"20",x"20",x"20"),
  1243 => (x"0a",x"64",x"25",x"20"),
  1244 => (x"00",x"00",x"00",x"00"),
  1245 => (x"20",x"20",x"20",x"20"),
  1246 => (x"20",x"20",x"20",x"20"),
  1247 => (x"75",x"6f",x"68",x"73"),
  1248 => (x"62",x"20",x"64",x"6c"),
  1249 => (x"20",x"20",x"3a",x"65"),
  1250 => (x"0a",x"64",x"25",x"20"),
  1251 => (x"00",x"00",x"00",x"00"),
  1252 => (x"5f",x"72",x"74",x"53"),
  1253 => (x"6f",x"4c",x"5f",x"31"),
  1254 => (x"20",x"20",x"3a",x"63"),
  1255 => (x"20",x"20",x"20",x"20"),
  1256 => (x"20",x"20",x"20",x"20"),
  1257 => (x"0a",x"73",x"25",x"20"),
  1258 => (x"00",x"00",x"00",x"00"),
  1259 => (x"20",x"20",x"20",x"20"),
  1260 => (x"20",x"20",x"20",x"20"),
  1261 => (x"75",x"6f",x"68",x"73"),
  1262 => (x"62",x"20",x"64",x"6c"),
  1263 => (x"20",x"20",x"3a",x"65"),
  1264 => (x"52",x"48",x"44",x"20"),
  1265 => (x"4f",x"54",x"53",x"59"),
  1266 => (x"50",x"20",x"45",x"4e"),
  1267 => (x"52",x"47",x"4f",x"52"),
  1268 => (x"20",x"2c",x"4d",x"41"),
  1269 => (x"54",x"53",x"27",x"31"),
  1270 => (x"52",x"54",x"53",x"20"),
  1271 => (x"0a",x"47",x"4e",x"49"),
  1272 => (x"00",x"00",x"00",x"00"),
  1273 => (x"5f",x"72",x"74",x"53"),
  1274 => (x"6f",x"4c",x"5f",x"32"),
  1275 => (x"20",x"20",x"3a",x"63"),
  1276 => (x"20",x"20",x"20",x"20"),
  1277 => (x"20",x"20",x"20",x"20"),
  1278 => (x"0a",x"73",x"25",x"20"),
  1279 => (x"00",x"00",x"00",x"00"),
  1280 => (x"20",x"20",x"20",x"20"),
  1281 => (x"20",x"20",x"20",x"20"),
  1282 => (x"75",x"6f",x"68",x"73"),
  1283 => (x"62",x"20",x"64",x"6c"),
  1284 => (x"20",x"20",x"3a",x"65"),
  1285 => (x"52",x"48",x"44",x"20"),
  1286 => (x"4f",x"54",x"53",x"59"),
  1287 => (x"50",x"20",x"45",x"4e"),
  1288 => (x"52",x"47",x"4f",x"52"),
  1289 => (x"20",x"2c",x"4d",x"41"),
  1290 => (x"44",x"4e",x"27",x"32"),
  1291 => (x"52",x"54",x"53",x"20"),
  1292 => (x"0a",x"47",x"4e",x"49"),
  1293 => (x"00",x"00",x"00",x"00"),
  1294 => (x"00",x"00",x"00",x"0a"),
  1295 => (x"72",x"65",x"73",x"55"),
  1296 => (x"6d",x"69",x"74",x"20"),
  1297 => (x"25",x"20",x"3a",x"65"),
  1298 => (x"0e",x"00",x"0a",x"64"),
  1299 => (x"c8",x"0e",x"5b",x"5e"),
  1300 => (x"66",x"cc",x"4b",x"66"),
  1301 => (x"c2",x"79",x"73",x"49"),
  1302 => (x"87",x"c4",x"05",x"ab"),
  1303 => (x"87",x"c2",x"4a",x"c1"),
  1304 => (x"9a",x"72",x"4a",x"c0"),
  1305 => (x"c3",x"87",x"c2",x"05"),
  1306 => (x"02",x"ab",x"c0",x"79"),
  1307 => (x"ab",x"c1",x"87",x"d8"),
  1308 => (x"c2",x"87",x"d7",x"02"),
  1309 => (x"e5",x"c0",x"02",x"ab"),
  1310 => (x"02",x"ab",x"c3",x"87"),
  1311 => (x"c4",x"87",x"e5",x"c0"),
  1312 => (x"87",x"de",x"02",x"ab"),
  1313 => (x"79",x"c0",x"87",x"de"),
  1314 => (x"d9",x"c1",x"87",x"da"),
  1315 => (x"c1",x"48",x"bf",x"c0"),
  1316 => (x"06",x"a8",x"b7",x"e4"),
  1317 => (x"79",x"c0",x"87",x"c4"),
  1318 => (x"79",x"c3",x"87",x"ca"),
  1319 => (x"79",x"c1",x"87",x"c6"),
  1320 => (x"79",x"c2",x"87",x"c2"),
  1321 => (x"4f",x"26",x"4b",x"26"),
  1322 => (x"48",x"66",x"c4",x"1e"),
  1323 => (x"c4",x"05",x"a8",x"c2"),
  1324 => (x"c2",x"48",x"c1",x"87"),
  1325 => (x"26",x"48",x"c0",x"87"),
  1326 => (x"66",x"c4",x"1e",x"4f"),
  1327 => (x"c8",x"81",x"c2",x"49"),
  1328 => (x"80",x"71",x"48",x"66"),
  1329 => (x"78",x"08",x"66",x"cc"),
  1330 => (x"0e",x"4f",x"26",x"08"),
  1331 => (x"5d",x"5c",x"5b",x"5e"),
  1332 => (x"c0",x"86",x"f4",x"0e"),
  1333 => (x"c5",x"4c",x"66",x"e4"),
  1334 => (x"c4",x"48",x"74",x"84"),
  1335 => (x"a6",x"c8",x"90",x"b7"),
  1336 => (x"48",x"66",x"dc",x"58"),
  1337 => (x"c4",x"80",x"66",x"c4"),
  1338 => (x"48",x"6e",x"58",x"a6"),
  1339 => (x"78",x"66",x"e8",x"c0"),
  1340 => (x"80",x"c1",x"48",x"74"),
  1341 => (x"c8",x"58",x"a6",x"cc"),
  1342 => (x"b7",x"c4",x"49",x"66"),
  1343 => (x"81",x"66",x"dc",x"91"),
  1344 => (x"79",x"66",x"e8",x"c0"),
  1345 => (x"81",x"de",x"49",x"74"),
  1346 => (x"dc",x"91",x"b7",x"c4"),
  1347 => (x"79",x"74",x"81",x"66"),
  1348 => (x"ac",x"b7",x"66",x"c8"),
  1349 => (x"87",x"e3",x"c0",x"01"),
  1350 => (x"c8",x"c3",x"49",x"74"),
  1351 => (x"e0",x"c0",x"91",x"b7"),
  1352 => (x"4d",x"c4",x"81",x"66"),
  1353 => (x"66",x"c4",x"4a",x"71"),
  1354 => (x"4b",x"66",x"c8",x"82"),
  1355 => (x"83",x"c1",x"8b",x"74"),
  1356 => (x"82",x"75",x"7a",x"74"),
  1357 => (x"9b",x"73",x"8b",x"c1"),
  1358 => (x"74",x"87",x"f5",x"01"),
  1359 => (x"b7",x"c8",x"c3",x"4a"),
  1360 => (x"66",x"e0",x"c0",x"92"),
  1361 => (x"c1",x"49",x"74",x"82"),
  1362 => (x"91",x"b7",x"c4",x"89"),
  1363 => (x"48",x"69",x"81",x"72"),
  1364 => (x"79",x"70",x"80",x"c1"),
  1365 => (x"81",x"d4",x"49",x"74"),
  1366 => (x"91",x"b7",x"c8",x"c3"),
  1367 => (x"81",x"66",x"e0",x"c0"),
  1368 => (x"6e",x"81",x"66",x"c4"),
  1369 => (x"d9",x"c1",x"79",x"bf"),
  1370 => (x"78",x"c5",x"48",x"c0"),
  1371 => (x"4d",x"26",x"8e",x"f4"),
  1372 => (x"4b",x"26",x"4c",x"26"),
  1373 => (x"5e",x"0e",x"4f",x"26"),
  1374 => (x"c8",x"97",x"0e",x"5b"),
  1375 => (x"4a",x"73",x"4b",x"66"),
  1376 => (x"ba",x"82",x"c0",x"fe"),
  1377 => (x"49",x"66",x"cc",x"97"),
  1378 => (x"b9",x"81",x"c0",x"fe"),
  1379 => (x"02",x"aa",x"b7",x"71"),
  1380 => (x"48",x"c0",x"87",x"c4"),
  1381 => (x"d9",x"c1",x"87",x"c7"),
  1382 => (x"c1",x"5b",x"97",x"cc"),
  1383 => (x"26",x"4b",x"26",x"48"),
  1384 => (x"5b",x"5e",x"0e",x"4f"),
  1385 => (x"f8",x"0e",x"5d",x"5c"),
  1386 => (x"dc",x"4d",x"c2",x"86"),
  1387 => (x"81",x"c1",x"49",x"66"),
  1388 => (x"c2",x"4c",x"66",x"d8"),
  1389 => (x"c2",x"4b",x"71",x"84"),
  1390 => (x"fe",x"49",x"13",x"83"),
  1391 => (x"c3",x"b9",x"81",x"c0"),
  1392 => (x"4a",x"14",x"99",x"ff"),
  1393 => (x"ba",x"82",x"c0",x"fe"),
  1394 => (x"5a",x"97",x"a6",x"c4"),
  1395 => (x"fe",x"4a",x"6e",x"97"),
  1396 => (x"fe",x"ba",x"82",x"c0"),
  1397 => (x"71",x"b9",x"81",x"c0"),
  1398 => (x"c7",x"02",x"aa",x"b7"),
  1399 => (x"48",x"a6",x"c4",x"87"),
  1400 => (x"87",x"cc",x"78",x"c0"),
  1401 => (x"48",x"c8",x"d9",x"c1"),
  1402 => (x"c4",x"50",x"6e",x"97"),
  1403 => (x"78",x"c1",x"48",x"a6"),
  1404 => (x"c2",x"05",x"66",x"c4"),
  1405 => (x"c2",x"85",x"c1",x"87"),
  1406 => (x"fe",x"06",x"ad",x"b7"),
  1407 => (x"66",x"d8",x"87",x"fb"),
  1408 => (x"49",x"66",x"dc",x"4a"),
  1409 => (x"87",x"ee",x"f7",x"fe"),
  1410 => (x"06",x"a8",x"b7",x"c0"),
  1411 => (x"48",x"75",x"87",x"cc"),
  1412 => (x"d9",x"c1",x"80",x"c7"),
  1413 => (x"48",x"c1",x"58",x"c4"),
  1414 => (x"48",x"c0",x"87",x"c2"),
  1415 => (x"4d",x"26",x"8e",x"f8"),
  1416 => (x"4b",x"26",x"4c",x"26"),
  1417 => (x"4b",x"26",x"4f",x"26"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
