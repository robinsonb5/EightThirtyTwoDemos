
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"c9",x"01"),
     1 => (x"cf",x"03",x"87",x"cc"),
     2 => (x"87",x"fd",x"00",x"87"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"36",x"27",x"4f",x"00"),
     5 => (x"4f",x"00",x"00",x"00"),
     6 => (x"0e",x"1e",x"18",x"0e"),
     7 => (x"00",x"00",x"44",x"27"),
     8 => (x"48",x"26",x"0f",x"00"),
     9 => (x"08",x"26",x"80",x"ff"),
    10 => (x"c0",x"c0",x"c2",x"4f"),
    11 => (x"05",x"2d",x"27",x"4e"),
    12 => (x"00",x"0f",x"00",x"00"),
    13 => (x"f0",x"c1",x"87",x"fd"),
    14 => (x"43",x"27",x"4e",x"c0"),
    15 => (x"0f",x"00",x"00",x"00"),
    16 => (x"4f",x"87",x"fd",x"00"),
    17 => (x"0e",x"1e",x"18",x"0e"),
    18 => (x"80",x"ff",x"48",x"26"),
    19 => (x"1e",x"4f",x"08",x"26"),
    20 => (x"ff",x"1e",x"1e",x"72"),
    21 => (x"48",x"6a",x"4a",x"c0"),
    22 => (x"c4",x"98",x"c0",x"c4"),
    23 => (x"02",x"6e",x"58",x"a6"),
    24 => (x"cc",x"87",x"f3",x"ff"),
    25 => (x"66",x"cc",x"7a",x"66"),
    26 => (x"4a",x"26",x"26",x"48"),
    27 => (x"5e",x"0e",x"4f",x"26"),
    28 => (x"5d",x"5c",x"5b",x"5a"),
    29 => (x"4d",x"66",x"d4",x"0e"),
    30 => (x"4b",x"15",x"4c",x"c0"),
    31 => (x"c0",x"02",x"9b",x"73"),
    32 => (x"4a",x"73",x"87",x"d6"),
    33 => (x"4f",x"27",x"1e",x"72"),
    34 => (x"0f",x"00",x"00",x"00"),
    35 => (x"84",x"c1",x"86",x"c4"),
    36 => (x"9b",x"73",x"4b",x"15"),
    37 => (x"87",x"ea",x"ff",x"05"),
    38 => (x"4d",x"26",x"48",x"74"),
    39 => (x"4b",x"26",x"4c",x"26"),
    40 => (x"4f",x"26",x"4a",x"26"),
    41 => (x"5b",x"5a",x"5e",x"0e"),
    42 => (x"1e",x"0e",x"5d",x"5c"),
    43 => (x"27",x"4d",x"66",x"d8"),
    44 => (x"00",x"00",x"15",x"f0"),
    45 => (x"27",x"49",x"76",x"4b"),
    46 => (x"00",x"00",x"0e",x"30"),
    47 => (x"75",x"4c",x"c0",x"79"),
    48 => (x"a9",x"b7",x"c0",x"49"),
    49 => (x"87",x"ce",x"c0",x"03"),
    50 => (x"27",x"1e",x"ed",x"c0"),
    51 => (x"00",x"00",x"00",x"4f"),
    52 => (x"c0",x"86",x"c4",x"0f"),
    53 => (x"9d",x"75",x"8d",x"0d"),
    54 => (x"87",x"c6",x"c0",x"05"),
    55 => (x"c0",x"53",x"f0",x"c0"),
    56 => (x"9d",x"75",x"87",x"f6"),
    57 => (x"87",x"f0",x"c0",x"02"),
    58 => (x"1e",x"72",x"49",x"75"),
    59 => (x"4a",x"66",x"e4",x"c0"),
    60 => (x"00",x"04",x"c8",x"27"),
    61 => (x"4a",x"26",x"0f",x"00"),
    62 => (x"4a",x"72",x"4a",x"71"),
    63 => (x"53",x"12",x"82",x"6e"),
    64 => (x"1e",x"72",x"49",x"75"),
    65 => (x"4a",x"66",x"e4",x"c0"),
    66 => (x"00",x"04",x"c8",x"27"),
    67 => (x"4a",x"26",x"0f",x"00"),
    68 => (x"9d",x"75",x"4d",x"70"),
    69 => (x"87",x"d0",x"ff",x"05"),
    70 => (x"f0",x"27",x"49",x"73"),
    71 => (x"b7",x"00",x"00",x"15"),
    72 => (x"e1",x"c0",x"02",x"a9"),
    73 => (x"dc",x"8b",x"c1",x"87"),
    74 => (x"97",x"49",x"bf",x"a6"),
    75 => (x"66",x"dc",x"51",x"6b"),
    76 => (x"c0",x"80",x"c1",x"48"),
    77 => (x"c1",x"58",x"a6",x"e0"),
    78 => (x"27",x"49",x"73",x"84"),
    79 => (x"00",x"00",x"15",x"f0"),
    80 => (x"ff",x"05",x"a9",x"b7"),
    81 => (x"a6",x"dc",x"87",x"df"),
    82 => (x"51",x"c0",x"49",x"bf"),
    83 => (x"26",x"26",x"48",x"74"),
    84 => (x"26",x"4c",x"26",x"4d"),
    85 => (x"26",x"4a",x"26",x"4b"),
    86 => (x"5a",x"5e",x"0e",x"4f"),
    87 => (x"0e",x"5d",x"5c",x"5b"),
    88 => (x"76",x"4c",x"c0",x"1e"),
    89 => (x"dc",x"79",x"c0",x"49"),
    90 => (x"66",x"d8",x"4b",x"a6"),
    91 => (x"48",x"66",x"d8",x"4a"),
    92 => (x"a6",x"dc",x"80",x"c1"),
    93 => (x"d8",x"4d",x"12",x"58"),
    94 => (x"75",x"2d",x"b7",x"35"),
    95 => (x"d7",x"c4",x"02",x"9d"),
    96 => (x"c3",x"02",x"6e",x"87"),
    97 => (x"49",x"76",x"87",x"e1"),
    98 => (x"4a",x"75",x"79",x"c0"),
    99 => (x"e3",x"c1",x"49",x"75"),
   100 => (x"e5",x"c2",x"02",x"a9"),
   101 => (x"c1",x"49",x"72",x"87"),
   102 => (x"c0",x"02",x"a9",x"e4"),
   103 => (x"49",x"72",x"87",x"de"),
   104 => (x"02",x"a9",x"ec",x"c1"),
   105 => (x"72",x"87",x"cc",x"c2"),
   106 => (x"a9",x"f3",x"c1",x"49"),
   107 => (x"87",x"ea",x"c1",x"02"),
   108 => (x"f8",x"c1",x"49",x"72"),
   109 => (x"f2",x"c0",x"02",x"a9"),
   110 => (x"87",x"d3",x"c2",x"87"),
   111 => (x"40",x"27",x"1e",x"ca"),
   112 => (x"1e",x"00",x"00",x"16"),
   113 => (x"4a",x"73",x"83",x"c4"),
   114 => (x"1e",x"6a",x"8a",x"c4"),
   115 => (x"00",x"00",x"a4",x"27"),
   116 => (x"86",x"cc",x"0f",x"00"),
   117 => (x"4c",x"74",x"4a",x"70"),
   118 => (x"40",x"27",x"84",x"72"),
   119 => (x"1e",x"00",x"00",x"16"),
   120 => (x"00",x"00",x"6e",x"27"),
   121 => (x"86",x"c4",x"0f",x"00"),
   122 => (x"d0",x"87",x"d6",x"c2"),
   123 => (x"16",x"40",x"27",x"1e"),
   124 => (x"c4",x"1e",x"00",x"00"),
   125 => (x"c4",x"4a",x"73",x"83"),
   126 => (x"27",x"1e",x"6a",x"8a"),
   127 => (x"00",x"00",x"00",x"a4"),
   128 => (x"70",x"86",x"cc",x"0f"),
   129 => (x"72",x"4c",x"74",x"4a"),
   130 => (x"16",x"40",x"27",x"84"),
   131 => (x"27",x"1e",x"00",x"00"),
   132 => (x"00",x"00",x"00",x"6e"),
   133 => (x"c1",x"86",x"c4",x"0f"),
   134 => (x"83",x"c4",x"87",x"e7"),
   135 => (x"8a",x"c4",x"4a",x"73"),
   136 => (x"6e",x"27",x"1e",x"6a"),
   137 => (x"0f",x"00",x"00",x"00"),
   138 => (x"4a",x"70",x"86",x"c4"),
   139 => (x"84",x"72",x"4c",x"74"),
   140 => (x"76",x"87",x"ce",x"c1"),
   141 => (x"c1",x"79",x"c1",x"49"),
   142 => (x"83",x"c4",x"87",x"c7"),
   143 => (x"8a",x"c4",x"4a",x"73"),
   144 => (x"4f",x"27",x"1e",x"6a"),
   145 => (x"0f",x"00",x"00",x"00"),
   146 => (x"84",x"c1",x"86",x"c4"),
   147 => (x"c0",x"87",x"f2",x"c0"),
   148 => (x"4f",x"27",x"1e",x"e5"),
   149 => (x"0f",x"00",x"00",x"00"),
   150 => (x"1e",x"75",x"86",x"c4"),
   151 => (x"00",x"00",x"4f",x"27"),
   152 => (x"86",x"c4",x"0f",x"00"),
   153 => (x"75",x"87",x"da",x"c0"),
   154 => (x"a9",x"e5",x"c0",x"49"),
   155 => (x"87",x"c7",x"c0",x"05"),
   156 => (x"79",x"c1",x"49",x"76"),
   157 => (x"75",x"87",x"ca",x"c0"),
   158 => (x"00",x"4f",x"27",x"1e"),
   159 => (x"c4",x"0f",x"00",x"00"),
   160 => (x"4a",x"66",x"d8",x"86"),
   161 => (x"c1",x"48",x"66",x"d8"),
   162 => (x"58",x"a6",x"dc",x"80"),
   163 => (x"35",x"d8",x"4d",x"12"),
   164 => (x"9d",x"75",x"2d",x"b7"),
   165 => (x"87",x"e9",x"fb",x"05"),
   166 => (x"26",x"26",x"48",x"74"),
   167 => (x"26",x"4c",x"26",x"4d"),
   168 => (x"26",x"4a",x"26",x"4b"),
   169 => (x"5a",x"5e",x"0e",x"4f"),
   170 => (x"66",x"d0",x"0e",x"5b"),
   171 => (x"7b",x"66",x"cc",x"4b"),
   172 => (x"27",x"1e",x"66",x"cc"),
   173 => (x"00",x"00",x"04",x"b4"),
   174 => (x"70",x"86",x"c4",x"0f"),
   175 => (x"05",x"9a",x"72",x"4a"),
   176 => (x"c3",x"87",x"c2",x"c0"),
   177 => (x"4a",x"66",x"cc",x"7b"),
   178 => (x"c0",x"49",x"66",x"cc"),
   179 => (x"c0",x"02",x"a9",x"b7"),
   180 => (x"49",x"72",x"87",x"e7"),
   181 => (x"02",x"a9",x"b7",x"c1"),
   182 => (x"72",x"87",x"e3",x"c0"),
   183 => (x"a9",x"b7",x"c2",x"49"),
   184 => (x"87",x"f3",x"c0",x"02"),
   185 => (x"b7",x"c3",x"49",x"72"),
   186 => (x"f1",x"c0",x"02",x"a9"),
   187 => (x"c4",x"49",x"72",x"87"),
   188 => (x"c0",x"02",x"a9",x"b7"),
   189 => (x"e5",x"c0",x"87",x"e6"),
   190 => (x"c0",x"7b",x"c0",x"87"),
   191 => (x"ec",x"27",x"87",x"e0"),
   192 => (x"bf",x"00",x"00",x"17"),
   193 => (x"b7",x"e4",x"c1",x"49"),
   194 => (x"c5",x"c0",x"06",x"a9"),
   195 => (x"c0",x"7b",x"c0",x"87"),
   196 => (x"7b",x"c3",x"87",x"cc"),
   197 => (x"c1",x"87",x"c7",x"c0"),
   198 => (x"87",x"c2",x"c0",x"7b"),
   199 => (x"4b",x"26",x"7b",x"c2"),
   200 => (x"4f",x"26",x"4a",x"26"),
   201 => (x"c8",x"1e",x"72",x"1e"),
   202 => (x"82",x"c2",x"4a",x"66"),
   203 => (x"72",x"48",x"66",x"cc"),
   204 => (x"49",x"66",x"d0",x"80"),
   205 => (x"4a",x"26",x"79",x"70"),
   206 => (x"5e",x"0e",x"4f",x"26"),
   207 => (x"5d",x"5c",x"5b",x"5a"),
   208 => (x"4d",x"66",x"dc",x"0e"),
   209 => (x"4a",x"75",x"85",x"c5"),
   210 => (x"4a",x"72",x"92",x"c4"),
   211 => (x"c0",x"82",x"66",x"d4"),
   212 => (x"72",x"7a",x"66",x"e0"),
   213 => (x"6a",x"83",x"c4",x"4b"),
   214 => (x"82",x"f8",x"c1",x"7b"),
   215 => (x"4c",x"75",x"7a",x"75"),
   216 => (x"82",x"c1",x"4a",x"75"),
   217 => (x"b7",x"72",x"49",x"75"),
   218 => (x"e3",x"c0",x"01",x"a9"),
   219 => (x"c3",x"4b",x"75",x"87"),
   220 => (x"4b",x"73",x"93",x"c8"),
   221 => (x"74",x"83",x"66",x"d8"),
   222 => (x"72",x"92",x"c4",x"4a"),
   223 => (x"75",x"82",x"73",x"4a"),
   224 => (x"75",x"84",x"c1",x"7a"),
   225 => (x"74",x"82",x"c1",x"4a"),
   226 => (x"a9",x"b7",x"72",x"49"),
   227 => (x"87",x"dd",x"ff",x"06"),
   228 => (x"c8",x"c3",x"4c",x"75"),
   229 => (x"d8",x"4c",x"74",x"94"),
   230 => (x"4a",x"75",x"84",x"66"),
   231 => (x"4b",x"74",x"92",x"c4"),
   232 => (x"8b",x"c4",x"83",x"72"),
   233 => (x"80",x"c1",x"48",x"6b"),
   234 => (x"66",x"d4",x"7b",x"70"),
   235 => (x"c0",x"83",x"72",x"4b"),
   236 => (x"72",x"84",x"e0",x"fe"),
   237 => (x"6b",x"82",x"74",x"4a"),
   238 => (x"17",x"ec",x"27",x"7a"),
   239 => (x"c5",x"49",x"00",x"00"),
   240 => (x"26",x"4d",x"26",x"79"),
   241 => (x"26",x"4b",x"26",x"4c"),
   242 => (x"0e",x"4f",x"26",x"4a"),
   243 => (x"5c",x"5b",x"5a",x"5e"),
   244 => (x"66",x"d0",x"97",x"0e"),
   245 => (x"d8",x"4b",x"74",x"4c"),
   246 => (x"97",x"2b",x"b7",x"33"),
   247 => (x"d8",x"4a",x"66",x"d4"),
   248 => (x"73",x"2a",x"b7",x"32"),
   249 => (x"a9",x"b7",x"72",x"49"),
   250 => (x"87",x"c5",x"c0",x"02"),
   251 => (x"ca",x"c0",x"48",x"c0"),
   252 => (x"16",x"e0",x"27",x"87"),
   253 => (x"74",x"49",x"00",x"00"),
   254 => (x"26",x"48",x"c1",x"51"),
   255 => (x"26",x"4b",x"26",x"4c"),
   256 => (x"0e",x"4f",x"26",x"4a"),
   257 => (x"0e",x"5b",x"5a",x"5e"),
   258 => (x"d4",x"4b",x"c2",x"1e"),
   259 => (x"82",x"c1",x"4a",x"66"),
   260 => (x"6a",x"97",x"82",x"73"),
   261 => (x"b7",x"32",x"d8",x"4a"),
   262 => (x"d4",x"1e",x"72",x"2a"),
   263 => (x"82",x"73",x"4a",x"66"),
   264 => (x"d8",x"4a",x"6a",x"97"),
   265 => (x"72",x"2a",x"b7",x"32"),
   266 => (x"03",x"cb",x"27",x"1e"),
   267 => (x"c8",x"0f",x"00",x"00"),
   268 => (x"72",x"4a",x"70",x"86"),
   269 => (x"c7",x"c0",x"05",x"9a"),
   270 => (x"c1",x"49",x"76",x"87"),
   271 => (x"83",x"c1",x"51",x"c1"),
   272 => (x"b7",x"c2",x"49",x"73"),
   273 => (x"c2",x"ff",x"06",x"a9"),
   274 => (x"4a",x"6e",x"97",x"87"),
   275 => (x"2a",x"b7",x"32",x"d8"),
   276 => (x"d7",x"c1",x"49",x"72"),
   277 => (x"c0",x"04",x"a9",x"b7"),
   278 => (x"6e",x"97",x"87",x"d3"),
   279 => (x"b7",x"32",x"d8",x"4a"),
   280 => (x"c1",x"49",x"72",x"2a"),
   281 => (x"03",x"a9",x"b7",x"da"),
   282 => (x"c7",x"87",x"c2",x"c0"),
   283 => (x"4a",x"6e",x"97",x"4b"),
   284 => (x"2a",x"b7",x"32",x"d8"),
   285 => (x"d2",x"c1",x"49",x"72"),
   286 => (x"c0",x"05",x"a9",x"b7"),
   287 => (x"48",x"c1",x"87",x"c5"),
   288 => (x"d4",x"87",x"ea",x"c0"),
   289 => (x"66",x"d4",x"1e",x"66"),
   290 => (x"05",x"12",x"27",x"1e"),
   291 => (x"c8",x"0f",x"00",x"00"),
   292 => (x"72",x"4a",x"70",x"86"),
   293 => (x"a9",x"b7",x"c0",x"49"),
   294 => (x"87",x"cf",x"c0",x"06"),
   295 => (x"80",x"c7",x"48",x"73"),
   296 => (x"00",x"17",x"f0",x"27"),
   297 => (x"48",x"c1",x"58",x"00"),
   298 => (x"c0",x"87",x"c2",x"c0"),
   299 => (x"4b",x"26",x"26",x"48"),
   300 => (x"4f",x"26",x"4a",x"26"),
   301 => (x"49",x"66",x"c4",x"1e"),
   302 => (x"05",x"a9",x"b7",x"c2"),
   303 => (x"c1",x"87",x"c5",x"c0"),
   304 => (x"87",x"c2",x"c0",x"48"),
   305 => (x"4f",x"26",x"48",x"c0"),
   306 => (x"72",x"1e",x"73",x"1e"),
   307 => (x"87",x"d9",x"02",x"9a"),
   308 => (x"4b",x"c1",x"48",x"c0"),
   309 => (x"82",x"01",x"a9",x"72"),
   310 => (x"87",x"f8",x"83",x"73"),
   311 => (x"89",x"03",x"a9",x"72"),
   312 => (x"c1",x"07",x"80",x"73"),
   313 => (x"f3",x"05",x"2b",x"2a"),
   314 => (x"26",x"4b",x"26",x"87"),
   315 => (x"1e",x"75",x"1e",x"4f"),
   316 => (x"a1",x"71",x"4d",x"c0"),
   317 => (x"c1",x"b9",x"ff",x"04"),
   318 => (x"72",x"07",x"bd",x"81"),
   319 => (x"ba",x"ff",x"04",x"a2"),
   320 => (x"07",x"bd",x"82",x"c1"),
   321 => (x"9d",x"75",x"87",x"c2"),
   322 => (x"c1",x"b8",x"ff",x"05"),
   323 => (x"4d",x"25",x"07",x"80"),
   324 => (x"c4",x"1e",x"4f",x"26"),
   325 => (x"66",x"c8",x"4a",x"66"),
   326 => (x"11",x"48",x"12",x"49"),
   327 => (x"88",x"87",x"c4",x"02"),
   328 => (x"26",x"87",x"f6",x"02"),
   329 => (x"c8",x"ff",x"1e",x"4f"),
   330 => (x"26",x"48",x"68",x"48"),
   331 => (x"5a",x"5e",x"0e",x"4f"),
   332 => (x"0e",x"5d",x"5c",x"5b"),
   333 => (x"66",x"c4",x"8e",x"d0"),
   334 => (x"16",x"e8",x"27",x"4c"),
   335 => (x"27",x"49",x"00",x"00"),
   336 => (x"00",x"00",x"16",x"f0"),
   337 => (x"16",x"68",x"27",x"79"),
   338 => (x"27",x"49",x"00",x"00"),
   339 => (x"00",x"00",x"16",x"b0"),
   340 => (x"16",x"b0",x"27",x"79"),
   341 => (x"27",x"49",x"00",x"00"),
   342 => (x"00",x"00",x"16",x"f0"),
   343 => (x"16",x"b4",x"27",x"79"),
   344 => (x"c0",x"49",x"00",x"00"),
   345 => (x"16",x"b8",x"27",x"79"),
   346 => (x"c2",x"49",x"00",x"00"),
   347 => (x"16",x"bc",x"27",x"79"),
   348 => (x"c0",x"49",x"00",x"00"),
   349 => (x"c0",x"27",x"79",x"e8"),
   350 => (x"49",x"00",x"00",x"16"),
   351 => (x"00",x"0f",x"ba",x"27"),
   352 => (x"1e",x"72",x"48",x"00"),
   353 => (x"10",x"4a",x"a1",x"df"),
   354 => (x"05",x"aa",x"71",x"51"),
   355 => (x"4a",x"26",x"87",x"f9"),
   356 => (x"00",x"16",x"70",x"27"),
   357 => (x"d9",x"27",x"49",x"00"),
   358 => (x"48",x"00",x"00",x"0f"),
   359 => (x"a1",x"df",x"1e",x"72"),
   360 => (x"71",x"51",x"10",x"4a"),
   361 => (x"87",x"f9",x"05",x"aa"),
   362 => (x"5c",x"27",x"4a",x"26"),
   363 => (x"49",x"00",x"00",x"1e"),
   364 => (x"f8",x"27",x"79",x"ca"),
   365 => (x"1e",x"00",x"00",x"0f"),
   366 => (x"00",x"01",x"59",x"27"),
   367 => (x"86",x"c4",x"0f",x"00"),
   368 => (x"00",x"0f",x"fa",x"27"),
   369 => (x"59",x"27",x"1e",x"00"),
   370 => (x"0f",x"00",x"00",x"01"),
   371 => (x"2a",x"27",x"86",x"c4"),
   372 => (x"1e",x"00",x"00",x"10"),
   373 => (x"00",x"01",x"59",x"27"),
   374 => (x"86",x"c4",x"0f",x"00"),
   375 => (x"00",x"15",x"de",x"27"),
   376 => (x"c0",x"02",x"bf",x"00"),
   377 => (x"41",x"27",x"87",x"df"),
   378 => (x"1e",x"00",x"00",x"0e"),
   379 => (x"00",x"01",x"59",x"27"),
   380 => (x"86",x"c4",x"0f",x"00"),
   381 => (x"00",x"0e",x"6d",x"27"),
   382 => (x"59",x"27",x"1e",x"00"),
   383 => (x"0f",x"00",x"00",x"01"),
   384 => (x"dc",x"c0",x"86",x"c4"),
   385 => (x"0e",x"6f",x"27",x"87"),
   386 => (x"27",x"1e",x"00",x"00"),
   387 => (x"00",x"00",x"01",x"59"),
   388 => (x"27",x"86",x"c4",x"0f"),
   389 => (x"00",x"00",x"0e",x"9e"),
   390 => (x"01",x"59",x"27",x"1e"),
   391 => (x"c4",x"0f",x"00",x"00"),
   392 => (x"15",x"e2",x"27",x"86"),
   393 => (x"1e",x"bf",x"00",x"00"),
   394 => (x"00",x"10",x"2c",x"27"),
   395 => (x"59",x"27",x"1e",x"00"),
   396 => (x"0f",x"00",x"00",x"01"),
   397 => (x"25",x"27",x"86",x"c8"),
   398 => (x"0f",x"00",x"00",x"05"),
   399 => (x"00",x"16",x"68",x"27"),
   400 => (x"4d",x"c1",x"58",x"00"),
   401 => (x"00",x"15",x"e2",x"27"),
   402 => (x"c0",x"49",x"bf",x"00"),
   403 => (x"c6",x"06",x"a9",x"b7"),
   404 => (x"1c",x"27",x"87",x"cf"),
   405 => (x"0f",x"00",x"00",x"0e"),
   406 => (x"00",x"0d",x"e0",x"27"),
   407 => (x"49",x"76",x"0f",x"00"),
   408 => (x"4c",x"c3",x"79",x"c2"),
   409 => (x"00",x"16",x"90",x"27"),
   410 => (x"bf",x"27",x"49",x"00"),
   411 => (x"48",x"00",x"00",x"0e"),
   412 => (x"a1",x"df",x"1e",x"72"),
   413 => (x"71",x"51",x"10",x"4a"),
   414 => (x"87",x"f9",x"05",x"aa"),
   415 => (x"a6",x"c8",x"4a",x"26"),
   416 => (x"27",x"79",x"c1",x"49"),
   417 => (x"00",x"00",x"16",x"90"),
   418 => (x"16",x"70",x"27",x"1e"),
   419 => (x"27",x"1e",x"00",x"00"),
   420 => (x"00",x"00",x"04",x"03"),
   421 => (x"70",x"86",x"c8",x"0f"),
   422 => (x"05",x"9a",x"72",x"4a"),
   423 => (x"c1",x"87",x"c5",x"c0"),
   424 => (x"87",x"c2",x"c0",x"4a"),
   425 => (x"f0",x"27",x"4a",x"c0"),
   426 => (x"49",x"00",x"00",x"17"),
   427 => (x"49",x"6e",x"79",x"72"),
   428 => (x"03",x"a9",x"b7",x"74"),
   429 => (x"6e",x"87",x"ed",x"c0"),
   430 => (x"72",x"92",x"c5",x"4a"),
   431 => (x"d0",x"88",x"74",x"48"),
   432 => (x"a6",x"cc",x"58",x"a6"),
   433 => (x"74",x"1e",x"72",x"4a"),
   434 => (x"1e",x"66",x"c8",x"1e"),
   435 => (x"00",x"03",x"24",x"27"),
   436 => (x"86",x"cc",x"0f",x"00"),
   437 => (x"80",x"c1",x"48",x"6e"),
   438 => (x"6e",x"58",x"a6",x"c4"),
   439 => (x"a9",x"b7",x"74",x"49"),
   440 => (x"87",x"d3",x"ff",x"04"),
   441 => (x"c4",x"1e",x"66",x"cc"),
   442 => (x"00",x"27",x"1e",x"66"),
   443 => (x"1e",x"00",x"00",x"18"),
   444 => (x"00",x"17",x"20",x"27"),
   445 => (x"3a",x"27",x"1e",x"00"),
   446 => (x"0f",x"00",x"00",x"03"),
   447 => (x"68",x"27",x"86",x"d0"),
   448 => (x"bf",x"00",x"00",x"16"),
   449 => (x"0c",x"c5",x"27",x"1e"),
   450 => (x"c4",x"0f",x"00",x"00"),
   451 => (x"49",x"a6",x"c4",x"86"),
   452 => (x"27",x"51",x"c1",x"c1"),
   453 => (x"00",x"00",x"17",x"e8"),
   454 => (x"d8",x"4a",x"bf",x"97"),
   455 => (x"72",x"2a",x"b7",x"32"),
   456 => (x"b7",x"c1",x"c1",x"49"),
   457 => (x"fb",x"c1",x"04",x"a9"),
   458 => (x"1e",x"c3",x"c1",x"87"),
   459 => (x"4a",x"66",x"c8",x"97"),
   460 => (x"2a",x"b7",x"32",x"d8"),
   461 => (x"cb",x"27",x"1e",x"72"),
   462 => (x"0f",x"00",x"00",x"03"),
   463 => (x"4a",x"70",x"86",x"c8"),
   464 => (x"72",x"49",x"66",x"c8"),
   465 => (x"c0",x"05",x"a9",x"b7"),
   466 => (x"a6",x"c8",x"87",x"f3"),
   467 => (x"c0",x"1e",x"72",x"4a"),
   468 => (x"02",x"a5",x"27",x"1e"),
   469 => (x"c8",x"0f",x"00",x"00"),
   470 => (x"16",x"90",x"27",x"86"),
   471 => (x"27",x"49",x"00",x"00"),
   472 => (x"00",x"00",x"0e",x"a0"),
   473 => (x"df",x"1e",x"72",x"48"),
   474 => (x"51",x"10",x"4a",x"a1"),
   475 => (x"f9",x"05",x"aa",x"71"),
   476 => (x"75",x"4a",x"26",x"87"),
   477 => (x"17",x"ec",x"27",x"4c"),
   478 => (x"75",x"49",x"00",x"00"),
   479 => (x"66",x"c4",x"97",x"79"),
   480 => (x"c4",x"80",x"c1",x"48"),
   481 => (x"97",x"50",x"08",x"a6"),
   482 => (x"d8",x"4b",x"66",x"c4"),
   483 => (x"27",x"2b",x"b7",x"33"),
   484 => (x"00",x"00",x"17",x"e8"),
   485 => (x"d8",x"4a",x"bf",x"97"),
   486 => (x"73",x"2a",x"b7",x"32"),
   487 => (x"a9",x"b7",x"72",x"49"),
   488 => (x"87",x"c5",x"fe",x"06"),
   489 => (x"49",x"74",x"94",x"6e"),
   490 => (x"66",x"d0",x"1e",x"72"),
   491 => (x"04",x"c8",x"27",x"4a"),
   492 => (x"26",x"0f",x"00",x"00"),
   493 => (x"c4",x"48",x"70",x"4a"),
   494 => (x"4a",x"74",x"58",x"a6"),
   495 => (x"c7",x"8a",x"66",x"cc"),
   496 => (x"6e",x"4c",x"72",x"92"),
   497 => (x"72",x"4a",x"76",x"8c"),
   498 => (x"0d",x"64",x"27",x"1e"),
   499 => (x"c4",x"0f",x"00",x"00"),
   500 => (x"75",x"85",x"c1",x"86"),
   501 => (x"15",x"e2",x"27",x"49"),
   502 => (x"b7",x"bf",x"00",x"00"),
   503 => (x"f1",x"f9",x"06",x"a9"),
   504 => (x"05",x"25",x"27",x"87"),
   505 => (x"27",x"0f",x"00",x"00"),
   506 => (x"00",x"00",x"16",x"e8"),
   507 => (x"10",x"59",x"27",x"58"),
   508 => (x"27",x"1e",x"00",x"00"),
   509 => (x"00",x"00",x"01",x"59"),
   510 => (x"27",x"86",x"c4",x"0f"),
   511 => (x"00",x"00",x"10",x"69"),
   512 => (x"01",x"59",x"27",x"1e"),
   513 => (x"c4",x"0f",x"00",x"00"),
   514 => (x"10",x"6b",x"27",x"86"),
   515 => (x"27",x"1e",x"00",x"00"),
   516 => (x"00",x"00",x"01",x"59"),
   517 => (x"27",x"86",x"c4",x"0f"),
   518 => (x"00",x"00",x"10",x"a1"),
   519 => (x"01",x"59",x"27",x"1e"),
   520 => (x"c4",x"0f",x"00",x"00"),
   521 => (x"17",x"ec",x"27",x"86"),
   522 => (x"1e",x"bf",x"00",x"00"),
   523 => (x"00",x"10",x"a3",x"27"),
   524 => (x"59",x"27",x"1e",x"00"),
   525 => (x"0f",x"00",x"00",x"01"),
   526 => (x"1e",x"c5",x"86",x"c8"),
   527 => (x"00",x"10",x"bc",x"27"),
   528 => (x"59",x"27",x"1e",x"00"),
   529 => (x"0f",x"00",x"00",x"01"),
   530 => (x"f0",x"27",x"86",x"c8"),
   531 => (x"bf",x"00",x"00",x"17"),
   532 => (x"10",x"d5",x"27",x"1e"),
   533 => (x"27",x"1e",x"00",x"00"),
   534 => (x"00",x"00",x"01",x"59"),
   535 => (x"c1",x"86",x"c8",x"0f"),
   536 => (x"10",x"ee",x"27",x"1e"),
   537 => (x"27",x"1e",x"00",x"00"),
   538 => (x"00",x"00",x"01",x"59"),
   539 => (x"27",x"86",x"c8",x"0f"),
   540 => (x"00",x"00",x"16",x"e0"),
   541 => (x"d8",x"4a",x"bf",x"97"),
   542 => (x"72",x"2a",x"b7",x"32"),
   543 => (x"11",x"07",x"27",x"1e"),
   544 => (x"27",x"1e",x"00",x"00"),
   545 => (x"00",x"00",x"01",x"59"),
   546 => (x"c1",x"86",x"c8",x"0f"),
   547 => (x"20",x"27",x"1e",x"c1"),
   548 => (x"1e",x"00",x"00",x"11"),
   549 => (x"00",x"01",x"59",x"27"),
   550 => (x"86",x"c8",x"0f",x"00"),
   551 => (x"00",x"17",x"e8",x"27"),
   552 => (x"4a",x"bf",x"97",x"00"),
   553 => (x"2a",x"b7",x"32",x"d8"),
   554 => (x"39",x"27",x"1e",x"72"),
   555 => (x"1e",x"00",x"00",x"11"),
   556 => (x"00",x"01",x"59",x"27"),
   557 => (x"86",x"c8",x"0f",x"00"),
   558 => (x"27",x"1e",x"c2",x"c1"),
   559 => (x"00",x"00",x"11",x"52"),
   560 => (x"01",x"59",x"27",x"1e"),
   561 => (x"c8",x"0f",x"00",x"00"),
   562 => (x"17",x"40",x"27",x"86"),
   563 => (x"1e",x"bf",x"00",x"00"),
   564 => (x"00",x"11",x"6b",x"27"),
   565 => (x"59",x"27",x"1e",x"00"),
   566 => (x"0f",x"00",x"00",x"01"),
   567 => (x"1e",x"c7",x"86",x"c8"),
   568 => (x"00",x"11",x"84",x"27"),
   569 => (x"59",x"27",x"1e",x"00"),
   570 => (x"0f",x"00",x"00",x"01"),
   571 => (x"5c",x"27",x"86",x"c8"),
   572 => (x"bf",x"00",x"00",x"1e"),
   573 => (x"11",x"9d",x"27",x"1e"),
   574 => (x"27",x"1e",x"00",x"00"),
   575 => (x"00",x"00",x"01",x"59"),
   576 => (x"27",x"86",x"c8",x"0f"),
   577 => (x"00",x"00",x"11",x"b6"),
   578 => (x"01",x"59",x"27",x"1e"),
   579 => (x"c4",x"0f",x"00",x"00"),
   580 => (x"11",x"e0",x"27",x"86"),
   581 => (x"27",x"1e",x"00",x"00"),
   582 => (x"00",x"00",x"01",x"59"),
   583 => (x"27",x"86",x"c4",x"0f"),
   584 => (x"00",x"00",x"16",x"68"),
   585 => (x"27",x"1e",x"bf",x"bf"),
   586 => (x"00",x"00",x"11",x"ec"),
   587 => (x"01",x"59",x"27",x"1e"),
   588 => (x"c8",x"0f",x"00",x"00"),
   589 => (x"12",x"05",x"27",x"86"),
   590 => (x"27",x"1e",x"00",x"00"),
   591 => (x"00",x"00",x"01",x"59"),
   592 => (x"27",x"86",x"c4",x"0f"),
   593 => (x"00",x"00",x"16",x"68"),
   594 => (x"82",x"c4",x"4a",x"bf"),
   595 => (x"36",x"27",x"1e",x"6a"),
   596 => (x"1e",x"00",x"00",x"12"),
   597 => (x"00",x"01",x"59",x"27"),
   598 => (x"86",x"c8",x"0f",x"00"),
   599 => (x"4f",x"27",x"1e",x"c0"),
   600 => (x"1e",x"00",x"00",x"12"),
   601 => (x"00",x"01",x"59",x"27"),
   602 => (x"86",x"c8",x"0f",x"00"),
   603 => (x"00",x"16",x"68",x"27"),
   604 => (x"c8",x"4a",x"bf",x"00"),
   605 => (x"27",x"1e",x"6a",x"82"),
   606 => (x"00",x"00",x"12",x"68"),
   607 => (x"01",x"59",x"27",x"1e"),
   608 => (x"c8",x"0f",x"00",x"00"),
   609 => (x"27",x"1e",x"c2",x"86"),
   610 => (x"00",x"00",x"12",x"81"),
   611 => (x"01",x"59",x"27",x"1e"),
   612 => (x"c8",x"0f",x"00",x"00"),
   613 => (x"16",x"68",x"27",x"86"),
   614 => (x"4a",x"bf",x"00",x"00"),
   615 => (x"1e",x"6a",x"82",x"cc"),
   616 => (x"00",x"12",x"9a",x"27"),
   617 => (x"59",x"27",x"1e",x"00"),
   618 => (x"0f",x"00",x"00",x"01"),
   619 => (x"1e",x"d1",x"86",x"c8"),
   620 => (x"00",x"12",x"b3",x"27"),
   621 => (x"59",x"27",x"1e",x"00"),
   622 => (x"0f",x"00",x"00",x"01"),
   623 => (x"68",x"27",x"86",x"c8"),
   624 => (x"bf",x"00",x"00",x"16"),
   625 => (x"72",x"82",x"d0",x"4a"),
   626 => (x"12",x"cc",x"27",x"1e"),
   627 => (x"27",x"1e",x"00",x"00"),
   628 => (x"00",x"00",x"01",x"59"),
   629 => (x"27",x"86",x"c8",x"0f"),
   630 => (x"00",x"00",x"12",x"e5"),
   631 => (x"01",x"59",x"27",x"1e"),
   632 => (x"c4",x"0f",x"00",x"00"),
   633 => (x"13",x"1a",x"27",x"86"),
   634 => (x"27",x"1e",x"00",x"00"),
   635 => (x"00",x"00",x"01",x"59"),
   636 => (x"27",x"86",x"c4",x"0f"),
   637 => (x"00",x"00",x"16",x"e8"),
   638 => (x"27",x"1e",x"bf",x"bf"),
   639 => (x"00",x"00",x"13",x"2b"),
   640 => (x"01",x"59",x"27",x"1e"),
   641 => (x"c8",x"0f",x"00",x"00"),
   642 => (x"13",x"44",x"27",x"86"),
   643 => (x"27",x"1e",x"00",x"00"),
   644 => (x"00",x"00",x"01",x"59"),
   645 => (x"27",x"86",x"c4",x"0f"),
   646 => (x"00",x"00",x"16",x"e8"),
   647 => (x"82",x"c4",x"4a",x"bf"),
   648 => (x"84",x"27",x"1e",x"6a"),
   649 => (x"1e",x"00",x"00",x"13"),
   650 => (x"00",x"01",x"59",x"27"),
   651 => (x"86",x"c8",x"0f",x"00"),
   652 => (x"9d",x"27",x"1e",x"c0"),
   653 => (x"1e",x"00",x"00",x"13"),
   654 => (x"00",x"01",x"59",x"27"),
   655 => (x"86",x"c8",x"0f",x"00"),
   656 => (x"00",x"16",x"e8",x"27"),
   657 => (x"c8",x"4a",x"bf",x"00"),
   658 => (x"27",x"1e",x"6a",x"82"),
   659 => (x"00",x"00",x"13",x"b6"),
   660 => (x"01",x"59",x"27",x"1e"),
   661 => (x"c8",x"0f",x"00",x"00"),
   662 => (x"27",x"1e",x"c1",x"86"),
   663 => (x"00",x"00",x"13",x"cf"),
   664 => (x"01",x"59",x"27",x"1e"),
   665 => (x"c8",x"0f",x"00",x"00"),
   666 => (x"16",x"e8",x"27",x"86"),
   667 => (x"4a",x"bf",x"00",x"00"),
   668 => (x"1e",x"6a",x"82",x"cc"),
   669 => (x"00",x"13",x"e8",x"27"),
   670 => (x"59",x"27",x"1e",x"00"),
   671 => (x"0f",x"00",x"00",x"01"),
   672 => (x"1e",x"d2",x"86",x"c8"),
   673 => (x"00",x"14",x"01",x"27"),
   674 => (x"59",x"27",x"1e",x"00"),
   675 => (x"0f",x"00",x"00",x"01"),
   676 => (x"e8",x"27",x"86",x"c8"),
   677 => (x"bf",x"00",x"00",x"16"),
   678 => (x"72",x"82",x"d0",x"4a"),
   679 => (x"14",x"1a",x"27",x"1e"),
   680 => (x"27",x"1e",x"00",x"00"),
   681 => (x"00",x"00",x"01",x"59"),
   682 => (x"27",x"86",x"c8",x"0f"),
   683 => (x"00",x"00",x"14",x"33"),
   684 => (x"01",x"59",x"27",x"1e"),
   685 => (x"c4",x"0f",x"00",x"00"),
   686 => (x"27",x"1e",x"6e",x"86"),
   687 => (x"00",x"00",x"14",x"68"),
   688 => (x"01",x"59",x"27",x"1e"),
   689 => (x"c8",x"0f",x"00",x"00"),
   690 => (x"27",x"1e",x"c5",x"86"),
   691 => (x"00",x"00",x"14",x"81"),
   692 => (x"01",x"59",x"27",x"1e"),
   693 => (x"c8",x"0f",x"00",x"00"),
   694 => (x"27",x"1e",x"74",x"86"),
   695 => (x"00",x"00",x"14",x"9a"),
   696 => (x"01",x"59",x"27",x"1e"),
   697 => (x"c8",x"0f",x"00",x"00"),
   698 => (x"27",x"1e",x"cd",x"86"),
   699 => (x"00",x"00",x"14",x"b3"),
   700 => (x"01",x"59",x"27",x"1e"),
   701 => (x"c8",x"0f",x"00",x"00"),
   702 => (x"1e",x"66",x"cc",x"86"),
   703 => (x"00",x"14",x"cc",x"27"),
   704 => (x"59",x"27",x"1e",x"00"),
   705 => (x"0f",x"00",x"00",x"01"),
   706 => (x"1e",x"c7",x"86",x"c8"),
   707 => (x"00",x"14",x"e5",x"27"),
   708 => (x"59",x"27",x"1e",x"00"),
   709 => (x"0f",x"00",x"00",x"01"),
   710 => (x"66",x"c8",x"86",x"c8"),
   711 => (x"14",x"fe",x"27",x"1e"),
   712 => (x"27",x"1e",x"00",x"00"),
   713 => (x"00",x"00",x"01",x"59"),
   714 => (x"c1",x"86",x"c8",x"0f"),
   715 => (x"15",x"17",x"27",x"1e"),
   716 => (x"27",x"1e",x"00",x"00"),
   717 => (x"00",x"00",x"01",x"59"),
   718 => (x"27",x"86",x"c8",x"0f"),
   719 => (x"00",x"00",x"16",x"70"),
   720 => (x"15",x"30",x"27",x"1e"),
   721 => (x"27",x"1e",x"00",x"00"),
   722 => (x"00",x"00",x"01",x"59"),
   723 => (x"27",x"86",x"c8",x"0f"),
   724 => (x"00",x"00",x"15",x"49"),
   725 => (x"01",x"59",x"27",x"1e"),
   726 => (x"c4",x"0f",x"00",x"00"),
   727 => (x"16",x"90",x"27",x"86"),
   728 => (x"27",x"1e",x"00",x"00"),
   729 => (x"00",x"00",x"15",x"7e"),
   730 => (x"01",x"59",x"27",x"1e"),
   731 => (x"c8",x"0f",x"00",x"00"),
   732 => (x"15",x"97",x"27",x"86"),
   733 => (x"27",x"1e",x"00",x"00"),
   734 => (x"00",x"00",x"01",x"59"),
   735 => (x"27",x"86",x"c4",x"0f"),
   736 => (x"00",x"00",x"15",x"cc"),
   737 => (x"01",x"59",x"27",x"1e"),
   738 => (x"c4",x"0f",x"00",x"00"),
   739 => (x"16",x"e4",x"27",x"86"),
   740 => (x"4a",x"bf",x"00",x"00"),
   741 => (x"00",x"16",x"64",x"27"),
   742 => (x"27",x"8a",x"bf",x"00"),
   743 => (x"00",x"00",x"16",x"6c"),
   744 => (x"72",x"79",x"72",x"49"),
   745 => (x"15",x"ce",x"27",x"1e"),
   746 => (x"27",x"1e",x"00",x"00"),
   747 => (x"00",x"00",x"01",x"59"),
   748 => (x"27",x"86",x"c8",x"0f"),
   749 => (x"00",x"00",x"16",x"6c"),
   750 => (x"f8",x"c1",x"49",x"bf"),
   751 => (x"c0",x"03",x"a9",x"b7"),
   752 => (x"de",x"27",x"87",x"ea"),
   753 => (x"1e",x"00",x"00",x"0e"),
   754 => (x"00",x"01",x"59",x"27"),
   755 => (x"86",x"c4",x"0f",x"00"),
   756 => (x"00",x"0f",x"14",x"27"),
   757 => (x"59",x"27",x"1e",x"00"),
   758 => (x"0f",x"00",x"00",x"01"),
   759 => (x"34",x"27",x"86",x"c4"),
   760 => (x"1e",x"00",x"00",x"0f"),
   761 => (x"00",x"01",x"59",x"27"),
   762 => (x"86",x"c4",x"0f",x"00"),
   763 => (x"00",x"16",x"6c",x"27"),
   764 => (x"72",x"4a",x"bf",x"00"),
   765 => (x"93",x"e8",x"cf",x"4b"),
   766 => (x"1e",x"72",x"49",x"73"),
   767 => (x"00",x"15",x"e2",x"27"),
   768 => (x"27",x"4a",x"bf",x"00"),
   769 => (x"00",x"00",x"04",x"c8"),
   770 => (x"70",x"4a",x"26",x"0f"),
   771 => (x"16",x"f0",x"27",x"48"),
   772 => (x"27",x"58",x"00",x"00"),
   773 => (x"00",x"00",x"15",x"e2"),
   774 => (x"4c",x"73",x"4b",x"bf"),
   775 => (x"74",x"94",x"e8",x"cf"),
   776 => (x"72",x"1e",x"72",x"49"),
   777 => (x"04",x"c8",x"27",x"4a"),
   778 => (x"26",x"0f",x"00",x"00"),
   779 => (x"27",x"48",x"70",x"4a"),
   780 => (x"00",x"00",x"16",x"64"),
   781 => (x"93",x"f9",x"c8",x"58"),
   782 => (x"1e",x"72",x"49",x"73"),
   783 => (x"c8",x"27",x"4a",x"72"),
   784 => (x"0f",x"00",x"00",x"04"),
   785 => (x"48",x"70",x"4a",x"26"),
   786 => (x"00",x"17",x"f8",x"27"),
   787 => (x"36",x"27",x"58",x"00"),
   788 => (x"1e",x"00",x"00",x"0f"),
   789 => (x"00",x"01",x"59",x"27"),
   790 => (x"86",x"c4",x"0f",x"00"),
   791 => (x"00",x"16",x"ec",x"27"),
   792 => (x"27",x"1e",x"bf",x"00"),
   793 => (x"00",x"00",x"0f",x"63"),
   794 => (x"01",x"59",x"27",x"1e"),
   795 => (x"c8",x"0f",x"00",x"00"),
   796 => (x"0f",x"68",x"27",x"86"),
   797 => (x"27",x"1e",x"00",x"00"),
   798 => (x"00",x"00",x"01",x"59"),
   799 => (x"27",x"86",x"c4",x"0f"),
   800 => (x"00",x"00",x"16",x"60"),
   801 => (x"95",x"27",x"1e",x"bf"),
   802 => (x"1e",x"00",x"00",x"0f"),
   803 => (x"00",x"01",x"59",x"27"),
   804 => (x"86",x"c8",x"0f",x"00"),
   805 => (x"00",x"17",x"f4",x"27"),
   806 => (x"27",x"1e",x"bf",x"00"),
   807 => (x"00",x"00",x"0f",x"9a"),
   808 => (x"01",x"59",x"27",x"1e"),
   809 => (x"c8",x"0f",x"00",x"00"),
   810 => (x"0f",x"b8",x"27",x"86"),
   811 => (x"27",x"1e",x"00",x"00"),
   812 => (x"00",x"00",x"01",x"59"),
   813 => (x"c0",x"86",x"c4",x"0f"),
   814 => (x"26",x"86",x"d0",x"48"),
   815 => (x"26",x"4c",x"26",x"4d"),
   816 => (x"26",x"4a",x"26",x"4b"),
   817 => (x"5a",x"5e",x"0e",x"4f"),
   818 => (x"0e",x"5d",x"5c",x"5b"),
   819 => (x"bf",x"bf",x"a6",x"d4"),
   820 => (x"27",x"4d",x"72",x"4a"),
   821 => (x"00",x"00",x"16",x"68"),
   822 => (x"1e",x"72",x"48",x"bf"),
   823 => (x"49",x"a2",x"f0",x"c0"),
   824 => (x"a9",x"72",x"52",x"10"),
   825 => (x"26",x"87",x"f9",x"05"),
   826 => (x"4c",x"66",x"d4",x"4a"),
   827 => (x"7c",x"c5",x"84",x"cc"),
   828 => (x"83",x"cc",x"4b",x"72"),
   829 => (x"a6",x"d4",x"7b",x"6c"),
   830 => (x"72",x"7a",x"bf",x"bf"),
   831 => (x"0d",x"a7",x"27",x"1e"),
   832 => (x"c4",x"0f",x"00",x"00"),
   833 => (x"6a",x"82",x"c4",x"86"),
   834 => (x"f4",x"c0",x"05",x"9a"),
   835 => (x"c8",x"4b",x"75",x"87"),
   836 => (x"cc",x"4a",x"75",x"83"),
   837 => (x"73",x"7a",x"c6",x"82"),
   838 => (x"4b",x"66",x"d8",x"1e"),
   839 => (x"1e",x"6b",x"83",x"c8"),
   840 => (x"00",x"02",x"a5",x"27"),
   841 => (x"86",x"c8",x"0f",x"00"),
   842 => (x"00",x"16",x"68",x"27"),
   843 => (x"7d",x"bf",x"bf",x"00"),
   844 => (x"1e",x"ca",x"1e",x"72"),
   845 => (x"24",x"27",x"1e",x"6a"),
   846 => (x"0f",x"00",x"00",x"03"),
   847 => (x"d9",x"c0",x"86",x"cc"),
   848 => (x"bf",x"a6",x"d4",x"87"),
   849 => (x"a6",x"d4",x"4a",x"bf"),
   850 => (x"72",x"48",x"49",x"bf"),
   851 => (x"a1",x"f0",x"c0",x"1e"),
   852 => (x"71",x"51",x"10",x"4a"),
   853 => (x"87",x"f9",x"05",x"aa"),
   854 => (x"4d",x"26",x"4a",x"26"),
   855 => (x"4b",x"26",x"4c",x"26"),
   856 => (x"4f",x"26",x"4a",x"26"),
   857 => (x"5b",x"5a",x"5e",x"0e"),
   858 => (x"a6",x"d0",x"1e",x"0e"),
   859 => (x"ca",x"4b",x"bf",x"bf"),
   860 => (x"16",x"e0",x"27",x"83"),
   861 => (x"bf",x"97",x"00",x"00"),
   862 => (x"b7",x"32",x"d8",x"4a"),
   863 => (x"c1",x"49",x"72",x"2a"),
   864 => (x"05",x"a9",x"b7",x"c1"),
   865 => (x"c1",x"87",x"d4",x"c0"),
   866 => (x"27",x"48",x"73",x"8b"),
   867 => (x"00",x"00",x"17",x"ec"),
   868 => (x"66",x"d0",x"88",x"bf"),
   869 => (x"76",x"79",x"70",x"49"),
   870 => (x"6e",x"79",x"c0",x"49"),
   871 => (x"87",x"d1",x"ff",x"05"),
   872 => (x"26",x"4b",x"26",x"26"),
   873 => (x"1e",x"4f",x"26",x"4a"),
   874 => (x"68",x"27",x"1e",x"72"),
   875 => (x"bf",x"00",x"00",x"16"),
   876 => (x"87",x"cc",x"c0",x"02"),
   877 => (x"49",x"bf",x"a6",x"c8"),
   878 => (x"00",x"16",x"68",x"27"),
   879 => (x"79",x"bf",x"bf",x"00"),
   880 => (x"00",x"16",x"68",x"27"),
   881 => (x"cc",x"4a",x"bf",x"00"),
   882 => (x"27",x"1e",x"72",x"82"),
   883 => (x"00",x"00",x"17",x"ec"),
   884 => (x"1e",x"ca",x"1e",x"bf"),
   885 => (x"00",x"03",x"24",x"27"),
   886 => (x"86",x"cc",x"0f",x"00"),
   887 => (x"4f",x"26",x"4a",x"26"),
   888 => (x"27",x"1e",x"72",x"1e"),
   889 => (x"00",x"00",x"16",x"e0"),
   890 => (x"d8",x"4a",x"bf",x"97"),
   891 => (x"72",x"2a",x"b7",x"32"),
   892 => (x"b7",x"c1",x"c1",x"49"),
   893 => (x"c5",x"c0",x"02",x"a9"),
   894 => (x"c0",x"4a",x"c0",x"87"),
   895 => (x"4a",x"c1",x"87",x"c2"),
   896 => (x"00",x"17",x"f0",x"27"),
   897 => (x"72",x"48",x"bf",x"00"),
   898 => (x"17",x"f4",x"27",x"b0"),
   899 => (x"27",x"58",x"00",x"00"),
   900 => (x"00",x"00",x"17",x"e8"),
   901 => (x"51",x"c2",x"c1",x"49"),
   902 => (x"4f",x"26",x"4a",x"26"),
   903 => (x"16",x"e0",x"27",x"1e"),
   904 => (x"c1",x"49",x"00",x"00"),
   905 => (x"f0",x"27",x"51",x"c1"),
   906 => (x"49",x"00",x"00",x"17"),
   907 => (x"4f",x"26",x"79",x"c0"),
   908 => (x"33",x"32",x"31",x"30"),
   909 => (x"37",x"36",x"35",x"34"),
   910 => (x"42",x"41",x"39",x"38"),
   911 => (x"46",x"45",x"44",x"43"),
   912 => (x"6f",x"72",x"50",x"00"),
   913 => (x"6d",x"61",x"72",x"67"),
   914 => (x"6d",x"6f",x"63",x"20"),
   915 => (x"65",x"6c",x"69",x"70"),
   916 => (x"69",x"77",x"20",x"64"),
   917 => (x"27",x"20",x"68",x"74"),
   918 => (x"69",x"67",x"65",x"72"),
   919 => (x"72",x"65",x"74",x"73"),
   920 => (x"74",x"61",x"20",x"27"),
   921 => (x"62",x"69",x"72",x"74"),
   922 => (x"0a",x"65",x"74",x"75"),
   923 => (x"50",x"00",x"0a",x"00"),
   924 => (x"72",x"67",x"6f",x"72"),
   925 => (x"63",x"20",x"6d",x"61"),
   926 => (x"69",x"70",x"6d",x"6f"),
   927 => (x"20",x"64",x"65",x"6c"),
   928 => (x"68",x"74",x"69",x"77"),
   929 => (x"20",x"74",x"75",x"6f"),
   930 => (x"67",x"65",x"72",x"27"),
   931 => (x"65",x"74",x"73",x"69"),
   932 => (x"61",x"20",x"27",x"72"),
   933 => (x"69",x"72",x"74",x"74"),
   934 => (x"65",x"74",x"75",x"62"),
   935 => (x"00",x"0a",x"00",x"0a"),
   936 => (x"59",x"52",x"48",x"44"),
   937 => (x"4e",x"4f",x"54",x"53"),
   938 => (x"52",x"50",x"20",x"45"),
   939 => (x"41",x"52",x"47",x"4f"),
   940 => (x"33",x"20",x"2c",x"4d"),
   941 => (x"20",x"44",x"52",x"27"),
   942 => (x"49",x"52",x"54",x"53"),
   943 => (x"44",x"00",x"47",x"4e"),
   944 => (x"53",x"59",x"52",x"48"),
   945 => (x"45",x"4e",x"4f",x"54"),
   946 => (x"4f",x"52",x"50",x"20"),
   947 => (x"4d",x"41",x"52",x"47"),
   948 => (x"27",x"32",x"20",x"2c"),
   949 => (x"53",x"20",x"44",x"4e"),
   950 => (x"4e",x"49",x"52",x"54"),
   951 => (x"65",x"4d",x"00",x"47"),
   952 => (x"72",x"75",x"73",x"61"),
   953 => (x"74",x"20",x"64",x"65"),
   954 => (x"20",x"65",x"6d",x"69"),
   955 => (x"20",x"6f",x"6f",x"74"),
   956 => (x"6c",x"61",x"6d",x"73"),
   957 => (x"6f",x"74",x"20",x"6c"),
   958 => (x"74",x"62",x"6f",x"20"),
   959 => (x"20",x"6e",x"69",x"61"),
   960 => (x"6e",x"61",x"65",x"6d"),
   961 => (x"66",x"67",x"6e",x"69"),
   962 => (x"72",x"20",x"6c",x"75"),
   963 => (x"6c",x"75",x"73",x"65"),
   964 => (x"00",x"0a",x"73",x"74"),
   965 => (x"61",x"65",x"6c",x"50"),
   966 => (x"69",x"20",x"65",x"73"),
   967 => (x"65",x"72",x"63",x"6e"),
   968 => (x"20",x"65",x"73",x"61"),
   969 => (x"62",x"6d",x"75",x"6e"),
   970 => (x"6f",x"20",x"72",x"65"),
   971 => (x"75",x"72",x"20",x"66"),
   972 => (x"00",x"0a",x"73",x"6e"),
   973 => (x"69",x"4d",x"00",x"0a"),
   974 => (x"73",x"6f",x"72",x"63"),
   975 => (x"6e",x"6f",x"63",x"65"),
   976 => (x"66",x"20",x"73",x"64"),
   977 => (x"6f",x"20",x"72",x"6f"),
   978 => (x"72",x"20",x"65",x"6e"),
   979 => (x"74",x"20",x"6e",x"75"),
   980 => (x"75",x"6f",x"72",x"68"),
   981 => (x"44",x"20",x"68",x"67"),
   982 => (x"73",x"79",x"72",x"68"),
   983 => (x"65",x"6e",x"6f",x"74"),
   984 => (x"25",x"00",x"20",x"3a"),
   985 => (x"00",x"0a",x"20",x"64"),
   986 => (x"79",x"72",x"68",x"44"),
   987 => (x"6e",x"6f",x"74",x"73"),
   988 => (x"70",x"20",x"73",x"65"),
   989 => (x"53",x"20",x"72",x"65"),
   990 => (x"6e",x"6f",x"63",x"65"),
   991 => (x"20",x"20",x"3a",x"64"),
   992 => (x"20",x"20",x"20",x"20"),
   993 => (x"20",x"20",x"20",x"20"),
   994 => (x"20",x"20",x"20",x"20"),
   995 => (x"20",x"20",x"20",x"20"),
   996 => (x"20",x"20",x"20",x"20"),
   997 => (x"20",x"64",x"25",x"00"),
   998 => (x"41",x"56",x"00",x"0a"),
   999 => (x"49",x"4d",x"20",x"58"),
  1000 => (x"72",x"20",x"53",x"50"),
  1001 => (x"6e",x"69",x"74",x"61"),
  1002 => (x"20",x"2a",x"20",x"67"),
  1003 => (x"30",x"30",x"30",x"31"),
  1004 => (x"25",x"20",x"3d",x"20"),
  1005 => (x"00",x"0a",x"20",x"64"),
  1006 => (x"48",x"44",x"00",x"0a"),
  1007 => (x"54",x"53",x"59",x"52"),
  1008 => (x"20",x"45",x"4e",x"4f"),
  1009 => (x"47",x"4f",x"52",x"50"),
  1010 => (x"2c",x"4d",x"41",x"52"),
  1011 => (x"4d",x"4f",x"53",x"20"),
  1012 => (x"54",x"53",x"20",x"45"),
  1013 => (x"47",x"4e",x"49",x"52"),
  1014 => (x"52",x"48",x"44",x"00"),
  1015 => (x"4f",x"54",x"53",x"59"),
  1016 => (x"50",x"20",x"45",x"4e"),
  1017 => (x"52",x"47",x"4f",x"52"),
  1018 => (x"20",x"2c",x"4d",x"41"),
  1019 => (x"54",x"53",x"27",x"31"),
  1020 => (x"52",x"54",x"53",x"20"),
  1021 => (x"00",x"47",x"4e",x"49"),
  1022 => (x"68",x"44",x"00",x"0a"),
  1023 => (x"74",x"73",x"79",x"72"),
  1024 => (x"20",x"65",x"6e",x"6f"),
  1025 => (x"63",x"6e",x"65",x"42"),
  1026 => (x"72",x"61",x"6d",x"68"),
  1027 => (x"56",x"20",x"2c",x"6b"),
  1028 => (x"69",x"73",x"72",x"65"),
  1029 => (x"32",x"20",x"6e",x"6f"),
  1030 => (x"28",x"20",x"31",x"2e"),
  1031 => (x"67",x"6e",x"61",x"4c"),
  1032 => (x"65",x"67",x"61",x"75"),
  1033 => (x"29",x"43",x"20",x"3a"),
  1034 => (x"00",x"0a",x"00",x"0a"),
  1035 => (x"63",x"65",x"78",x"45"),
  1036 => (x"6f",x"69",x"74",x"75"),
  1037 => (x"74",x"73",x"20",x"6e"),
  1038 => (x"73",x"74",x"72",x"61"),
  1039 => (x"64",x"25",x"20",x"2c"),
  1040 => (x"6e",x"75",x"72",x"20"),
  1041 => (x"68",x"74",x"20",x"73"),
  1042 => (x"67",x"75",x"6f",x"72"),
  1043 => (x"68",x"44",x"20",x"68"),
  1044 => (x"74",x"73",x"79",x"72"),
  1045 => (x"0a",x"65",x"6e",x"6f"),
  1046 => (x"65",x"78",x"45",x"00"),
  1047 => (x"69",x"74",x"75",x"63"),
  1048 => (x"65",x"20",x"6e",x"6f"),
  1049 => (x"0a",x"73",x"64",x"6e"),
  1050 => (x"46",x"00",x"0a",x"00"),
  1051 => (x"6c",x"61",x"6e",x"69"),
  1052 => (x"6c",x"61",x"76",x"20"),
  1053 => (x"20",x"73",x"65",x"75"),
  1054 => (x"74",x"20",x"66",x"6f"),
  1055 => (x"76",x"20",x"65",x"68"),
  1056 => (x"61",x"69",x"72",x"61"),
  1057 => (x"73",x"65",x"6c",x"62"),
  1058 => (x"65",x"73",x"75",x"20"),
  1059 => (x"6e",x"69",x"20",x"64"),
  1060 => (x"65",x"68",x"74",x"20"),
  1061 => (x"6e",x"65",x"62",x"20"),
  1062 => (x"61",x"6d",x"68",x"63"),
  1063 => (x"0a",x"3a",x"6b",x"72"),
  1064 => (x"49",x"00",x"0a",x"00"),
  1065 => (x"47",x"5f",x"74",x"6e"),
  1066 => (x"3a",x"62",x"6f",x"6c"),
  1067 => (x"20",x"20",x"20",x"20"),
  1068 => (x"20",x"20",x"20",x"20"),
  1069 => (x"20",x"20",x"20",x"20"),
  1070 => (x"00",x"0a",x"64",x"25"),
  1071 => (x"20",x"20",x"20",x"20"),
  1072 => (x"20",x"20",x"20",x"20"),
  1073 => (x"75",x"6f",x"68",x"73"),
  1074 => (x"62",x"20",x"64",x"6c"),
  1075 => (x"20",x"20",x"3a",x"65"),
  1076 => (x"0a",x"64",x"25",x"20"),
  1077 => (x"6f",x"6f",x"42",x"00"),
  1078 => (x"6c",x"47",x"5f",x"6c"),
  1079 => (x"20",x"3a",x"62",x"6f"),
  1080 => (x"20",x"20",x"20",x"20"),
  1081 => (x"20",x"20",x"20",x"20"),
  1082 => (x"64",x"25",x"20",x"20"),
  1083 => (x"20",x"20",x"00",x"0a"),
  1084 => (x"20",x"20",x"20",x"20"),
  1085 => (x"68",x"73",x"20",x"20"),
  1086 => (x"64",x"6c",x"75",x"6f"),
  1087 => (x"3a",x"65",x"62",x"20"),
  1088 => (x"25",x"20",x"20",x"20"),
  1089 => (x"43",x"00",x"0a",x"64"),
  1090 => (x"5f",x"31",x"5f",x"68"),
  1091 => (x"62",x"6f",x"6c",x"47"),
  1092 => (x"20",x"20",x"20",x"3a"),
  1093 => (x"20",x"20",x"20",x"20"),
  1094 => (x"20",x"20",x"20",x"20"),
  1095 => (x"00",x"0a",x"63",x"25"),
  1096 => (x"20",x"20",x"20",x"20"),
  1097 => (x"20",x"20",x"20",x"20"),
  1098 => (x"75",x"6f",x"68",x"73"),
  1099 => (x"62",x"20",x"64",x"6c"),
  1100 => (x"20",x"20",x"3a",x"65"),
  1101 => (x"0a",x"63",x"25",x"20"),
  1102 => (x"5f",x"68",x"43",x"00"),
  1103 => (x"6c",x"47",x"5f",x"32"),
  1104 => (x"20",x"3a",x"62",x"6f"),
  1105 => (x"20",x"20",x"20",x"20"),
  1106 => (x"20",x"20",x"20",x"20"),
  1107 => (x"63",x"25",x"20",x"20"),
  1108 => (x"20",x"20",x"00",x"0a"),
  1109 => (x"20",x"20",x"20",x"20"),
  1110 => (x"68",x"73",x"20",x"20"),
  1111 => (x"64",x"6c",x"75",x"6f"),
  1112 => (x"3a",x"65",x"62",x"20"),
  1113 => (x"25",x"20",x"20",x"20"),
  1114 => (x"41",x"00",x"0a",x"63"),
  1115 => (x"31",x"5f",x"72",x"72"),
  1116 => (x"6f",x"6c",x"47",x"5f"),
  1117 => (x"5d",x"38",x"5b",x"62"),
  1118 => (x"20",x"20",x"20",x"3a"),
  1119 => (x"20",x"20",x"20",x"20"),
  1120 => (x"00",x"0a",x"64",x"25"),
  1121 => (x"20",x"20",x"20",x"20"),
  1122 => (x"20",x"20",x"20",x"20"),
  1123 => (x"75",x"6f",x"68",x"73"),
  1124 => (x"62",x"20",x"64",x"6c"),
  1125 => (x"20",x"20",x"3a",x"65"),
  1126 => (x"0a",x"64",x"25",x"20"),
  1127 => (x"72",x"72",x"41",x"00"),
  1128 => (x"47",x"5f",x"32",x"5f"),
  1129 => (x"5b",x"62",x"6f",x"6c"),
  1130 => (x"37",x"5b",x"5d",x"38"),
  1131 => (x"20",x"20",x"3a",x"5d"),
  1132 => (x"64",x"25",x"20",x"20"),
  1133 => (x"20",x"20",x"00",x"0a"),
  1134 => (x"20",x"20",x"20",x"20"),
  1135 => (x"68",x"73",x"20",x"20"),
  1136 => (x"64",x"6c",x"75",x"6f"),
  1137 => (x"3a",x"65",x"62",x"20"),
  1138 => (x"4e",x"20",x"20",x"20"),
  1139 => (x"65",x"62",x"6d",x"75"),
  1140 => (x"66",x"4f",x"5f",x"72"),
  1141 => (x"6e",x"75",x"52",x"5f"),
  1142 => (x"20",x"2b",x"20",x"73"),
  1143 => (x"00",x"0a",x"30",x"31"),
  1144 => (x"5f",x"72",x"74",x"50"),
  1145 => (x"62",x"6f",x"6c",x"47"),
  1146 => (x"00",x"0a",x"3e",x"2d"),
  1147 => (x"74",x"50",x"20",x"20"),
  1148 => (x"6f",x"43",x"5f",x"72"),
  1149 => (x"20",x"3a",x"70",x"6d"),
  1150 => (x"20",x"20",x"20",x"20"),
  1151 => (x"20",x"20",x"20",x"20"),
  1152 => (x"0a",x"64",x"25",x"20"),
  1153 => (x"20",x"20",x"20",x"00"),
  1154 => (x"20",x"20",x"20",x"20"),
  1155 => (x"6f",x"68",x"73",x"20"),
  1156 => (x"20",x"64",x"6c",x"75"),
  1157 => (x"20",x"3a",x"65",x"62"),
  1158 => (x"69",x"28",x"20",x"20"),
  1159 => (x"65",x"6c",x"70",x"6d"),
  1160 => (x"74",x"6e",x"65",x"6d"),
  1161 => (x"6f",x"69",x"74",x"61"),
  1162 => (x"65",x"64",x"2d",x"6e"),
  1163 => (x"64",x"6e",x"65",x"70"),
  1164 => (x"29",x"74",x"6e",x"65"),
  1165 => (x"20",x"20",x"00",x"0a"),
  1166 => (x"63",x"73",x"69",x"44"),
  1167 => (x"20",x"20",x"3a",x"72"),
  1168 => (x"20",x"20",x"20",x"20"),
  1169 => (x"20",x"20",x"20",x"20"),
  1170 => (x"25",x"20",x"20",x"20"),
  1171 => (x"20",x"00",x"0a",x"64"),
  1172 => (x"20",x"20",x"20",x"20"),
  1173 => (x"73",x"20",x"20",x"20"),
  1174 => (x"6c",x"75",x"6f",x"68"),
  1175 => (x"65",x"62",x"20",x"64"),
  1176 => (x"20",x"20",x"20",x"3a"),
  1177 => (x"00",x"0a",x"64",x"25"),
  1178 => (x"6e",x"45",x"20",x"20"),
  1179 => (x"43",x"5f",x"6d",x"75"),
  1180 => (x"3a",x"70",x"6d",x"6f"),
  1181 => (x"20",x"20",x"20",x"20"),
  1182 => (x"20",x"20",x"20",x"20"),
  1183 => (x"0a",x"64",x"25",x"20"),
  1184 => (x"20",x"20",x"20",x"00"),
  1185 => (x"20",x"20",x"20",x"20"),
  1186 => (x"6f",x"68",x"73",x"20"),
  1187 => (x"20",x"64",x"6c",x"75"),
  1188 => (x"20",x"3a",x"65",x"62"),
  1189 => (x"64",x"25",x"20",x"20"),
  1190 => (x"20",x"20",x"00",x"0a"),
  1191 => (x"5f",x"74",x"6e",x"49"),
  1192 => (x"70",x"6d",x"6f",x"43"),
  1193 => (x"20",x"20",x"20",x"3a"),
  1194 => (x"20",x"20",x"20",x"20"),
  1195 => (x"25",x"20",x"20",x"20"),
  1196 => (x"20",x"00",x"0a",x"64"),
  1197 => (x"20",x"20",x"20",x"20"),
  1198 => (x"73",x"20",x"20",x"20"),
  1199 => (x"6c",x"75",x"6f",x"68"),
  1200 => (x"65",x"62",x"20",x"64"),
  1201 => (x"20",x"20",x"20",x"3a"),
  1202 => (x"00",x"0a",x"64",x"25"),
  1203 => (x"74",x"53",x"20",x"20"),
  1204 => (x"6f",x"43",x"5f",x"72"),
  1205 => (x"20",x"3a",x"70",x"6d"),
  1206 => (x"20",x"20",x"20",x"20"),
  1207 => (x"20",x"20",x"20",x"20"),
  1208 => (x"0a",x"73",x"25",x"20"),
  1209 => (x"20",x"20",x"20",x"00"),
  1210 => (x"20",x"20",x"20",x"20"),
  1211 => (x"6f",x"68",x"73",x"20"),
  1212 => (x"20",x"64",x"6c",x"75"),
  1213 => (x"20",x"3a",x"65",x"62"),
  1214 => (x"48",x"44",x"20",x"20"),
  1215 => (x"54",x"53",x"59",x"52"),
  1216 => (x"20",x"45",x"4e",x"4f"),
  1217 => (x"47",x"4f",x"52",x"50"),
  1218 => (x"2c",x"4d",x"41",x"52"),
  1219 => (x"4d",x"4f",x"53",x"20"),
  1220 => (x"54",x"53",x"20",x"45"),
  1221 => (x"47",x"4e",x"49",x"52"),
  1222 => (x"65",x"4e",x"00",x"0a"),
  1223 => (x"50",x"5f",x"74",x"78"),
  1224 => (x"47",x"5f",x"72",x"74"),
  1225 => (x"2d",x"62",x"6f",x"6c"),
  1226 => (x"20",x"00",x"0a",x"3e"),
  1227 => (x"72",x"74",x"50",x"20"),
  1228 => (x"6d",x"6f",x"43",x"5f"),
  1229 => (x"20",x"20",x"3a",x"70"),
  1230 => (x"20",x"20",x"20",x"20"),
  1231 => (x"20",x"20",x"20",x"20"),
  1232 => (x"00",x"0a",x"64",x"25"),
  1233 => (x"20",x"20",x"20",x"20"),
  1234 => (x"20",x"20",x"20",x"20"),
  1235 => (x"75",x"6f",x"68",x"73"),
  1236 => (x"62",x"20",x"64",x"6c"),
  1237 => (x"20",x"20",x"3a",x"65"),
  1238 => (x"6d",x"69",x"28",x"20"),
  1239 => (x"6d",x"65",x"6c",x"70"),
  1240 => (x"61",x"74",x"6e",x"65"),
  1241 => (x"6e",x"6f",x"69",x"74"),
  1242 => (x"70",x"65",x"64",x"2d"),
  1243 => (x"65",x"64",x"6e",x"65"),
  1244 => (x"2c",x"29",x"74",x"6e"),
  1245 => (x"6d",x"61",x"73",x"20"),
  1246 => (x"73",x"61",x"20",x"65"),
  1247 => (x"6f",x"62",x"61",x"20"),
  1248 => (x"00",x"0a",x"65",x"76"),
  1249 => (x"69",x"44",x"20",x"20"),
  1250 => (x"3a",x"72",x"63",x"73"),
  1251 => (x"20",x"20",x"20",x"20"),
  1252 => (x"20",x"20",x"20",x"20"),
  1253 => (x"20",x"20",x"20",x"20"),
  1254 => (x"0a",x"64",x"25",x"20"),
  1255 => (x"20",x"20",x"20",x"00"),
  1256 => (x"20",x"20",x"20",x"20"),
  1257 => (x"6f",x"68",x"73",x"20"),
  1258 => (x"20",x"64",x"6c",x"75"),
  1259 => (x"20",x"3a",x"65",x"62"),
  1260 => (x"64",x"25",x"20",x"20"),
  1261 => (x"20",x"20",x"00",x"0a"),
  1262 => (x"6d",x"75",x"6e",x"45"),
  1263 => (x"6d",x"6f",x"43",x"5f"),
  1264 => (x"20",x"20",x"3a",x"70"),
  1265 => (x"20",x"20",x"20",x"20"),
  1266 => (x"25",x"20",x"20",x"20"),
  1267 => (x"20",x"00",x"0a",x"64"),
  1268 => (x"20",x"20",x"20",x"20"),
  1269 => (x"73",x"20",x"20",x"20"),
  1270 => (x"6c",x"75",x"6f",x"68"),
  1271 => (x"65",x"62",x"20",x"64"),
  1272 => (x"20",x"20",x"20",x"3a"),
  1273 => (x"00",x"0a",x"64",x"25"),
  1274 => (x"6e",x"49",x"20",x"20"),
  1275 => (x"6f",x"43",x"5f",x"74"),
  1276 => (x"20",x"3a",x"70",x"6d"),
  1277 => (x"20",x"20",x"20",x"20"),
  1278 => (x"20",x"20",x"20",x"20"),
  1279 => (x"0a",x"64",x"25",x"20"),
  1280 => (x"20",x"20",x"20",x"00"),
  1281 => (x"20",x"20",x"20",x"20"),
  1282 => (x"6f",x"68",x"73",x"20"),
  1283 => (x"20",x"64",x"6c",x"75"),
  1284 => (x"20",x"3a",x"65",x"62"),
  1285 => (x"64",x"25",x"20",x"20"),
  1286 => (x"20",x"20",x"00",x"0a"),
  1287 => (x"5f",x"72",x"74",x"53"),
  1288 => (x"70",x"6d",x"6f",x"43"),
  1289 => (x"20",x"20",x"20",x"3a"),
  1290 => (x"20",x"20",x"20",x"20"),
  1291 => (x"25",x"20",x"20",x"20"),
  1292 => (x"20",x"00",x"0a",x"73"),
  1293 => (x"20",x"20",x"20",x"20"),
  1294 => (x"73",x"20",x"20",x"20"),
  1295 => (x"6c",x"75",x"6f",x"68"),
  1296 => (x"65",x"62",x"20",x"64"),
  1297 => (x"20",x"20",x"20",x"3a"),
  1298 => (x"59",x"52",x"48",x"44"),
  1299 => (x"4e",x"4f",x"54",x"53"),
  1300 => (x"52",x"50",x"20",x"45"),
  1301 => (x"41",x"52",x"47",x"4f"),
  1302 => (x"53",x"20",x"2c",x"4d"),
  1303 => (x"20",x"45",x"4d",x"4f"),
  1304 => (x"49",x"52",x"54",x"53"),
  1305 => (x"00",x"0a",x"47",x"4e"),
  1306 => (x"5f",x"74",x"6e",x"49"),
  1307 => (x"6f",x"4c",x"5f",x"31"),
  1308 => (x"20",x"20",x"3a",x"63"),
  1309 => (x"20",x"20",x"20",x"20"),
  1310 => (x"20",x"20",x"20",x"20"),
  1311 => (x"0a",x"64",x"25",x"20"),
  1312 => (x"20",x"20",x"20",x"00"),
  1313 => (x"20",x"20",x"20",x"20"),
  1314 => (x"6f",x"68",x"73",x"20"),
  1315 => (x"20",x"64",x"6c",x"75"),
  1316 => (x"20",x"3a",x"65",x"62"),
  1317 => (x"64",x"25",x"20",x"20"),
  1318 => (x"6e",x"49",x"00",x"0a"),
  1319 => (x"5f",x"32",x"5f",x"74"),
  1320 => (x"3a",x"63",x"6f",x"4c"),
  1321 => (x"20",x"20",x"20",x"20"),
  1322 => (x"20",x"20",x"20",x"20"),
  1323 => (x"25",x"20",x"20",x"20"),
  1324 => (x"20",x"00",x"0a",x"64"),
  1325 => (x"20",x"20",x"20",x"20"),
  1326 => (x"73",x"20",x"20",x"20"),
  1327 => (x"6c",x"75",x"6f",x"68"),
  1328 => (x"65",x"62",x"20",x"64"),
  1329 => (x"20",x"20",x"20",x"3a"),
  1330 => (x"00",x"0a",x"64",x"25"),
  1331 => (x"5f",x"74",x"6e",x"49"),
  1332 => (x"6f",x"4c",x"5f",x"33"),
  1333 => (x"20",x"20",x"3a",x"63"),
  1334 => (x"20",x"20",x"20",x"20"),
  1335 => (x"20",x"20",x"20",x"20"),
  1336 => (x"0a",x"64",x"25",x"20"),
  1337 => (x"20",x"20",x"20",x"00"),
  1338 => (x"20",x"20",x"20",x"20"),
  1339 => (x"6f",x"68",x"73",x"20"),
  1340 => (x"20",x"64",x"6c",x"75"),
  1341 => (x"20",x"3a",x"65",x"62"),
  1342 => (x"64",x"25",x"20",x"20"),
  1343 => (x"6e",x"45",x"00",x"0a"),
  1344 => (x"4c",x"5f",x"6d",x"75"),
  1345 => (x"20",x"3a",x"63",x"6f"),
  1346 => (x"20",x"20",x"20",x"20"),
  1347 => (x"20",x"20",x"20",x"20"),
  1348 => (x"25",x"20",x"20",x"20"),
  1349 => (x"20",x"00",x"0a",x"64"),
  1350 => (x"20",x"20",x"20",x"20"),
  1351 => (x"73",x"20",x"20",x"20"),
  1352 => (x"6c",x"75",x"6f",x"68"),
  1353 => (x"65",x"62",x"20",x"64"),
  1354 => (x"20",x"20",x"20",x"3a"),
  1355 => (x"00",x"0a",x"64",x"25"),
  1356 => (x"5f",x"72",x"74",x"53"),
  1357 => (x"6f",x"4c",x"5f",x"31"),
  1358 => (x"20",x"20",x"3a",x"63"),
  1359 => (x"20",x"20",x"20",x"20"),
  1360 => (x"20",x"20",x"20",x"20"),
  1361 => (x"0a",x"73",x"25",x"20"),
  1362 => (x"20",x"20",x"20",x"00"),
  1363 => (x"20",x"20",x"20",x"20"),
  1364 => (x"6f",x"68",x"73",x"20"),
  1365 => (x"20",x"64",x"6c",x"75"),
  1366 => (x"20",x"3a",x"65",x"62"),
  1367 => (x"48",x"44",x"20",x"20"),
  1368 => (x"54",x"53",x"59",x"52"),
  1369 => (x"20",x"45",x"4e",x"4f"),
  1370 => (x"47",x"4f",x"52",x"50"),
  1371 => (x"2c",x"4d",x"41",x"52"),
  1372 => (x"53",x"27",x"31",x"20"),
  1373 => (x"54",x"53",x"20",x"54"),
  1374 => (x"47",x"4e",x"49",x"52"),
  1375 => (x"74",x"53",x"00",x"0a"),
  1376 => (x"5f",x"32",x"5f",x"72"),
  1377 => (x"3a",x"63",x"6f",x"4c"),
  1378 => (x"20",x"20",x"20",x"20"),
  1379 => (x"20",x"20",x"20",x"20"),
  1380 => (x"25",x"20",x"20",x"20"),
  1381 => (x"20",x"00",x"0a",x"73"),
  1382 => (x"20",x"20",x"20",x"20"),
  1383 => (x"73",x"20",x"20",x"20"),
  1384 => (x"6c",x"75",x"6f",x"68"),
  1385 => (x"65",x"62",x"20",x"64"),
  1386 => (x"20",x"20",x"20",x"3a"),
  1387 => (x"59",x"52",x"48",x"44"),
  1388 => (x"4e",x"4f",x"54",x"53"),
  1389 => (x"52",x"50",x"20",x"45"),
  1390 => (x"41",x"52",x"47",x"4f"),
  1391 => (x"32",x"20",x"2c",x"4d"),
  1392 => (x"20",x"44",x"4e",x"27"),
  1393 => (x"49",x"52",x"54",x"53"),
  1394 => (x"00",x"0a",x"47",x"4e"),
  1395 => (x"73",x"55",x"00",x"0a"),
  1396 => (x"74",x"20",x"72",x"65"),
  1397 => (x"3a",x"65",x"6d",x"69"),
  1398 => (x"0a",x"64",x"25",x"20"),
  1399 => (x"00",x"00",x"00",x"00"),
  1400 => (x"61",x"a8",x"00",x"00"),
  1401 => (x"61",x"a8",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
