
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"44",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"36"),
    10 => (x"c0",x"c0",x"c2",x"4f"),
    11 => (x"15",x"00",x"27",x"4e"),
    12 => (x"00",x"0f",x"00",x"00"),
    13 => (x"f0",x"c1",x"87",x"fd"),
    14 => (x"43",x"27",x"4e",x"c0"),
    15 => (x"0f",x"00",x"00",x"00"),
    16 => (x"4f",x"87",x"fd",x"00"),
    17 => (x"ff",x"1e",x"1e",x"4f"),
    18 => (x"48",x"69",x"49",x"c0"),
    19 => (x"c4",x"98",x"c0",x"c4"),
    20 => (x"02",x"6e",x"58",x"a6"),
    21 => (x"c8",x"87",x"f3",x"ff"),
    22 => (x"26",x"48",x"79",x"66"),
    23 => (x"87",x"c6",x"c0",x"c0"),
    24 => (x"4c",x"26",x"4d",x"26"),
    25 => (x"4f",x"26",x"4b",x"26"),
    26 => (x"5c",x"5b",x"5e",x"0e"),
    27 => (x"4c",x"66",x"cc",x"0e"),
    28 => (x"4a",x"14",x"4b",x"c0"),
    29 => (x"c0",x"02",x"9a",x"72"),
    30 => (x"49",x"72",x"87",x"d9"),
    31 => (x"71",x"99",x"ff",x"c3"),
    32 => (x"00",x"45",x"27",x"1e"),
    33 => (x"c4",x"0f",x"00",x"00"),
    34 => (x"14",x"83",x"c1",x"86"),
    35 => (x"05",x"9a",x"72",x"4a"),
    36 => (x"73",x"87",x"e7",x"ff"),
    37 => (x"c9",x"ff",x"ff",x"48"),
    38 => (x"5b",x"5e",x"0e",x"87"),
    39 => (x"f0",x"0e",x"5d",x"5c"),
    40 => (x"c4",x"4b",x"c0",x"86"),
    41 => (x"78",x"c0",x"48",x"a6"),
    42 => (x"4c",x"a6",x"e4",x"c0"),
    43 => (x"49",x"66",x"e0",x"c0"),
    44 => (x"c0",x"80",x"c1",x"48"),
    45 => (x"11",x"58",x"a6",x"e4"),
    46 => (x"b7",x"32",x"d8",x"4a"),
    47 => (x"02",x"9a",x"72",x"2a"),
    48 => (x"c4",x"87",x"ef",x"c4"),
    49 => (x"f9",x"c3",x"02",x"66"),
    50 => (x"48",x"a6",x"c4",x"87"),
    51 => (x"49",x"72",x"78",x"c0"),
    52 => (x"02",x"aa",x"f0",x"c0"),
    53 => (x"c1",x"87",x"c1",x"c3"),
    54 => (x"c3",x"02",x"a9",x"e3"),
    55 => (x"e4",x"c1",x"87",x"c2"),
    56 => (x"e3",x"c0",x"02",x"a9"),
    57 => (x"a9",x"ec",x"c1",x"87"),
    58 => (x"87",x"ec",x"c2",x"02"),
    59 => (x"02",x"a9",x"f0",x"c1"),
    60 => (x"c1",x"87",x"d5",x"c0"),
    61 => (x"c2",x"02",x"a9",x"f3"),
    62 => (x"f5",x"c1",x"87",x"c8"),
    63 => (x"c7",x"c0",x"02",x"a9"),
    64 => (x"a9",x"f8",x"c1",x"87"),
    65 => (x"87",x"ed",x"c2",x"05"),
    66 => (x"49",x"74",x"84",x"c4"),
    67 => (x"48",x"76",x"89",x"c4"),
    68 => (x"02",x"6e",x"78",x"69"),
    69 => (x"c8",x"87",x"db",x"c1"),
    70 => (x"78",x"c0",x"48",x"a6"),
    71 => (x"c0",x"48",x"a6",x"cc"),
    72 => (x"dc",x"49",x"6e",x"78"),
    73 => (x"4a",x"71",x"29",x"b7"),
    74 => (x"48",x"6e",x"9a",x"cf"),
    75 => (x"a6",x"c4",x"30",x"c4"),
    76 => (x"02",x"9a",x"72",x"58"),
    77 => (x"c8",x"87",x"c5",x"c0"),
    78 => (x"78",x"c1",x"48",x"a6"),
    79 => (x"c0",x"06",x"aa",x"c9"),
    80 => (x"f7",x"c0",x"87",x"c6"),
    81 => (x"87",x"c3",x"c0",x"82"),
    82 => (x"c8",x"82",x"f0",x"c0"),
    83 => (x"cc",x"c0",x"02",x"66"),
    84 => (x"27",x"1e",x"72",x"87"),
    85 => (x"00",x"00",x"00",x"45"),
    86 => (x"c1",x"86",x"c4",x"0f"),
    87 => (x"48",x"66",x"cc",x"83"),
    88 => (x"a6",x"d0",x"80",x"c1"),
    89 => (x"48",x"66",x"cc",x"58"),
    90 => (x"04",x"a8",x"b7",x"c8"),
    91 => (x"c1",x"87",x"f2",x"fe"),
    92 => (x"f0",x"c0",x"87",x"e9"),
    93 => (x"00",x"45",x"27",x"1e"),
    94 => (x"c4",x"0f",x"00",x"00"),
    95 => (x"c1",x"83",x"c1",x"86"),
    96 => (x"84",x"c4",x"87",x"d9"),
    97 => (x"89",x"c4",x"49",x"74"),
    98 => (x"68",x"27",x"1e",x"69"),
    99 => (x"0f",x"00",x"00",x"00"),
   100 => (x"49",x"70",x"86",x"c4"),
   101 => (x"87",x"c3",x"c1",x"83"),
   102 => (x"c1",x"48",x"a6",x"c4"),
   103 => (x"87",x"fb",x"c0",x"78"),
   104 => (x"49",x"74",x"84",x"c4"),
   105 => (x"1e",x"69",x"89",x"c4"),
   106 => (x"00",x"00",x"45",x"27"),
   107 => (x"86",x"c4",x"0f",x"00"),
   108 => (x"e6",x"c0",x"83",x"c1"),
   109 => (x"27",x"1e",x"72",x"87"),
   110 => (x"00",x"00",x"00",x"45"),
   111 => (x"c0",x"86",x"c4",x"0f"),
   112 => (x"e5",x"c0",x"87",x"d9"),
   113 => (x"c8",x"c0",x"05",x"aa"),
   114 => (x"48",x"a6",x"c4",x"87"),
   115 => (x"ca",x"c0",x"78",x"c1"),
   116 => (x"27",x"1e",x"72",x"87"),
   117 => (x"00",x"00",x"00",x"45"),
   118 => (x"c0",x"86",x"c4",x"0f"),
   119 => (x"48",x"49",x"66",x"e0"),
   120 => (x"e4",x"c0",x"80",x"c1"),
   121 => (x"4a",x"11",x"58",x"a6"),
   122 => (x"2a",x"b7",x"32",x"d8"),
   123 => (x"fb",x"05",x"9a",x"72"),
   124 => (x"48",x"73",x"87",x"d1"),
   125 => (x"4d",x"26",x"8e",x"f0"),
   126 => (x"4b",x"26",x"4c",x"26"),
   127 => (x"00",x"00",x"4f",x"26"),
   128 => (x"75",x"1e",x"00",x"00"),
   129 => (x"4d",x"d4",x"ff",x"1e"),
   130 => (x"7d",x"49",x"ff",x"c3"),
   131 => (x"38",x"c8",x"48",x"6d"),
   132 => (x"b0",x"6d",x"7d",x"71"),
   133 => (x"7d",x"71",x"38",x"c8"),
   134 => (x"38",x"c8",x"b0",x"6d"),
   135 => (x"b0",x"6d",x"7d",x"71"),
   136 => (x"4d",x"26",x"38",x"c8"),
   137 => (x"75",x"1e",x"4f",x"26"),
   138 => (x"4d",x"d4",x"ff",x"1e"),
   139 => (x"7d",x"49",x"ff",x"c3"),
   140 => (x"30",x"c8",x"48",x"6d"),
   141 => (x"b0",x"6d",x"7d",x"71"),
   142 => (x"7d",x"71",x"30",x"c8"),
   143 => (x"30",x"c8",x"b0",x"6d"),
   144 => (x"b0",x"6d",x"7d",x"71"),
   145 => (x"4f",x"26",x"4d",x"26"),
   146 => (x"ff",x"1e",x"75",x"1e"),
   147 => (x"66",x"cc",x"4d",x"d4"),
   148 => (x"48",x"66",x"c8",x"49"),
   149 => (x"67",x"e6",x"fe",x"7d"),
   150 => (x"07",x"31",x"c9",x"02"),
   151 => (x"7d",x"09",x"39",x"d8"),
   152 => (x"7d",x"09",x"39",x"09"),
   153 => (x"7d",x"09",x"39",x"09"),
   154 => (x"7d",x"09",x"39",x"09"),
   155 => (x"7d",x"70",x"38",x"d0"),
   156 => (x"49",x"c0",x"f1",x"c9"),
   157 => (x"6d",x"48",x"ff",x"c3"),
   158 => (x"c7",x"05",x"a8",x"08"),
   159 => (x"c1",x"7d",x"08",x"87"),
   160 => (x"87",x"f3",x"05",x"89"),
   161 => (x"4f",x"26",x"4d",x"26"),
   162 => (x"49",x"d4",x"ff",x"1e"),
   163 => (x"ff",x"48",x"c8",x"c3"),
   164 => (x"fa",x"05",x"80",x"79"),
   165 => (x"0e",x"4f",x"26",x"87"),
   166 => (x"5c",x"5b",x"5a",x"5e"),
   167 => (x"ff",x"c0",x"0e",x"5d"),
   168 => (x"4d",x"f7",x"c1",x"f0"),
   169 => (x"c0",x"c0",x"c0",x"c1"),
   170 => (x"27",x"4b",x"c0",x"c0"),
   171 => (x"00",x"00",x"02",x"88"),
   172 => (x"df",x"f8",x"c4",x"0f"),
   173 => (x"75",x"1e",x"c0",x"4c"),
   174 => (x"02",x"48",x"27",x"1e"),
   175 => (x"c8",x"0f",x"00",x"00"),
   176 => (x"c1",x"4a",x"70",x"86"),
   177 => (x"c0",x"05",x"aa",x"b7"),
   178 => (x"d4",x"ff",x"87",x"ef"),
   179 => (x"79",x"ff",x"c3",x"49"),
   180 => (x"e1",x"c0",x"1e",x"73"),
   181 => (x"1e",x"e9",x"c1",x"f0"),
   182 => (x"00",x"02",x"48",x"27"),
   183 => (x"86",x"c8",x"0f",x"00"),
   184 => (x"9a",x"72",x"4a",x"70"),
   185 => (x"87",x"cb",x"c0",x"05"),
   186 => (x"c3",x"49",x"d4",x"ff"),
   187 => (x"48",x"c1",x"79",x"ff"),
   188 => (x"27",x"87",x"d0",x"c0"),
   189 => (x"00",x"00",x"02",x"88"),
   190 => (x"74",x"8c",x"c1",x"0f"),
   191 => (x"f4",x"fe",x"05",x"9c"),
   192 => (x"26",x"48",x"c0",x"87"),
   193 => (x"26",x"4c",x"26",x"4d"),
   194 => (x"26",x"4a",x"26",x"4b"),
   195 => (x"5a",x"5e",x"0e",x"4f"),
   196 => (x"c0",x"0e",x"5c",x"5b"),
   197 => (x"c1",x"c1",x"f0",x"ff"),
   198 => (x"49",x"d4",x"ff",x"4c"),
   199 => (x"27",x"79",x"ff",x"c3"),
   200 => (x"00",x"00",x"16",x"40"),
   201 => (x"00",x"68",x"27",x"1e"),
   202 => (x"c4",x"0f",x"00",x"00"),
   203 => (x"c0",x"4b",x"d3",x"86"),
   204 => (x"27",x"1e",x"74",x"1e"),
   205 => (x"00",x"00",x"02",x"48"),
   206 => (x"70",x"86",x"c8",x"0f"),
   207 => (x"05",x"9a",x"72",x"4a"),
   208 => (x"ff",x"87",x"cb",x"c0"),
   209 => (x"ff",x"c3",x"49",x"d4"),
   210 => (x"c0",x"48",x"c1",x"79"),
   211 => (x"88",x"27",x"87",x"d0"),
   212 => (x"0f",x"00",x"00",x"02"),
   213 => (x"9b",x"73",x"8b",x"c1"),
   214 => (x"87",x"d3",x"ff",x"05"),
   215 => (x"4c",x"26",x"48",x"c0"),
   216 => (x"4a",x"26",x"4b",x"26"),
   217 => (x"5e",x"0e",x"4f",x"26"),
   218 => (x"5d",x"5c",x"5b",x"5a"),
   219 => (x"ff",x"c3",x"1e",x"0e"),
   220 => (x"4c",x"d4",x"ff",x"4d"),
   221 => (x"00",x"02",x"88",x"27"),
   222 => (x"ea",x"c6",x"0f",x"00"),
   223 => (x"f0",x"e1",x"c0",x"1e"),
   224 => (x"27",x"1e",x"c8",x"c1"),
   225 => (x"00",x"00",x"02",x"48"),
   226 => (x"70",x"86",x"c8",x"0f"),
   227 => (x"27",x"1e",x"72",x"4a"),
   228 => (x"00",x"00",x"04",x"c5"),
   229 => (x"00",x"99",x"27",x"1e"),
   230 => (x"c8",x"0f",x"00",x"00"),
   231 => (x"aa",x"b7",x"c1",x"86"),
   232 => (x"87",x"cb",x"c0",x"02"),
   233 => (x"00",x"03",x"0d",x"27"),
   234 => (x"48",x"c0",x"0f",x"00"),
   235 => (x"27",x"87",x"c9",x"c3"),
   236 => (x"00",x"00",x"02",x"26"),
   237 => (x"cf",x"4a",x"70",x"0f"),
   238 => (x"c6",x"9a",x"ff",x"ff"),
   239 => (x"02",x"aa",x"b7",x"ea"),
   240 => (x"27",x"87",x"cb",x"c0"),
   241 => (x"00",x"00",x"03",x"0d"),
   242 => (x"c2",x"48",x"c0",x"0f"),
   243 => (x"7c",x"75",x"87",x"ea"),
   244 => (x"f1",x"c0",x"49",x"76"),
   245 => (x"02",x"97",x"27",x"79"),
   246 => (x"70",x"0f",x"00",x"00"),
   247 => (x"02",x"9a",x"72",x"4a"),
   248 => (x"c0",x"87",x"eb",x"c1"),
   249 => (x"f0",x"ff",x"c0",x"1e"),
   250 => (x"27",x"1e",x"fa",x"c1"),
   251 => (x"00",x"00",x"02",x"48"),
   252 => (x"70",x"86",x"c8",x"0f"),
   253 => (x"05",x"9b",x"73",x"4b"),
   254 => (x"73",x"87",x"c3",x"c1"),
   255 => (x"04",x"83",x"27",x"1e"),
   256 => (x"27",x"1e",x"00",x"00"),
   257 => (x"00",x"00",x"00",x"99"),
   258 => (x"75",x"86",x"c8",x"0f"),
   259 => (x"75",x"4b",x"6c",x"7c"),
   260 => (x"27",x"1e",x"73",x"9b"),
   261 => (x"00",x"00",x"04",x"8f"),
   262 => (x"00",x"99",x"27",x"1e"),
   263 => (x"c8",x"0f",x"00",x"00"),
   264 => (x"75",x"7c",x"75",x"86"),
   265 => (x"75",x"7c",x"75",x"7c"),
   266 => (x"c1",x"4a",x"73",x"7c"),
   267 => (x"9a",x"72",x"9a",x"c0"),
   268 => (x"87",x"c5",x"c0",x"02"),
   269 => (x"ff",x"c0",x"48",x"c1"),
   270 => (x"c0",x"48",x"c0",x"87"),
   271 => (x"1e",x"73",x"87",x"fa"),
   272 => (x"00",x"04",x"9d",x"27"),
   273 => (x"99",x"27",x"1e",x"00"),
   274 => (x"0f",x"00",x"00",x"00"),
   275 => (x"49",x"6e",x"86",x"c8"),
   276 => (x"05",x"a9",x"b7",x"c2"),
   277 => (x"27",x"87",x"d3",x"c0"),
   278 => (x"00",x"00",x"04",x"a9"),
   279 => (x"00",x"99",x"27",x"1e"),
   280 => (x"c4",x"0f",x"00",x"00"),
   281 => (x"c0",x"48",x"c0",x"86"),
   282 => (x"48",x"6e",x"87",x"ce"),
   283 => (x"a6",x"c4",x"88",x"c1"),
   284 => (x"fd",x"05",x"6e",x"58"),
   285 => (x"48",x"c0",x"87",x"df"),
   286 => (x"26",x"4d",x"26",x"26"),
   287 => (x"26",x"4b",x"26",x"4c"),
   288 => (x"43",x"4f",x"26",x"4a"),
   289 => (x"38",x"35",x"44",x"4d"),
   290 => (x"0a",x"64",x"25",x"20"),
   291 => (x"43",x"00",x"20",x"20"),
   292 => (x"38",x"35",x"44",x"4d"),
   293 => (x"25",x"20",x"32",x"5f"),
   294 => (x"20",x"20",x"0a",x"64"),
   295 => (x"44",x"4d",x"43",x"00"),
   296 => (x"25",x"20",x"38",x"35"),
   297 => (x"20",x"20",x"0a",x"64"),
   298 => (x"48",x"44",x"53",x"00"),
   299 => (x"6e",x"49",x"20",x"43"),
   300 => (x"61",x"69",x"74",x"69"),
   301 => (x"61",x"7a",x"69",x"6c"),
   302 => (x"6e",x"6f",x"69",x"74"),
   303 => (x"72",x"72",x"65",x"20"),
   304 => (x"0a",x"21",x"72",x"6f"),
   305 => (x"64",x"6d",x"63",x"00"),
   306 => (x"44",x"4d",x"43",x"5f"),
   307 => (x"65",x"72",x"20",x"38"),
   308 => (x"6e",x"6f",x"70",x"73"),
   309 => (x"20",x"3a",x"65",x"73"),
   310 => (x"00",x"0a",x"64",x"25"),
   311 => (x"5b",x"5a",x"5e",x"0e"),
   312 => (x"1e",x"0e",x"5d",x"5c"),
   313 => (x"c8",x"4c",x"d0",x"ff"),
   314 => (x"27",x"4b",x"c0",x"c0"),
   315 => (x"00",x"00",x"01",x"fe"),
   316 => (x"27",x"79",x"c1",x"49"),
   317 => (x"00",x"00",x"05",x"f9"),
   318 => (x"00",x"68",x"27",x"1e"),
   319 => (x"c4",x"0f",x"00",x"00"),
   320 => (x"6c",x"4d",x"c7",x"86"),
   321 => (x"c4",x"98",x"73",x"48"),
   322 => (x"02",x"6e",x"58",x"a6"),
   323 => (x"6c",x"87",x"cc",x"c0"),
   324 => (x"c4",x"98",x"73",x"48"),
   325 => (x"05",x"6e",x"58",x"a6"),
   326 => (x"c0",x"87",x"f4",x"ff"),
   327 => (x"02",x"88",x"27",x"7c"),
   328 => (x"6c",x"0f",x"00",x"00"),
   329 => (x"c4",x"98",x"73",x"48"),
   330 => (x"02",x"6e",x"58",x"a6"),
   331 => (x"6c",x"87",x"cc",x"c0"),
   332 => (x"c4",x"98",x"73",x"48"),
   333 => (x"05",x"6e",x"58",x"a6"),
   334 => (x"c1",x"87",x"f4",x"ff"),
   335 => (x"c0",x"1e",x"c0",x"7c"),
   336 => (x"c0",x"c1",x"d0",x"e5"),
   337 => (x"02",x"48",x"27",x"1e"),
   338 => (x"c8",x"0f",x"00",x"00"),
   339 => (x"c1",x"4a",x"70",x"86"),
   340 => (x"c0",x"05",x"aa",x"b7"),
   341 => (x"4d",x"c1",x"87",x"c2"),
   342 => (x"05",x"ad",x"b7",x"c2"),
   343 => (x"27",x"87",x"d3",x"c0"),
   344 => (x"00",x"00",x"05",x"f4"),
   345 => (x"00",x"68",x"27",x"1e"),
   346 => (x"c4",x"0f",x"00",x"00"),
   347 => (x"c1",x"48",x"c0",x"86"),
   348 => (x"8d",x"c1",x"87",x"f7"),
   349 => (x"fe",x"05",x"9d",x"75"),
   350 => (x"66",x"27",x"87",x"c9"),
   351 => (x"0f",x"00",x"00",x"03"),
   352 => (x"00",x"02",x"02",x"27"),
   353 => (x"fe",x"27",x"58",x"00"),
   354 => (x"bf",x"00",x"00",x"01"),
   355 => (x"87",x"d0",x"c0",x"05"),
   356 => (x"ff",x"c0",x"1e",x"c1"),
   357 => (x"1e",x"d0",x"c1",x"f0"),
   358 => (x"00",x"02",x"48",x"27"),
   359 => (x"86",x"c8",x"0f",x"00"),
   360 => (x"c3",x"49",x"d4",x"ff"),
   361 => (x"8f",x"27",x"79",x"ff"),
   362 => (x"0f",x"00",x"00",x"08"),
   363 => (x"00",x"17",x"e0",x"27"),
   364 => (x"dc",x"27",x"58",x"00"),
   365 => (x"bf",x"00",x"00",x"17"),
   366 => (x"05",x"fd",x"27",x"1e"),
   367 => (x"27",x"1e",x"00",x"00"),
   368 => (x"00",x"00",x"00",x"99"),
   369 => (x"6c",x"86",x"c8",x"0f"),
   370 => (x"c4",x"98",x"73",x"48"),
   371 => (x"02",x"6e",x"58",x"a6"),
   372 => (x"6c",x"87",x"cc",x"c0"),
   373 => (x"c4",x"98",x"73",x"48"),
   374 => (x"05",x"6e",x"58",x"a6"),
   375 => (x"c0",x"87",x"f4",x"ff"),
   376 => (x"49",x"d4",x"ff",x"7c"),
   377 => (x"c1",x"79",x"ff",x"c3"),
   378 => (x"4d",x"26",x"26",x"48"),
   379 => (x"4b",x"26",x"4c",x"26"),
   380 => (x"4f",x"26",x"4a",x"26"),
   381 => (x"52",x"52",x"45",x"49"),
   382 => (x"49",x"50",x"53",x"00"),
   383 => (x"20",x"44",x"53",x"00"),
   384 => (x"64",x"72",x"61",x"63"),
   385 => (x"7a",x"69",x"73",x"20"),
   386 => (x"73",x"69",x"20",x"65"),
   387 => (x"0a",x"64",x"25",x"20"),
   388 => (x"5a",x"5e",x"0e",x"00"),
   389 => (x"0e",x"5d",x"5c",x"5b"),
   390 => (x"4d",x"ff",x"c3",x"1e"),
   391 => (x"75",x"4c",x"d4",x"ff"),
   392 => (x"bf",x"d0",x"ff",x"7c"),
   393 => (x"c0",x"c0",x"c8",x"48"),
   394 => (x"58",x"a6",x"c4",x"98"),
   395 => (x"d2",x"c0",x"02",x"6e"),
   396 => (x"c0",x"c0",x"c8",x"87"),
   397 => (x"bf",x"d0",x"ff",x"4a"),
   398 => (x"c4",x"98",x"72",x"48"),
   399 => (x"05",x"6e",x"58",x"a6"),
   400 => (x"ff",x"87",x"f2",x"ff"),
   401 => (x"c1",x"c4",x"49",x"d0"),
   402 => (x"d8",x"7c",x"75",x"79"),
   403 => (x"ff",x"c0",x"1e",x"66"),
   404 => (x"1e",x"d8",x"c1",x"f0"),
   405 => (x"00",x"02",x"48",x"27"),
   406 => (x"86",x"c8",x"0f",x"00"),
   407 => (x"9a",x"72",x"4a",x"70"),
   408 => (x"87",x"d3",x"c0",x"02"),
   409 => (x"00",x"07",x"19",x"27"),
   410 => (x"68",x"27",x"1e",x"00"),
   411 => (x"0f",x"00",x"00",x"00"),
   412 => (x"48",x"c1",x"86",x"c4"),
   413 => (x"75",x"87",x"d7",x"c2"),
   414 => (x"7c",x"fe",x"c3",x"7c"),
   415 => (x"79",x"c0",x"49",x"76"),
   416 => (x"4a",x"bf",x"66",x"dc"),
   417 => (x"b7",x"d8",x"4b",x"72"),
   418 => (x"75",x"48",x"73",x"2b"),
   419 => (x"72",x"7c",x"70",x"98"),
   420 => (x"2b",x"b7",x"d0",x"4b"),
   421 => (x"98",x"75",x"48",x"73"),
   422 => (x"4b",x"72",x"7c",x"70"),
   423 => (x"73",x"2b",x"b7",x"c8"),
   424 => (x"70",x"98",x"75",x"48"),
   425 => (x"75",x"48",x"72",x"7c"),
   426 => (x"dc",x"7c",x"70",x"98"),
   427 => (x"80",x"c4",x"48",x"66"),
   428 => (x"58",x"a6",x"e0",x"c0"),
   429 => (x"80",x"c1",x"48",x"6e"),
   430 => (x"6e",x"58",x"a6",x"c4"),
   431 => (x"b7",x"c0",x"c2",x"49"),
   432 => (x"fb",x"fe",x"04",x"a9"),
   433 => (x"75",x"7c",x"75",x"87"),
   434 => (x"d8",x"7c",x"75",x"7c"),
   435 => (x"75",x"4b",x"e0",x"da"),
   436 => (x"75",x"4a",x"6c",x"7c"),
   437 => (x"05",x"9a",x"72",x"9a"),
   438 => (x"c1",x"87",x"c8",x"c0"),
   439 => (x"05",x"9b",x"73",x"8b"),
   440 => (x"75",x"87",x"ec",x"ff"),
   441 => (x"bf",x"d0",x"ff",x"7c"),
   442 => (x"c0",x"c0",x"c8",x"48"),
   443 => (x"58",x"a6",x"c4",x"98"),
   444 => (x"d2",x"c0",x"02",x"6e"),
   445 => (x"c0",x"c0",x"c8",x"87"),
   446 => (x"bf",x"d0",x"ff",x"4a"),
   447 => (x"c4",x"98",x"72",x"48"),
   448 => (x"05",x"6e",x"58",x"a6"),
   449 => (x"ff",x"87",x"f2",x"ff"),
   450 => (x"79",x"c0",x"49",x"d0"),
   451 => (x"26",x"26",x"48",x"c0"),
   452 => (x"26",x"4c",x"26",x"4d"),
   453 => (x"26",x"4a",x"26",x"4b"),
   454 => (x"69",x"72",x"57",x"4f"),
   455 => (x"66",x"20",x"65",x"74"),
   456 => (x"65",x"6c",x"69",x"61"),
   457 => (x"0e",x"00",x"0a",x"64"),
   458 => (x"5c",x"5b",x"5a",x"5e"),
   459 => (x"d8",x"1e",x"0e",x"5d"),
   460 => (x"66",x"dc",x"4c",x"66"),
   461 => (x"c0",x"49",x"76",x"4b"),
   462 => (x"cd",x"ee",x"c5",x"79"),
   463 => (x"d4",x"ff",x"4d",x"df"),
   464 => (x"79",x"ff",x"c3",x"49"),
   465 => (x"4a",x"bf",x"d4",x"ff"),
   466 => (x"c3",x"9a",x"ff",x"c3"),
   467 => (x"05",x"aa",x"b7",x"fe"),
   468 => (x"27",x"87",x"e5",x"c1"),
   469 => (x"00",x"00",x"17",x"d8"),
   470 => (x"c4",x"79",x"c0",x"49"),
   471 => (x"c0",x"04",x"ab",x"b7"),
   472 => (x"02",x"27",x"87",x"e4"),
   473 => (x"0f",x"00",x"00",x"02"),
   474 => (x"7c",x"72",x"4a",x"70"),
   475 => (x"d8",x"27",x"84",x"c4"),
   476 => (x"bf",x"00",x"00",x"17"),
   477 => (x"27",x"80",x"72",x"48"),
   478 => (x"00",x"00",x"17",x"dc"),
   479 => (x"c4",x"8b",x"c4",x"58"),
   480 => (x"ff",x"03",x"ab",x"b7"),
   481 => (x"b7",x"c0",x"87",x"dc"),
   482 => (x"e5",x"c0",x"06",x"ab"),
   483 => (x"4d",x"d4",x"ff",x"87"),
   484 => (x"6d",x"7d",x"ff",x"c3"),
   485 => (x"7c",x"97",x"72",x"4a"),
   486 => (x"d8",x"27",x"84",x"c1"),
   487 => (x"bf",x"00",x"00",x"17"),
   488 => (x"27",x"80",x"72",x"48"),
   489 => (x"00",x"00",x"17",x"dc"),
   490 => (x"c0",x"8b",x"c1",x"58"),
   491 => (x"ff",x"01",x"ab",x"b7"),
   492 => (x"4d",x"c1",x"87",x"de"),
   493 => (x"79",x"c1",x"49",x"76"),
   494 => (x"9d",x"75",x"8d",x"c1"),
   495 => (x"87",x"fe",x"fd",x"05"),
   496 => (x"c3",x"49",x"d4",x"ff"),
   497 => (x"48",x"6e",x"79",x"ff"),
   498 => (x"26",x"4d",x"26",x"26"),
   499 => (x"26",x"4b",x"26",x"4c"),
   500 => (x"0e",x"4f",x"26",x"4a"),
   501 => (x"5c",x"5b",x"5a",x"5e"),
   502 => (x"ff",x"1e",x"0e",x"5d"),
   503 => (x"c0",x"c8",x"4b",x"d0"),
   504 => (x"4c",x"c0",x"4a",x"c0"),
   505 => (x"c3",x"49",x"d4",x"ff"),
   506 => (x"48",x"6b",x"79",x"ff"),
   507 => (x"a6",x"c4",x"98",x"72"),
   508 => (x"c0",x"02",x"6e",x"58"),
   509 => (x"48",x"6b",x"87",x"cc"),
   510 => (x"a6",x"c4",x"98",x"72"),
   511 => (x"ff",x"05",x"6e",x"58"),
   512 => (x"c1",x"c4",x"87",x"f4"),
   513 => (x"49",x"d4",x"ff",x"7b"),
   514 => (x"d8",x"79",x"ff",x"c3"),
   515 => (x"ff",x"c0",x"1e",x"66"),
   516 => (x"1e",x"d1",x"c1",x"f0"),
   517 => (x"00",x"02",x"48",x"27"),
   518 => (x"86",x"c8",x"0f",x"00"),
   519 => (x"9d",x"75",x"4d",x"70"),
   520 => (x"87",x"d6",x"c0",x"02"),
   521 => (x"66",x"dc",x"1e",x"75"),
   522 => (x"08",x"6f",x"27",x"1e"),
   523 => (x"27",x"1e",x"00",x"00"),
   524 => (x"00",x"00",x"00",x"99"),
   525 => (x"c0",x"86",x"cc",x"0f"),
   526 => (x"c0",x"c8",x"87",x"e8"),
   527 => (x"66",x"e0",x"c0",x"1e"),
   528 => (x"87",x"e3",x"fb",x"1e"),
   529 => (x"4c",x"70",x"86",x"c8"),
   530 => (x"98",x"72",x"48",x"6b"),
   531 => (x"6e",x"58",x"a6",x"c4"),
   532 => (x"87",x"cc",x"c0",x"02"),
   533 => (x"98",x"72",x"48",x"6b"),
   534 => (x"6e",x"58",x"a6",x"c4"),
   535 => (x"87",x"f4",x"ff",x"05"),
   536 => (x"48",x"74",x"7b",x"c0"),
   537 => (x"26",x"4d",x"26",x"26"),
   538 => (x"26",x"4b",x"26",x"4c"),
   539 => (x"52",x"4f",x"26",x"4a"),
   540 => (x"20",x"64",x"61",x"65"),
   541 => (x"6d",x"6d",x"6f",x"63"),
   542 => (x"20",x"64",x"6e",x"61"),
   543 => (x"6c",x"69",x"61",x"66"),
   544 => (x"61",x"20",x"64",x"65"),
   545 => (x"64",x"25",x"20",x"74"),
   546 => (x"64",x"25",x"28",x"20"),
   547 => (x"0e",x"00",x"0a",x"29"),
   548 => (x"5c",x"5b",x"5a",x"5e"),
   549 => (x"c0",x"1e",x"0e",x"5d"),
   550 => (x"f0",x"ff",x"c0",x"1e"),
   551 => (x"27",x"1e",x"c9",x"c1"),
   552 => (x"00",x"00",x"02",x"48"),
   553 => (x"d2",x"86",x"c8",x"0f"),
   554 => (x"17",x"e8",x"27",x"1e"),
   555 => (x"f9",x"1e",x"00",x"00"),
   556 => (x"86",x"c8",x"87",x"f5"),
   557 => (x"85",x"c1",x"4d",x"c0"),
   558 => (x"04",x"ad",x"b7",x"d2"),
   559 => (x"27",x"87",x"f7",x"ff"),
   560 => (x"00",x"00",x"17",x"e8"),
   561 => (x"c3",x"4a",x"bf",x"97"),
   562 => (x"c0",x"c1",x"9a",x"c0"),
   563 => (x"c0",x"05",x"aa",x"b7"),
   564 => (x"ef",x"27",x"87",x"f2"),
   565 => (x"97",x"00",x"00",x"17"),
   566 => (x"32",x"d0",x"4a",x"bf"),
   567 => (x"00",x"17",x"f0",x"27"),
   568 => (x"4b",x"bf",x"97",x"00"),
   569 => (x"4a",x"72",x"33",x"c8"),
   570 => (x"f1",x"27",x"b2",x"73"),
   571 => (x"97",x"00",x"00",x"17"),
   572 => (x"4a",x"72",x"4b",x"bf"),
   573 => (x"ff",x"cf",x"b2",x"73"),
   574 => (x"72",x"9a",x"ff",x"ff"),
   575 => (x"ca",x"85",x"c1",x"4d"),
   576 => (x"87",x"cb",x"c3",x"35"),
   577 => (x"00",x"17",x"f1",x"27"),
   578 => (x"4a",x"bf",x"97",x"00"),
   579 => (x"9a",x"c6",x"32",x"c1"),
   580 => (x"00",x"17",x"f2",x"27"),
   581 => (x"4b",x"bf",x"97",x"00"),
   582 => (x"72",x"2b",x"b7",x"c7"),
   583 => (x"27",x"b2",x"73",x"4a"),
   584 => (x"00",x"00",x"17",x"ed"),
   585 => (x"73",x"4b",x"bf",x"97"),
   586 => (x"c4",x"98",x"cf",x"48"),
   587 => (x"ee",x"27",x"58",x"a6"),
   588 => (x"97",x"00",x"00",x"17"),
   589 => (x"9b",x"c3",x"4b",x"bf"),
   590 => (x"ef",x"27",x"33",x"ca"),
   591 => (x"97",x"00",x"00",x"17"),
   592 => (x"34",x"c2",x"4c",x"bf"),
   593 => (x"b3",x"74",x"4b",x"73"),
   594 => (x"00",x"17",x"f0",x"27"),
   595 => (x"4c",x"bf",x"97",x"00"),
   596 => (x"c6",x"9c",x"c0",x"c3"),
   597 => (x"4b",x"73",x"2c",x"b7"),
   598 => (x"1e",x"73",x"b3",x"74"),
   599 => (x"72",x"1e",x"66",x"c4"),
   600 => (x"09",x"dc",x"27",x"1e"),
   601 => (x"27",x"1e",x"00",x"00"),
   602 => (x"00",x"00",x"00",x"99"),
   603 => (x"c2",x"86",x"d0",x"0f"),
   604 => (x"72",x"48",x"c1",x"82"),
   605 => (x"72",x"4a",x"70",x"30"),
   606 => (x"0a",x"09",x"27",x"1e"),
   607 => (x"27",x"1e",x"00",x"00"),
   608 => (x"00",x"00",x"00",x"99"),
   609 => (x"c1",x"86",x"c8",x"0f"),
   610 => (x"c4",x"30",x"6e",x"48"),
   611 => (x"83",x"c1",x"58",x"a6"),
   612 => (x"95",x"72",x"4d",x"73"),
   613 => (x"1e",x"75",x"1e",x"6e"),
   614 => (x"00",x"0a",x"12",x"27"),
   615 => (x"99",x"27",x"1e",x"00"),
   616 => (x"0f",x"00",x"00",x"00"),
   617 => (x"49",x"6e",x"86",x"cc"),
   618 => (x"a9",x"b7",x"c0",x"c8"),
   619 => (x"87",x"cf",x"c0",x"06"),
   620 => (x"35",x"c1",x"4a",x"6e"),
   621 => (x"c8",x"2a",x"b7",x"c1"),
   622 => (x"01",x"aa",x"b7",x"c0"),
   623 => (x"75",x"87",x"f3",x"ff"),
   624 => (x"0a",x"28",x"27",x"1e"),
   625 => (x"27",x"1e",x"00",x"00"),
   626 => (x"00",x"00",x"00",x"99"),
   627 => (x"75",x"86",x"c8",x"0f"),
   628 => (x"4d",x"26",x"26",x"48"),
   629 => (x"4b",x"26",x"4c",x"26"),
   630 => (x"4f",x"26",x"4a",x"26"),
   631 => (x"69",x"73",x"5f",x"63"),
   632 => (x"6d",x"5f",x"65",x"7a"),
   633 => (x"3a",x"74",x"6c",x"75"),
   634 => (x"2c",x"64",x"25",x"20"),
   635 => (x"61",x"65",x"72",x"20"),
   636 => (x"6c",x"62",x"5f",x"64"),
   637 => (x"6e",x"65",x"6c",x"5f"),
   638 => (x"64",x"25",x"20",x"3a"),
   639 => (x"73",x"63",x"20",x"2c"),
   640 => (x"3a",x"65",x"7a",x"69"),
   641 => (x"0a",x"64",x"25",x"20"),
   642 => (x"6c",x"75",x"4d",x"00"),
   643 => (x"64",x"25",x"20",x"74"),
   644 => (x"64",x"25",x"00",x"0a"),
   645 => (x"6f",x"6c",x"62",x"20"),
   646 => (x"20",x"73",x"6b",x"63"),
   647 => (x"73",x"20",x"66",x"6f"),
   648 => (x"20",x"65",x"7a",x"69"),
   649 => (x"00",x"0a",x"64",x"25"),
   650 => (x"62",x"20",x"64",x"25"),
   651 => (x"6b",x"63",x"6f",x"6c"),
   652 => (x"66",x"6f",x"20",x"73"),
   653 => (x"32",x"31",x"35",x"20"),
   654 => (x"74",x"79",x"62",x"20"),
   655 => (x"00",x"0a",x"73",x"65"),
   656 => (x"0e",x"5b",x"5e",x"0e"),
   657 => (x"66",x"d0",x"4b",x"c0"),
   658 => (x"a8",x"b7",x"c0",x"48"),
   659 => (x"87",x"f8",x"c0",x"06"),
   660 => (x"bf",x"97",x"66",x"c8"),
   661 => (x"b7",x"32",x"d8",x"4a"),
   662 => (x"48",x"66",x"c8",x"2a"),
   663 => (x"a6",x"cc",x"80",x"c1"),
   664 => (x"97",x"66",x"cc",x"58"),
   665 => (x"31",x"d8",x"49",x"bf"),
   666 => (x"66",x"cc",x"29",x"b7"),
   667 => (x"d0",x"80",x"c1",x"48"),
   668 => (x"b7",x"71",x"58",x"a6"),
   669 => (x"c5",x"c0",x"02",x"aa"),
   670 => (x"c0",x"48",x"c1",x"87"),
   671 => (x"83",x"c1",x"87",x"cc"),
   672 => (x"ab",x"b7",x"66",x"d0"),
   673 => (x"87",x"c8",x"ff",x"04"),
   674 => (x"c0",x"c0",x"48",x"c0"),
   675 => (x"4d",x"26",x"87",x"c4"),
   676 => (x"4b",x"26",x"4c",x"26"),
   677 => (x"5e",x"0e",x"4f",x"26"),
   678 => (x"0e",x"5d",x"5c",x"5b"),
   679 => (x"00",x"1a",x"08",x"27"),
   680 => (x"78",x"c0",x"48",x"00"),
   681 => (x"00",x"17",x"18",x"27"),
   682 => (x"68",x"27",x"1e",x"00"),
   683 => (x"0f",x"00",x"00",x"00"),
   684 => (x"00",x"27",x"86",x"c4"),
   685 => (x"1e",x"00",x"00",x"18"),
   686 => (x"d3",x"27",x"1e",x"c0"),
   687 => (x"0f",x"00",x"00",x"07"),
   688 => (x"98",x"70",x"86",x"c8"),
   689 => (x"87",x"d3",x"c0",x"05"),
   690 => (x"00",x"16",x"44",x"27"),
   691 => (x"68",x"27",x"1e",x"00"),
   692 => (x"0f",x"00",x"00",x"00"),
   693 => (x"48",x"c0",x"86",x"c4"),
   694 => (x"27",x"87",x"d9",x"ce"),
   695 => (x"00",x"00",x"17",x"25"),
   696 => (x"00",x"68",x"27",x"1e"),
   697 => (x"c4",x"0f",x"00",x"00"),
   698 => (x"27",x"4b",x"c0",x"86"),
   699 => (x"00",x"00",x"1a",x"34"),
   700 => (x"c8",x"78",x"c1",x"48"),
   701 => (x"17",x"3c",x"27",x"1e"),
   702 => (x"27",x"1e",x"00",x"00"),
   703 => (x"00",x"00",x"18",x"36"),
   704 => (x"0a",x"40",x"27",x"1e"),
   705 => (x"cc",x"0f",x"00",x"00"),
   706 => (x"05",x"98",x"70",x"86"),
   707 => (x"27",x"87",x"c8",x"c0"),
   708 => (x"00",x"00",x"1a",x"34"),
   709 => (x"c8",x"78",x"c0",x"48"),
   710 => (x"17",x"45",x"27",x"1e"),
   711 => (x"27",x"1e",x"00",x"00"),
   712 => (x"00",x"00",x"18",x"52"),
   713 => (x"0a",x"40",x"27",x"1e"),
   714 => (x"cc",x"0f",x"00",x"00"),
   715 => (x"05",x"98",x"70",x"86"),
   716 => (x"27",x"87",x"c8",x"c0"),
   717 => (x"00",x"00",x"1a",x"34"),
   718 => (x"27",x"78",x"c0",x"48"),
   719 => (x"00",x"00",x"1a",x"34"),
   720 => (x"4e",x"27",x"1e",x"bf"),
   721 => (x"1e",x"00",x"00",x"17"),
   722 => (x"00",x"00",x"99",x"27"),
   723 => (x"86",x"c8",x"0f",x"00"),
   724 => (x"00",x"1a",x"34",x"27"),
   725 => (x"c2",x"02",x"bf",x"00"),
   726 => (x"00",x"27",x"87",x"fc"),
   727 => (x"4d",x"00",x"00",x"18"),
   728 => (x"00",x"19",x"be",x"27"),
   729 => (x"fe",x"27",x"4c",x"00"),
   730 => (x"9f",x"00",x"00",x"19"),
   731 => (x"1e",x"71",x"49",x"bf"),
   732 => (x"00",x"19",x"fe",x"27"),
   733 => (x"00",x"27",x"49",x"00"),
   734 => (x"89",x"00",x"00",x"18"),
   735 => (x"1e",x"d0",x"1e",x"71"),
   736 => (x"27",x"1e",x"c0",x"c8"),
   737 => (x"00",x"00",x"16",x"76"),
   738 => (x"00",x"99",x"27",x"1e"),
   739 => (x"d4",x"0f",x"00",x"00"),
   740 => (x"c8",x"49",x"74",x"86"),
   741 => (x"27",x"4b",x"69",x"81"),
   742 => (x"00",x"00",x"19",x"fe"),
   743 => (x"c5",x"49",x"bf",x"9f"),
   744 => (x"05",x"a9",x"ea",x"d6"),
   745 => (x"74",x"87",x"d3",x"c0"),
   746 => (x"69",x"81",x"c8",x"49"),
   747 => (x"11",x"86",x"27",x"1e"),
   748 => (x"c4",x"0f",x"00",x"00"),
   749 => (x"c0",x"4b",x"70",x"86"),
   750 => (x"49",x"75",x"87",x"e3"),
   751 => (x"9f",x"81",x"fe",x"c7"),
   752 => (x"e9",x"ca",x"49",x"69"),
   753 => (x"c0",x"02",x"a9",x"d5"),
   754 => (x"58",x"27",x"87",x"d3"),
   755 => (x"1e",x"00",x"00",x"16"),
   756 => (x"00",x"00",x"68",x"27"),
   757 => (x"86",x"c4",x"0f",x"00"),
   758 => (x"d7",x"ca",x"48",x"c0"),
   759 => (x"27",x"1e",x"73",x"87"),
   760 => (x"00",x"00",x"16",x"b3"),
   761 => (x"00",x"99",x"27",x"1e"),
   762 => (x"c8",x"0f",x"00",x"00"),
   763 => (x"18",x"00",x"27",x"86"),
   764 => (x"73",x"1e",x"00",x"00"),
   765 => (x"07",x"d3",x"27",x"1e"),
   766 => (x"c8",x"0f",x"00",x"00"),
   767 => (x"05",x"98",x"70",x"86"),
   768 => (x"c0",x"87",x"c5",x"c0"),
   769 => (x"87",x"ec",x"c9",x"48"),
   770 => (x"00",x"16",x"cb",x"27"),
   771 => (x"68",x"27",x"1e",x"00"),
   772 => (x"0f",x"00",x"00",x"00"),
   773 => (x"61",x"27",x"86",x"c4"),
   774 => (x"1e",x"00",x"00",x"17"),
   775 => (x"00",x"00",x"99",x"27"),
   776 => (x"86",x"c4",x"0f",x"00"),
   777 => (x"79",x"27",x"1e",x"c8"),
   778 => (x"1e",x"00",x"00",x"17"),
   779 => (x"00",x"18",x"52",x"27"),
   780 => (x"40",x"27",x"1e",x"00"),
   781 => (x"0f",x"00",x"00",x"0a"),
   782 => (x"98",x"70",x"86",x"cc"),
   783 => (x"87",x"cb",x"c0",x"05"),
   784 => (x"00",x"1a",x"08",x"27"),
   785 => (x"78",x"c1",x"48",x"00"),
   786 => (x"c8",x"87",x"ef",x"c0"),
   787 => (x"17",x"82",x"27",x"1e"),
   788 => (x"27",x"1e",x"00",x"00"),
   789 => (x"00",x"00",x"18",x"36"),
   790 => (x"0a",x"40",x"27",x"1e"),
   791 => (x"cc",x"0f",x"00",x"00"),
   792 => (x"02",x"98",x"70",x"86"),
   793 => (x"27",x"87",x"d3",x"c0"),
   794 => (x"00",x"00",x"16",x"f2"),
   795 => (x"00",x"99",x"27",x"1e"),
   796 => (x"c4",x"0f",x"00",x"00"),
   797 => (x"c7",x"48",x"c0",x"86"),
   798 => (x"fe",x"27",x"87",x"fa"),
   799 => (x"97",x"00",x"00",x"19"),
   800 => (x"d5",x"c1",x"49",x"bf"),
   801 => (x"cf",x"c0",x"05",x"a9"),
   802 => (x"19",x"ff",x"27",x"87"),
   803 => (x"bf",x"97",x"00",x"00"),
   804 => (x"a9",x"ea",x"c2",x"49"),
   805 => (x"87",x"c5",x"c0",x"02"),
   806 => (x"d7",x"c7",x"48",x"c0"),
   807 => (x"18",x"00",x"27",x"87"),
   808 => (x"bf",x"97",x"00",x"00"),
   809 => (x"a9",x"e9",x"c3",x"49"),
   810 => (x"87",x"d4",x"c0",x"02"),
   811 => (x"00",x"18",x"00",x"27"),
   812 => (x"49",x"bf",x"97",x"00"),
   813 => (x"02",x"a9",x"eb",x"c3"),
   814 => (x"c0",x"87",x"c5",x"c0"),
   815 => (x"87",x"f4",x"c6",x"48"),
   816 => (x"00",x"18",x"0b",x"27"),
   817 => (x"49",x"bf",x"97",x"00"),
   818 => (x"c0",x"05",x"99",x"71"),
   819 => (x"0c",x"27",x"87",x"ce"),
   820 => (x"97",x"00",x"00",x"18"),
   821 => (x"a9",x"c2",x"49",x"bf"),
   822 => (x"87",x"c5",x"c0",x"02"),
   823 => (x"d3",x"c6",x"48",x"c0"),
   824 => (x"18",x"0d",x"27",x"87"),
   825 => (x"bf",x"97",x"00",x"00"),
   826 => (x"1a",x"04",x"27",x"48"),
   827 => (x"27",x"58",x"00",x"00"),
   828 => (x"00",x"00",x"1a",x"00"),
   829 => (x"4a",x"71",x"49",x"bf"),
   830 => (x"08",x"27",x"8a",x"c1"),
   831 => (x"5a",x"00",x"00",x"1a"),
   832 => (x"1e",x"71",x"1e",x"72"),
   833 => (x"00",x"17",x"8b",x"27"),
   834 => (x"99",x"27",x"1e",x"00"),
   835 => (x"0f",x"00",x"00",x"00"),
   836 => (x"0e",x"27",x"86",x"cc"),
   837 => (x"97",x"00",x"00",x"18"),
   838 => (x"81",x"73",x"49",x"bf"),
   839 => (x"00",x"18",x"0f",x"27"),
   840 => (x"4a",x"bf",x"97",x"00"),
   841 => (x"48",x"72",x"32",x"c8"),
   842 => (x"18",x"27",x"80",x"71"),
   843 => (x"58",x"00",x"00",x"1a"),
   844 => (x"00",x"18",x"10",x"27"),
   845 => (x"48",x"bf",x"97",x"00"),
   846 => (x"00",x"1a",x"2c",x"27"),
   847 => (x"08",x"27",x"58",x"00"),
   848 => (x"bf",x"00",x"00",x"1a"),
   849 => (x"87",x"c3",x"c3",x"02"),
   850 => (x"0f",x"27",x"1e",x"c8"),
   851 => (x"1e",x"00",x"00",x"17"),
   852 => (x"00",x"18",x"52",x"27"),
   853 => (x"40",x"27",x"1e",x"00"),
   854 => (x"0f",x"00",x"00",x"0a"),
   855 => (x"98",x"70",x"86",x"cc"),
   856 => (x"87",x"c5",x"c0",x"02"),
   857 => (x"cb",x"c4",x"48",x"c0"),
   858 => (x"1a",x"00",x"27",x"87"),
   859 => (x"4a",x"bf",x"00",x"00"),
   860 => (x"30",x"c4",x"48",x"72"),
   861 => (x"00",x"1a",x"30",x"27"),
   862 => (x"28",x"27",x"58",x"00"),
   863 => (x"5a",x"00",x"00",x"1a"),
   864 => (x"00",x"18",x"25",x"27"),
   865 => (x"49",x"bf",x"97",x"00"),
   866 => (x"24",x"27",x"31",x"c8"),
   867 => (x"97",x"00",x"00",x"18"),
   868 => (x"81",x"73",x"4b",x"bf"),
   869 => (x"00",x"18",x"26",x"27"),
   870 => (x"4b",x"bf",x"97",x"00"),
   871 => (x"81",x"73",x"33",x"d0"),
   872 => (x"00",x"18",x"27",x"27"),
   873 => (x"4b",x"bf",x"97",x"00"),
   874 => (x"81",x"73",x"33",x"d8"),
   875 => (x"00",x"1a",x"34",x"27"),
   876 => (x"28",x"27",x"59",x"00"),
   877 => (x"bf",x"00",x"00",x"1a"),
   878 => (x"1a",x"14",x"27",x"91"),
   879 => (x"81",x"bf",x"00",x"00"),
   880 => (x"00",x"1a",x"1c",x"27"),
   881 => (x"2d",x"27",x"59",x"00"),
   882 => (x"97",x"00",x"00",x"18"),
   883 => (x"33",x"c8",x"4b",x"bf"),
   884 => (x"00",x"18",x"2c",x"27"),
   885 => (x"4c",x"bf",x"97",x"00"),
   886 => (x"2e",x"27",x"83",x"74"),
   887 => (x"97",x"00",x"00",x"18"),
   888 => (x"34",x"d0",x"4c",x"bf"),
   889 => (x"2f",x"27",x"83",x"74"),
   890 => (x"97",x"00",x"00",x"18"),
   891 => (x"9c",x"cf",x"4c",x"bf"),
   892 => (x"83",x"74",x"34",x"d8"),
   893 => (x"00",x"1a",x"20",x"27"),
   894 => (x"8b",x"c2",x"5b",x"00"),
   895 => (x"48",x"72",x"92",x"73"),
   896 => (x"24",x"27",x"80",x"71"),
   897 => (x"58",x"00",x"00",x"1a"),
   898 => (x"27",x"87",x"e7",x"c1"),
   899 => (x"00",x"00",x"18",x"12"),
   900 => (x"c8",x"49",x"bf",x"97"),
   901 => (x"18",x"11",x"27",x"31"),
   902 => (x"bf",x"97",x"00",x"00"),
   903 => (x"27",x"81",x"72",x"4a"),
   904 => (x"00",x"00",x"1a",x"30"),
   905 => (x"c7",x"31",x"c5",x"59"),
   906 => (x"29",x"c9",x"81",x"ff"),
   907 => (x"00",x"1a",x"28",x"27"),
   908 => (x"17",x"27",x"59",x"00"),
   909 => (x"97",x"00",x"00",x"18"),
   910 => (x"32",x"c8",x"4a",x"bf"),
   911 => (x"00",x"18",x"16",x"27"),
   912 => (x"4b",x"bf",x"97",x"00"),
   913 => (x"34",x"27",x"82",x"73"),
   914 => (x"5a",x"00",x"00",x"1a"),
   915 => (x"00",x"1a",x"28",x"27"),
   916 => (x"27",x"92",x"bf",x"00"),
   917 => (x"00",x"00",x"1a",x"14"),
   918 => (x"24",x"27",x"82",x"bf"),
   919 => (x"5a",x"00",x"00",x"1a"),
   920 => (x"00",x"1a",x"1c",x"27"),
   921 => (x"78",x"c0",x"48",x"00"),
   922 => (x"80",x"71",x"48",x"72"),
   923 => (x"00",x"1a",x"1c",x"27"),
   924 => (x"48",x"c1",x"58",x"00"),
   925 => (x"87",x"d6",x"f0",x"ff"),
   926 => (x"5c",x"5b",x"5e",x"0e"),
   927 => (x"1a",x"08",x"27",x"0e"),
   928 => (x"02",x"bf",x"00",x"00"),
   929 => (x"cc",x"87",x"cf",x"c0"),
   930 => (x"b7",x"c7",x"4a",x"66"),
   931 => (x"4b",x"66",x"cc",x"2a"),
   932 => (x"c0",x"9b",x"ff",x"c1"),
   933 => (x"66",x"cc",x"87",x"cc"),
   934 => (x"2a",x"b7",x"c8",x"4a"),
   935 => (x"c3",x"4b",x"66",x"cc"),
   936 => (x"00",x"27",x"9b",x"ff"),
   937 => (x"1e",x"00",x"00",x"18"),
   938 => (x"00",x"1a",x"14",x"27"),
   939 => (x"72",x"49",x"bf",x"00"),
   940 => (x"27",x"1e",x"71",x"81"),
   941 => (x"00",x"00",x"07",x"d3"),
   942 => (x"70",x"86",x"c8",x"0f"),
   943 => (x"c5",x"c0",x"05",x"98"),
   944 => (x"c0",x"48",x"c0",x"87"),
   945 => (x"08",x"27",x"87",x"ee"),
   946 => (x"bf",x"00",x"00",x"1a"),
   947 => (x"87",x"d5",x"c0",x"02"),
   948 => (x"91",x"c4",x"49",x"73"),
   949 => (x"00",x"18",x"00",x"27"),
   950 => (x"4c",x"69",x"81",x"00"),
   951 => (x"ff",x"ff",x"ff",x"cf"),
   952 => (x"cd",x"c0",x"9c",x"ff"),
   953 => (x"c2",x"49",x"73",x"87"),
   954 => (x"18",x"00",x"27",x"91"),
   955 => (x"9f",x"81",x"00",x"00"),
   956 => (x"48",x"74",x"4c",x"69"),
   957 => (x"87",x"d8",x"ee",x"ff"),
   958 => (x"5c",x"5b",x"5e",x"0e"),
   959 => (x"86",x"f4",x"0e",x"5d"),
   960 => (x"48",x"76",x"4b",x"c0"),
   961 => (x"00",x"1a",x"1c",x"27"),
   962 => (x"c4",x"78",x"bf",x"00"),
   963 => (x"20",x"27",x"48",x"a6"),
   964 => (x"bf",x"00",x"00",x"1a"),
   965 => (x"1a",x"08",x"27",x"78"),
   966 => (x"02",x"bf",x"00",x"00"),
   967 => (x"27",x"87",x"cc",x"c0"),
   968 => (x"00",x"00",x"1a",x"00"),
   969 => (x"31",x"c4",x"49",x"bf"),
   970 => (x"27",x"87",x"c9",x"c0"),
   971 => (x"00",x"00",x"1a",x"24"),
   972 => (x"31",x"c4",x"49",x"bf"),
   973 => (x"c0",x"59",x"a6",x"cc"),
   974 => (x"48",x"66",x"c8",x"4d"),
   975 => (x"c3",x"06",x"a8",x"c0"),
   976 => (x"49",x"75",x"87",x"c2"),
   977 => (x"99",x"71",x"99",x"cf"),
   978 => (x"87",x"e2",x"c0",x"05"),
   979 => (x"00",x"18",x"00",x"27"),
   980 => (x"66",x"c8",x"1e",x"00"),
   981 => (x"80",x"c1",x"48",x"49"),
   982 => (x"71",x"58",x"a6",x"cc"),
   983 => (x"07",x"d3",x"27",x"1e"),
   984 => (x"c8",x"0f",x"00",x"00"),
   985 => (x"18",x"00",x"27",x"86"),
   986 => (x"c0",x"4b",x"00",x"00"),
   987 => (x"e0",x"c0",x"87",x"c3"),
   988 => (x"49",x"6b",x"97",x"83"),
   989 => (x"c2",x"02",x"99",x"71"),
   990 => (x"6b",x"97",x"87",x"c1"),
   991 => (x"a9",x"e5",x"c3",x"49"),
   992 => (x"87",x"f7",x"c1",x"02"),
   993 => (x"81",x"cb",x"49",x"73"),
   994 => (x"d8",x"49",x"69",x"97"),
   995 => (x"05",x"99",x"71",x"99"),
   996 => (x"73",x"87",x"e8",x"c1"),
   997 => (x"00",x"68",x"27",x"1e"),
   998 => (x"c4",x"0f",x"00",x"00"),
   999 => (x"c0",x"1e",x"cb",x"86"),
  1000 => (x"73",x"1e",x"66",x"e4"),
  1001 => (x"0a",x"40",x"27",x"1e"),
  1002 => (x"cc",x"0f",x"00",x"00"),
  1003 => (x"05",x"98",x"70",x"86"),
  1004 => (x"73",x"87",x"c8",x"c1"),
  1005 => (x"66",x"82",x"dc",x"4a"),
  1006 => (x"6a",x"81",x"c4",x"49"),
  1007 => (x"da",x"4a",x"73",x"79"),
  1008 => (x"49",x"66",x"dc",x"82"),
  1009 => (x"6a",x"9f",x"81",x"c8"),
  1010 => (x"71",x"79",x"70",x"48"),
  1011 => (x"1a",x"08",x"27",x"4c"),
  1012 => (x"02",x"bf",x"00",x"00"),
  1013 => (x"73",x"87",x"d2",x"c0"),
  1014 => (x"9f",x"81",x"d4",x"49"),
  1015 => (x"ff",x"c0",x"49",x"69"),
  1016 => (x"4a",x"71",x"99",x"ff"),
  1017 => (x"c2",x"c0",x"32",x"d0"),
  1018 => (x"72",x"4a",x"c0",x"87"),
  1019 => (x"70",x"80",x"6c",x"48"),
  1020 => (x"48",x"66",x"dc",x"7c"),
  1021 => (x"48",x"c1",x"78",x"c0"),
  1022 => (x"c1",x"87",x"c9",x"c1"),
  1023 => (x"ad",x"66",x"c8",x"85"),
  1024 => (x"87",x"fe",x"fc",x"04"),
  1025 => (x"00",x"1a",x"08",x"27"),
  1026 => (x"c0",x"02",x"bf",x"00"),
  1027 => (x"1e",x"6e",x"87",x"f4"),
  1028 => (x"00",x"0e",x"78",x"27"),
  1029 => (x"86",x"c4",x"0f",x"00"),
  1030 => (x"6e",x"58",x"a6",x"c4"),
  1031 => (x"ff",x"ff",x"cf",x"49"),
  1032 => (x"a9",x"99",x"f8",x"ff"),
  1033 => (x"87",x"da",x"c0",x"02"),
  1034 => (x"89",x"c2",x"49",x"6e"),
  1035 => (x"00",x"1a",x"00",x"27"),
  1036 => (x"27",x"91",x"bf",x"00"),
  1037 => (x"00",x"00",x"1a",x"18"),
  1038 => (x"80",x"71",x"48",x"bf"),
  1039 => (x"fb",x"58",x"a6",x"c8"),
  1040 => (x"48",x"c0",x"87",x"f5"),
  1041 => (x"e9",x"ff",x"8e",x"f4"),
  1042 => (x"73",x"1e",x"87",x"c4"),
  1043 => (x"bf",x"66",x"c8",x"1e"),
  1044 => (x"c8",x"81",x"c1",x"49"),
  1045 => (x"09",x"79",x"09",x"66"),
  1046 => (x"00",x"1a",x"04",x"27"),
  1047 => (x"71",x"99",x"bf",x"00"),
  1048 => (x"d2",x"c0",x"05",x"99"),
  1049 => (x"4b",x"66",x"c8",x"87"),
  1050 => (x"1e",x"6b",x"83",x"c8"),
  1051 => (x"00",x"0e",x"78",x"27"),
  1052 => (x"86",x"c4",x"0f",x"00"),
  1053 => (x"c1",x"7b",x"49",x"70"),
  1054 => (x"d5",x"e8",x"ff",x"48"),
  1055 => (x"18",x"27",x"1e",x"87"),
  1056 => (x"bf",x"00",x"00",x"1a"),
  1057 => (x"4a",x"66",x"c4",x"49"),
  1058 => (x"4a",x"6a",x"82",x"c8"),
  1059 => (x"00",x"27",x"8a",x"c2"),
  1060 => (x"bf",x"00",x"00",x"1a"),
  1061 => (x"27",x"81",x"72",x"92"),
  1062 => (x"00",x"00",x"1a",x"04"),
  1063 => (x"66",x"c4",x"4a",x"bf"),
  1064 => (x"81",x"72",x"9a",x"bf"),
  1065 => (x"71",x"1e",x"66",x"c8"),
  1066 => (x"07",x"d3",x"27",x"1e"),
  1067 => (x"c8",x"0f",x"00",x"00"),
  1068 => (x"05",x"98",x"70",x"86"),
  1069 => (x"c0",x"87",x"c5",x"c0"),
  1070 => (x"87",x"c2",x"c0",x"48"),
  1071 => (x"e7",x"ff",x"48",x"c1"),
  1072 => (x"5e",x"0e",x"87",x"d2"),
  1073 => (x"cc",x"0e",x"5c",x"5b"),
  1074 => (x"38",x"27",x"1e",x"66"),
  1075 => (x"1e",x"00",x"00",x"1a"),
  1076 => (x"00",x"0e",x"f8",x"27"),
  1077 => (x"86",x"c8",x"0f",x"00"),
  1078 => (x"c1",x"02",x"98",x"70"),
  1079 => (x"3c",x"27",x"87",x"e4"),
  1080 => (x"bf",x"00",x"00",x"1a"),
  1081 => (x"81",x"ff",x"c7",x"49"),
  1082 => (x"4c",x"71",x"29",x"c9"),
  1083 => (x"5e",x"27",x"4b",x"c0"),
  1084 => (x"1e",x"00",x"00",x"11"),
  1085 => (x"00",x"00",x"68",x"27"),
  1086 => (x"86",x"c4",x"0f",x"00"),
  1087 => (x"06",x"ac",x"b7",x"c0"),
  1088 => (x"d0",x"87",x"d5",x"c1"),
  1089 => (x"38",x"27",x"1e",x"66"),
  1090 => (x"1e",x"00",x"00",x"1a"),
  1091 => (x"00",x"10",x"7d",x"27"),
  1092 => (x"86",x"c8",x"0f",x"00"),
  1093 => (x"c0",x"05",x"98",x"70"),
  1094 => (x"48",x"c0",x"87",x"c5"),
  1095 => (x"27",x"87",x"fb",x"c0"),
  1096 => (x"00",x"00",x"1a",x"38"),
  1097 => (x"10",x"4a",x"27",x"1e"),
  1098 => (x"c4",x"0f",x"00",x"00"),
  1099 => (x"48",x"66",x"d0",x"86"),
  1100 => (x"d4",x"80",x"c0",x"c8"),
  1101 => (x"83",x"c1",x"58",x"a6"),
  1102 => (x"04",x"ab",x"b7",x"74"),
  1103 => (x"c0",x"87",x"c4",x"ff"),
  1104 => (x"66",x"cc",x"87",x"d6"),
  1105 => (x"11",x"77",x"27",x"1e"),
  1106 => (x"27",x"1e",x"00",x"00"),
  1107 => (x"00",x"00",x"00",x"99"),
  1108 => (x"c0",x"86",x"c8",x"0f"),
  1109 => (x"87",x"c2",x"c0",x"48"),
  1110 => (x"e4",x"ff",x"48",x"c1"),
  1111 => (x"70",x"4f",x"87",x"f2"),
  1112 => (x"64",x"65",x"6e",x"65"),
  1113 => (x"6c",x"69",x"66",x"20"),
  1114 => (x"6c",x"20",x"2c",x"65"),
  1115 => (x"69",x"64",x"61",x"6f"),
  1116 => (x"2e",x"2e",x"67",x"6e"),
  1117 => (x"43",x"00",x"0a",x"2e"),
  1118 => (x"74",x"27",x"6e",x"61"),
  1119 => (x"65",x"70",x"6f",x"20"),
  1120 => (x"73",x"25",x"20",x"6e"),
  1121 => (x"c4",x"1e",x"00",x"0a"),
  1122 => (x"29",x"d8",x"49",x"66"),
  1123 => (x"c4",x"99",x"ff",x"c3"),
  1124 => (x"2a",x"c8",x"4a",x"66"),
  1125 => (x"9a",x"c0",x"fc",x"cf"),
  1126 => (x"66",x"c4",x"b1",x"72"),
  1127 => (x"c0",x"32",x"c8",x"4a"),
  1128 => (x"c0",x"c0",x"f0",x"ff"),
  1129 => (x"c4",x"b1",x"72",x"9a"),
  1130 => (x"32",x"d8",x"4a",x"66"),
  1131 => (x"c0",x"c0",x"c0",x"ff"),
  1132 => (x"b1",x"72",x"9a",x"c0"),
  1133 => (x"c0",x"c0",x"48",x"71"),
  1134 => (x"4d",x"26",x"87",x"c6"),
  1135 => (x"4b",x"26",x"4c",x"26"),
  1136 => (x"c4",x"1e",x"4f",x"26"),
  1137 => (x"2a",x"c8",x"4a",x"66"),
  1138 => (x"72",x"9a",x"ff",x"c3"),
  1139 => (x"49",x"66",x"c4",x"4a"),
  1140 => (x"fc",x"cf",x"31",x"c8"),
  1141 => (x"ff",x"cf",x"99",x"c0"),
  1142 => (x"b1",x"72",x"9a",x"ff"),
  1143 => (x"ff",x"cf",x"49",x"71"),
  1144 => (x"48",x"71",x"99",x"ff"),
  1145 => (x"87",x"d8",x"ff",x"ff"),
  1146 => (x"49",x"66",x"c4",x"1e"),
  1147 => (x"ff",x"cf",x"29",x"d0"),
  1148 => (x"49",x"71",x"99",x"ff"),
  1149 => (x"d0",x"4a",x"66",x"c4"),
  1150 => (x"c0",x"c0",x"f0",x"32"),
  1151 => (x"71",x"b1",x"72",x"9a"),
  1152 => (x"fb",x"fe",x"ff",x"48"),
  1153 => (x"1e",x"73",x"1e",x"87"),
  1154 => (x"c0",x"c0",x"c0",x"d0"),
  1155 => (x"0f",x"73",x"4b",x"c0"),
  1156 => (x"c0",x"87",x"fd",x"ff"),
  1157 => (x"26",x"87",x"c4",x"c0"),
  1158 => (x"26",x"4c",x"26",x"4d"),
  1159 => (x"1e",x"4f",x"26",x"4b"),
  1160 => (x"c3",x"49",x"66",x"c8"),
  1161 => (x"f7",x"c0",x"99",x"df"),
  1162 => (x"a9",x"b7",x"c0",x"89"),
  1163 => (x"87",x"c3",x"c0",x"03"),
  1164 => (x"c4",x"81",x"e7",x"c0"),
  1165 => (x"30",x"c4",x"48",x"66"),
  1166 => (x"c4",x"58",x"a6",x"c8"),
  1167 => (x"b0",x"71",x"48",x"66"),
  1168 => (x"c4",x"58",x"a6",x"c8"),
  1169 => (x"ff",x"ff",x"48",x"66"),
  1170 => (x"5e",x"0e",x"87",x"d3"),
  1171 => (x"d0",x"0e",x"5c",x"5b"),
  1172 => (x"c0",x"c0",x"c0",x"c0"),
  1173 => (x"1a",x"44",x"27",x"4c"),
  1174 => (x"48",x"bf",x"00",x"00"),
  1175 => (x"48",x"27",x"80",x"c1"),
  1176 => (x"58",x"00",x"00",x"1a"),
  1177 => (x"49",x"66",x"cc",x"97"),
  1178 => (x"29",x"b7",x"31",x"d8"),
  1179 => (x"05",x"a9",x"d3",x"c1"),
  1180 => (x"27",x"87",x"e9",x"c0"),
  1181 => (x"00",x"00",x"1a",x"44"),
  1182 => (x"27",x"78",x"c0",x"48"),
  1183 => (x"00",x"00",x"1a",x"48"),
  1184 => (x"27",x"78",x"c0",x"48"),
  1185 => (x"00",x"00",x"1a",x"50"),
  1186 => (x"27",x"78",x"c0",x"48"),
  1187 => (x"00",x"00",x"1a",x"54"),
  1188 => (x"ff",x"78",x"c0",x"48"),
  1189 => (x"d3",x"c1",x"48",x"c0"),
  1190 => (x"87",x"e0",x"c9",x"78"),
  1191 => (x"00",x"1a",x"44",x"27"),
  1192 => (x"c1",x"48",x"bf",x"00"),
  1193 => (x"d4",x"c1",x"05",x"a8"),
  1194 => (x"48",x"c0",x"ff",x"87"),
  1195 => (x"97",x"78",x"f4",x"c1"),
  1196 => (x"d8",x"49",x"66",x"cc"),
  1197 => (x"71",x"29",x"b7",x"31"),
  1198 => (x"1a",x"54",x"27",x"1e"),
  1199 => (x"1e",x"bf",x"00",x"00"),
  1200 => (x"00",x"12",x"1f",x"27"),
  1201 => (x"86",x"c8",x"0f",x"00"),
  1202 => (x"00",x"1a",x"58",x"27"),
  1203 => (x"54",x"27",x"58",x"00"),
  1204 => (x"bf",x"00",x"00",x"1a"),
  1205 => (x"aa",x"b7",x"c3",x"4a"),
  1206 => (x"87",x"c6",x"c0",x"06"),
  1207 => (x"88",x"72",x"48",x"ca"),
  1208 => (x"49",x"72",x"4a",x"70"),
  1209 => (x"48",x"71",x"81",x"c1"),
  1210 => (x"50",x"27",x"30",x"c1"),
  1211 => (x"58",x"00",x"00",x"1a"),
  1212 => (x"f0",x"c0",x"48",x"72"),
  1213 => (x"08",x"c0",x"ff",x"80"),
  1214 => (x"ff",x"c7",x"08",x"78"),
  1215 => (x"1a",x"54",x"27",x"87"),
  1216 => (x"48",x"bf",x"00",x"00"),
  1217 => (x"01",x"a8",x"b7",x"c9"),
  1218 => (x"27",x"87",x"f1",x"c7"),
  1219 => (x"00",x"00",x"1a",x"54"),
  1220 => (x"b7",x"c0",x"48",x"bf"),
  1221 => (x"e3",x"c7",x"06",x"a8"),
  1222 => (x"1a",x"54",x"27",x"87"),
  1223 => (x"48",x"bf",x"00",x"00"),
  1224 => (x"ff",x"80",x"f0",x"c0"),
  1225 => (x"08",x"78",x"08",x"c0"),
  1226 => (x"00",x"1a",x"44",x"27"),
  1227 => (x"c3",x"48",x"bf",x"00"),
  1228 => (x"c0",x"01",x"a8",x"b7"),
  1229 => (x"cc",x"97",x"87",x"e2"),
  1230 => (x"31",x"d8",x"49",x"66"),
  1231 => (x"1e",x"71",x"29",x"b7"),
  1232 => (x"00",x"1a",x"50",x"27"),
  1233 => (x"27",x"1e",x"bf",x"00"),
  1234 => (x"00",x"00",x"12",x"1f"),
  1235 => (x"27",x"86",x"c8",x"0f"),
  1236 => (x"00",x"00",x"1a",x"54"),
  1237 => (x"87",x"e4",x"c6",x"58"),
  1238 => (x"00",x"1a",x"4c",x"27"),
  1239 => (x"c3",x"49",x"bf",x"00"),
  1240 => (x"1a",x"44",x"27",x"81"),
  1241 => (x"b7",x"bf",x"00",x"00"),
  1242 => (x"ea",x"c0",x"04",x"a9"),
  1243 => (x"66",x"cc",x"97",x"87"),
  1244 => (x"b7",x"31",x"d8",x"49"),
  1245 => (x"27",x"1e",x"71",x"29"),
  1246 => (x"00",x"00",x"1a",x"48"),
  1247 => (x"1f",x"27",x"1e",x"bf"),
  1248 => (x"0f",x"00",x"00",x"12"),
  1249 => (x"4c",x"27",x"86",x"c8"),
  1250 => (x"58",x"00",x"00",x"1a"),
  1251 => (x"00",x"1a",x"58",x"27"),
  1252 => (x"78",x"c1",x"48",x"00"),
  1253 => (x"27",x"87",x"e5",x"c5"),
  1254 => (x"00",x"00",x"1a",x"54"),
  1255 => (x"b7",x"c0",x"48",x"bf"),
  1256 => (x"c1",x"c3",x"06",x"a8"),
  1257 => (x"1a",x"54",x"27",x"87"),
  1258 => (x"48",x"bf",x"00",x"00"),
  1259 => (x"01",x"a8",x"b7",x"c3"),
  1260 => (x"27",x"87",x"f3",x"c2"),
  1261 => (x"00",x"00",x"1a",x"50"),
  1262 => (x"31",x"c1",x"49",x"bf"),
  1263 => (x"1a",x"44",x"27",x"81"),
  1264 => (x"b7",x"bf",x"00",x"00"),
  1265 => (x"f7",x"c1",x"04",x"a9"),
  1266 => (x"66",x"cc",x"97",x"87"),
  1267 => (x"b7",x"31",x"d8",x"49"),
  1268 => (x"27",x"1e",x"71",x"29"),
  1269 => (x"00",x"00",x"1a",x"5c"),
  1270 => (x"1f",x"27",x"1e",x"bf"),
  1271 => (x"0f",x"00",x"00",x"12"),
  1272 => (x"60",x"27",x"86",x"c8"),
  1273 => (x"58",x"00",x"00",x"1a"),
  1274 => (x"00",x"1a",x"58",x"27"),
  1275 => (x"c1",x"49",x"bf",x"00"),
  1276 => (x"1a",x"5c",x"27",x"89"),
  1277 => (x"c0",x"59",x"00",x"00"),
  1278 => (x"c3",x"03",x"a9",x"b7"),
  1279 => (x"48",x"27",x"87",x"fe"),
  1280 => (x"bf",x"00",x"00",x"1a"),
  1281 => (x"1a",x"5c",x"27",x"49"),
  1282 => (x"bf",x"97",x"00",x"00"),
  1283 => (x"1a",x"48",x"27",x"51"),
  1284 => (x"49",x"bf",x"00",x"00"),
  1285 => (x"4c",x"27",x"81",x"c1"),
  1286 => (x"59",x"00",x"00",x"1a"),
  1287 => (x"00",x"1a",x"60",x"27"),
  1288 => (x"a9",x"b7",x"bf",x"00"),
  1289 => (x"87",x"cd",x"c0",x"06"),
  1290 => (x"00",x"1a",x"60",x"27"),
  1291 => (x"48",x"27",x"48",x"00"),
  1292 => (x"bf",x"00",x"00",x"1a"),
  1293 => (x"1a",x"58",x"27",x"78"),
  1294 => (x"c1",x"48",x"00",x"00"),
  1295 => (x"87",x"fc",x"c2",x"78"),
  1296 => (x"00",x"1a",x"58",x"27"),
  1297 => (x"c2",x"05",x"bf",x"00"),
  1298 => (x"5c",x"27",x"87",x"f2"),
  1299 => (x"bf",x"00",x"00",x"1a"),
  1300 => (x"27",x"31",x"c4",x"49"),
  1301 => (x"00",x"00",x"1a",x"60"),
  1302 => (x"1a",x"48",x"27",x"59"),
  1303 => (x"09",x"bf",x"00",x"00"),
  1304 => (x"c2",x"09",x"79",x"97"),
  1305 => (x"54",x"27",x"87",x"d6"),
  1306 => (x"bf",x"00",x"00",x"1a"),
  1307 => (x"a8",x"b7",x"c7",x"48"),
  1308 => (x"87",x"f9",x"c1",x"04"),
  1309 => (x"f4",x"fe",x"4b",x"c0"),
  1310 => (x"27",x"78",x"c1",x"48"),
  1311 => (x"00",x"00",x"1a",x"60"),
  1312 => (x"1e",x"74",x"1e",x"bf"),
  1313 => (x"00",x"17",x"af",x"27"),
  1314 => (x"99",x"27",x"1e",x"00"),
  1315 => (x"0f",x"00",x"00",x"00"),
  1316 => (x"4c",x"27",x"86",x"cc"),
  1317 => (x"5c",x"00",x"00",x"1a"),
  1318 => (x"00",x"1a",x"48",x"27"),
  1319 => (x"27",x"48",x"bf",x"00"),
  1320 => (x"00",x"00",x"1a",x"60"),
  1321 => (x"03",x"a8",x"b7",x"bf"),
  1322 => (x"27",x"87",x"e3",x"c0"),
  1323 => (x"00",x"00",x"1a",x"48"),
  1324 => (x"27",x"83",x"bf",x"bf"),
  1325 => (x"00",x"00",x"1a",x"48"),
  1326 => (x"81",x"c4",x"49",x"bf"),
  1327 => (x"00",x"1a",x"4c",x"27"),
  1328 => (x"60",x"27",x"59",x"00"),
  1329 => (x"bf",x"00",x"00",x"1a"),
  1330 => (x"ff",x"04",x"a9",x"b7"),
  1331 => (x"1e",x"73",x"87",x"dd"),
  1332 => (x"00",x"17",x"ce",x"27"),
  1333 => (x"99",x"27",x"1e",x"00"),
  1334 => (x"0f",x"00",x"00",x"00"),
  1335 => (x"c0",x"ff",x"86",x"c8"),
  1336 => (x"78",x"c2",x"c1",x"48"),
  1337 => (x"00",x"12",x"05",x"27"),
  1338 => (x"cf",x"c0",x"0f",x"00"),
  1339 => (x"1a",x"54",x"27",x"87"),
  1340 => (x"48",x"bf",x"00",x"00"),
  1341 => (x"ff",x"80",x"f0",x"c0"),
  1342 => (x"08",x"78",x"08",x"c0"),
  1343 => (x"87",x"d9",x"f4",x"ff"),
  1344 => (x"5c",x"5b",x"5e",x"0e"),
  1345 => (x"02",x"27",x"0e",x"5d"),
  1346 => (x"1e",x"00",x"00",x"16"),
  1347 => (x"00",x"00",x"68",x"27"),
  1348 => (x"86",x"c4",x"0f",x"00"),
  1349 => (x"00",x"04",x"dc",x"27"),
  1350 => (x"98",x"70",x"0f",x"00"),
  1351 => (x"87",x"d1",x"c0",x"02"),
  1352 => (x"00",x"0a",x"96",x"27"),
  1353 => (x"98",x"70",x"0f",x"00"),
  1354 => (x"87",x"c5",x"c0",x"02"),
  1355 => (x"c2",x"c0",x"49",x"c1"),
  1356 => (x"71",x"49",x"c0",x"87"),
  1357 => (x"16",x"18",x"27",x"4d"),
  1358 => (x"27",x"1e",x"00",x"00"),
  1359 => (x"00",x"00",x"00",x"68"),
  1360 => (x"27",x"86",x"c4",x"0f"),
  1361 => (x"00",x"00",x"1a",x"60"),
  1362 => (x"c0",x"78",x"c0",x"48"),
  1363 => (x"45",x"27",x"1e",x"ee"),
  1364 => (x"0f",x"00",x"00",x"00"),
  1365 => (x"f4",x"c3",x"86",x"c4"),
  1366 => (x"ff",x"4a",x"ff",x"c8"),
  1367 => (x"74",x"4c",x"bf",x"c0"),
  1368 => (x"99",x"c0",x"c8",x"49"),
  1369 => (x"c1",x"02",x"99",x"71"),
  1370 => (x"4b",x"74",x"87",x"df"),
  1371 => (x"db",x"9b",x"ff",x"c3"),
  1372 => (x"c5",x"c1",x"05",x"ab"),
  1373 => (x"02",x"9d",x"75",x"87"),
  1374 => (x"d0",x"87",x"f1",x"c0"),
  1375 => (x"c0",x"c0",x"c0",x"c0"),
  1376 => (x"15",x"e6",x"27",x"1e"),
  1377 => (x"27",x"1e",x"00",x"00"),
  1378 => (x"00",x"00",x"10",x"c2"),
  1379 => (x"70",x"86",x"c8",x"0f"),
  1380 => (x"d7",x"c0",x"02",x"98"),
  1381 => (x"15",x"da",x"27",x"87"),
  1382 => (x"27",x"1e",x"00",x"00"),
  1383 => (x"00",x"00",x"00",x"68"),
  1384 => (x"27",x"86",x"c4",x"0f"),
  1385 => (x"00",x"00",x"12",x"05"),
  1386 => (x"87",x"ce",x"c0",x"0f"),
  1387 => (x"00",x"15",x"f2",x"27"),
  1388 => (x"68",x"27",x"1e",x"00"),
  1389 => (x"0f",x"00",x"00",x"00"),
  1390 => (x"1e",x"73",x"86",x"c4"),
  1391 => (x"00",x"12",x"4a",x"27"),
  1392 => (x"86",x"c4",x"0f",x"00"),
  1393 => (x"c0",x"c9",x"f4",x"c3"),
  1394 => (x"c1",x"49",x"72",x"4a"),
  1395 => (x"05",x"99",x"71",x"8a"),
  1396 => (x"fd",x"87",x"c8",x"fe"),
  1397 => (x"f0",x"ff",x"87",x"f5"),
  1398 => (x"6f",x"42",x"87",x"fd"),
  1399 => (x"6e",x"69",x"74",x"6f"),
  1400 => (x"2e",x"2e",x"2e",x"67"),
  1401 => (x"4f",x"42",x"00",x"0a"),
  1402 => (x"33",x"38",x"54",x"4f"),
  1403 => (x"49",x"42",x"20",x"32"),
  1404 => (x"44",x"53",x"00",x"4e"),
  1405 => (x"6f",x"6f",x"62",x"20"),
  1406 => (x"61",x"66",x"20",x"74"),
  1407 => (x"64",x"65",x"6c",x"69"),
  1408 => (x"6e",x"49",x"00",x"0a"),
  1409 => (x"61",x"69",x"74",x"69"),
  1410 => (x"69",x"7a",x"69",x"6c"),
  1411 => (x"53",x"20",x"67",x"6e"),
  1412 => (x"61",x"63",x"20",x"44"),
  1413 => (x"00",x"0a",x"64",x"72"),
  1414 => (x"33",x"32",x"53",x"52"),
  1415 => (x"6f",x"62",x"20",x"32"),
  1416 => (x"2d",x"20",x"74",x"6f"),
  1417 => (x"65",x"72",x"70",x"20"),
  1418 => (x"45",x"20",x"73",x"73"),
  1419 => (x"74",x"20",x"43",x"53"),
  1420 => (x"6f",x"62",x"20",x"6f"),
  1421 => (x"66",x"20",x"74",x"6f"),
  1422 => (x"20",x"6d",x"6f",x"72"),
  1423 => (x"00",x"2e",x"44",x"53"),
  1424 => (x"00",x"44",x"4d",x"43"),
  1425 => (x"64",x"61",x"65",x"52"),
  1426 => (x"20",x"66",x"6f",x"20"),
  1427 => (x"20",x"52",x"42",x"4d"),
  1428 => (x"6c",x"69",x"61",x"66"),
  1429 => (x"00",x"0a",x"64",x"65"),
  1430 => (x"70",x"20",x"6f",x"4e"),
  1431 => (x"69",x"74",x"72",x"61"),
  1432 => (x"6e",x"6f",x"69",x"74"),
  1433 => (x"67",x"69",x"73",x"20"),
  1434 => (x"75",x"74",x"61",x"6e"),
  1435 => (x"66",x"20",x"65",x"72"),
  1436 => (x"64",x"6e",x"75",x"6f"),
  1437 => (x"42",x"4d",x"00",x"0a"),
  1438 => (x"7a",x"69",x"73",x"52"),
  1439 => (x"25",x"20",x"3a",x"65"),
  1440 => (x"70",x"20",x"2c",x"64"),
  1441 => (x"69",x"74",x"72",x"61"),
  1442 => (x"6e",x"6f",x"69",x"74"),
  1443 => (x"65",x"7a",x"69",x"73"),
  1444 => (x"64",x"25",x"20",x"3a"),
  1445 => (x"66",x"6f",x"20",x"2c"),
  1446 => (x"74",x"65",x"73",x"66"),
  1447 => (x"20",x"66",x"6f",x"20"),
  1448 => (x"3a",x"67",x"69",x"73"),
  1449 => (x"2c",x"64",x"25",x"20"),
  1450 => (x"67",x"69",x"73",x"20"),
  1451 => (x"25",x"78",x"30",x"20"),
  1452 => (x"52",x"00",x"0a",x"78"),
  1453 => (x"69",x"64",x"61",x"65"),
  1454 => (x"62",x"20",x"67",x"6e"),
  1455 => (x"20",x"74",x"6f",x"6f"),
  1456 => (x"74",x"63",x"65",x"73"),
  1457 => (x"25",x"20",x"72",x"6f"),
  1458 => (x"52",x"00",x"0a",x"64"),
  1459 => (x"20",x"64",x"61",x"65"),
  1460 => (x"74",x"6f",x"6f",x"62"),
  1461 => (x"63",x"65",x"73",x"20"),
  1462 => (x"20",x"72",x"6f",x"74"),
  1463 => (x"6d",x"6f",x"72",x"66"),
  1464 => (x"72",x"69",x"66",x"20"),
  1465 => (x"70",x"20",x"74",x"73"),
  1466 => (x"69",x"74",x"72",x"61"),
  1467 => (x"6e",x"6f",x"69",x"74"),
  1468 => (x"6e",x"55",x"00",x"0a"),
  1469 => (x"70",x"70",x"75",x"73"),
  1470 => (x"65",x"74",x"72",x"6f"),
  1471 => (x"61",x"70",x"20",x"64"),
  1472 => (x"74",x"69",x"74",x"72"),
  1473 => (x"20",x"6e",x"6f",x"69"),
  1474 => (x"65",x"70",x"79",x"74"),
  1475 => (x"46",x"00",x"0d",x"21"),
  1476 => (x"32",x"33",x"54",x"41"),
  1477 => (x"00",x"20",x"20",x"20"),
  1478 => (x"64",x"61",x"65",x"52"),
  1479 => (x"20",x"67",x"6e",x"69"),
  1480 => (x"0a",x"52",x"42",x"4d"),
  1481 => (x"52",x"42",x"4d",x"00"),
  1482 => (x"63",x"75",x"73",x"20"),
  1483 => (x"73",x"73",x"65",x"63"),
  1484 => (x"6c",x"6c",x"75",x"66"),
  1485 => (x"65",x"72",x"20",x"79"),
  1486 => (x"00",x"0a",x"64",x"61"),
  1487 => (x"31",x"54",x"41",x"46"),
  1488 => (x"20",x"20",x"20",x"36"),
  1489 => (x"54",x"41",x"46",x"00"),
  1490 => (x"20",x"20",x"32",x"33"),
  1491 => (x"61",x"50",x"00",x"20"),
  1492 => (x"74",x"69",x"74",x"72"),
  1493 => (x"63",x"6e",x"6f",x"69"),
  1494 => (x"74",x"6e",x"75",x"6f"),
  1495 => (x"0a",x"64",x"25",x"20"),
  1496 => (x"6e",x"75",x"48",x"00"),
  1497 => (x"67",x"6e",x"69",x"74"),
  1498 => (x"72",x"6f",x"66",x"20"),
  1499 => (x"6c",x"69",x"66",x"20"),
  1500 => (x"73",x"79",x"73",x"65"),
  1501 => (x"0a",x"6d",x"65",x"74"),
  1502 => (x"54",x"41",x"46",x"00"),
  1503 => (x"20",x"20",x"32",x"33"),
  1504 => (x"41",x"46",x"00",x"20"),
  1505 => (x"20",x"36",x"31",x"54"),
  1506 => (x"43",x"00",x"20",x"20"),
  1507 => (x"74",x"73",x"75",x"6c"),
  1508 => (x"73",x"20",x"72",x"65"),
  1509 => (x"3a",x"65",x"7a",x"69"),
  1510 => (x"2c",x"64",x"25",x"20"),
  1511 => (x"75",x"6c",x"43",x"20"),
  1512 => (x"72",x"65",x"74",x"73"),
  1513 => (x"73",x"61",x"6d",x"20"),
  1514 => (x"25",x"20",x"2c",x"6b"),
  1515 => (x"43",x"00",x"0a",x"64"),
  1516 => (x"6b",x"63",x"65",x"68"),
  1517 => (x"6d",x"6d",x"75",x"73"),
  1518 => (x"20",x"67",x"6e",x"69"),
  1519 => (x"6d",x"6f",x"72",x"66"),
  1520 => (x"20",x"64",x"25",x"20"),
  1521 => (x"25",x"20",x"6f",x"74"),
  1522 => (x"2e",x"2e",x"2e",x"64"),
  1523 => (x"64",x"25",x"00",x"20"),
  1524 => (x"64",x"25",x"00",x"0a"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
