
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"d7",x"01"),
     1 => (x"58",x"0e",x"87",x"da"),
     2 => (x"27",x"0e",x"59",x"5e"),
     3 => (x"00",x"00",x"00",x"41"),
     4 => (x"26",x"49",x"26",x"0f"),
     5 => (x"26",x"80",x"ff",x"48"),
     6 => (x"26",x"27",x"4f",x"08"),
     7 => (x"4f",x"00",x"00",x"00"),
     8 => (x"00",x"00",x"33",x"27"),
     9 => (x"c0",x"c2",x"4f",x"00"),
    10 => (x"2d",x"27",x"4e",x"c0"),
    11 => (x"0f",x"00",x"00",x"16"),
    12 => (x"c1",x"87",x"fd",x"00"),
    13 => (x"27",x"4e",x"c0",x"f0"),
    14 => (x"00",x"00",x"00",x"40"),
    15 => (x"87",x"fd",x"00",x"0f"),
    16 => (x"72",x"1e",x"4f",x"4f"),
    17 => (x"c0",x"ff",x"1e",x"1e"),
    18 => (x"c4",x"48",x"6a",x"4a"),
    19 => (x"a6",x"c4",x"98",x"c0"),
    20 => (x"ff",x"02",x"6e",x"58"),
    21 => (x"66",x"cc",x"87",x"f3"),
    22 => (x"48",x"66",x"cc",x"7a"),
    23 => (x"26",x"4a",x"26",x"26"),
    24 => (x"5a",x"5e",x"0e",x"4f"),
    25 => (x"0e",x"5d",x"5c",x"5b"),
    26 => (x"c0",x"4b",x"66",x"d4"),
    27 => (x"74",x"4c",x"13",x"4d"),
    28 => (x"d9",x"c0",x"02",x"9c"),
    29 => (x"c3",x"4a",x"74",x"87"),
    30 => (x"1e",x"72",x"9a",x"ff"),
    31 => (x"00",x"00",x"42",x"27"),
    32 => (x"86",x"c4",x"0f",x"00"),
    33 => (x"4c",x"13",x"85",x"c1"),
    34 => (x"ff",x"05",x"9c",x"74"),
    35 => (x"48",x"75",x"87",x"e7"),
    36 => (x"4c",x"26",x"4d",x"26"),
    37 => (x"4a",x"26",x"4b",x"26"),
    38 => (x"5e",x"0e",x"4f",x"26"),
    39 => (x"5d",x"5c",x"5b",x"5a"),
    40 => (x"c0",x"8e",x"d0",x"0e"),
    41 => (x"49",x"a6",x"c4",x"4c"),
    42 => (x"e8",x"c0",x"79",x"c0"),
    43 => (x"e4",x"c0",x"4b",x"a6"),
    44 => (x"e4",x"c0",x"4a",x"66"),
    45 => (x"80",x"c1",x"48",x"66"),
    46 => (x"58",x"a6",x"e8",x"c0"),
    47 => (x"c0",x"c1",x"48",x"12"),
    48 => (x"90",x"c0",x"c0",x"c0"),
    49 => (x"90",x"b7",x"c0",x"c4"),
    50 => (x"58",x"a6",x"c4",x"48"),
    51 => (x"c0",x"c5",x"02",x"6e"),
    52 => (x"02",x"66",x"c4",x"87"),
    53 => (x"c4",x"87",x"fc",x"c3"),
    54 => (x"79",x"c0",x"49",x"a6"),
    55 => (x"49",x"6e",x"4a",x"6e"),
    56 => (x"02",x"a9",x"f0",x"c0"),
    57 => (x"c1",x"87",x"c2",x"c3"),
    58 => (x"c3",x"02",x"aa",x"e3"),
    59 => (x"e4",x"c1",x"87",x"c3"),
    60 => (x"e3",x"c0",x"02",x"aa"),
    61 => (x"aa",x"ec",x"c1",x"87"),
    62 => (x"87",x"ed",x"c2",x"02"),
    63 => (x"02",x"aa",x"f0",x"c1"),
    64 => (x"c1",x"87",x"d5",x"c0"),
    65 => (x"c2",x"02",x"aa",x"f3"),
    66 => (x"f5",x"c1",x"87",x"c8"),
    67 => (x"c7",x"c0",x"02",x"aa"),
    68 => (x"aa",x"f8",x"c1",x"87"),
    69 => (x"87",x"ee",x"c2",x"05"),
    70 => (x"4a",x"73",x"83",x"c4"),
    71 => (x"49",x"76",x"8a",x"c4"),
    72 => (x"02",x"6e",x"79",x"6a"),
    73 => (x"c8",x"87",x"db",x"c1"),
    74 => (x"79",x"c0",x"49",x"a6"),
    75 => (x"c0",x"49",x"a6",x"cc"),
    76 => (x"dc",x"4a",x"6e",x"79"),
    77 => (x"4d",x"72",x"2a",x"b7"),
    78 => (x"48",x"6e",x"9d",x"cf"),
    79 => (x"a6",x"c4",x"30",x"c4"),
    80 => (x"02",x"9d",x"75",x"58"),
    81 => (x"c8",x"87",x"c5",x"c0"),
    82 => (x"79",x"c1",x"49",x"a6"),
    83 => (x"c0",x"06",x"ad",x"c9"),
    84 => (x"f7",x"c0",x"87",x"c6"),
    85 => (x"87",x"c3",x"c0",x"85"),
    86 => (x"c8",x"85",x"f0",x"c0"),
    87 => (x"cc",x"c0",x"02",x"66"),
    88 => (x"27",x"1e",x"75",x"87"),
    89 => (x"00",x"00",x"00",x"42"),
    90 => (x"c1",x"86",x"c4",x"0f"),
    91 => (x"48",x"66",x"cc",x"84"),
    92 => (x"a6",x"d0",x"80",x"c1"),
    93 => (x"49",x"66",x"cc",x"58"),
    94 => (x"04",x"a9",x"b7",x"c8"),
    95 => (x"c1",x"87",x"f2",x"fe"),
    96 => (x"f0",x"c0",x"87",x"ec"),
    97 => (x"00",x"42",x"27",x"1e"),
    98 => (x"c4",x"0f",x"00",x"00"),
    99 => (x"c1",x"84",x"c1",x"86"),
   100 => (x"83",x"c4",x"87",x"dc"),
   101 => (x"8a",x"c4",x"4a",x"73"),
   102 => (x"61",x"27",x"1e",x"6a"),
   103 => (x"0f",x"00",x"00",x"00"),
   104 => (x"4a",x"70",x"86",x"c4"),
   105 => (x"c5",x"c1",x"84",x"72"),
   106 => (x"49",x"a6",x"c4",x"87"),
   107 => (x"fd",x"c0",x"79",x"c1"),
   108 => (x"73",x"83",x"c4",x"87"),
   109 => (x"6a",x"8a",x"c4",x"4a"),
   110 => (x"00",x"42",x"27",x"1e"),
   111 => (x"c4",x"0f",x"00",x"00"),
   112 => (x"c0",x"84",x"c1",x"86"),
   113 => (x"1e",x"6e",x"87",x"e8"),
   114 => (x"00",x"00",x"42",x"27"),
   115 => (x"86",x"c4",x"0f",x"00"),
   116 => (x"6e",x"87",x"db",x"c0"),
   117 => (x"a9",x"e5",x"c0",x"49"),
   118 => (x"87",x"c8",x"c0",x"05"),
   119 => (x"c1",x"49",x"a6",x"c4"),
   120 => (x"87",x"ca",x"c0",x"79"),
   121 => (x"42",x"27",x"1e",x"6e"),
   122 => (x"0f",x"00",x"00",x"00"),
   123 => (x"e4",x"c0",x"86",x"c4"),
   124 => (x"e4",x"c0",x"4a",x"66"),
   125 => (x"80",x"c1",x"48",x"66"),
   126 => (x"58",x"a6",x"e8",x"c0"),
   127 => (x"c0",x"c1",x"48",x"12"),
   128 => (x"90",x"c0",x"c0",x"c0"),
   129 => (x"90",x"b7",x"c0",x"c4"),
   130 => (x"58",x"a6",x"c4",x"48"),
   131 => (x"c0",x"fb",x"05",x"6e"),
   132 => (x"d0",x"48",x"74",x"87"),
   133 => (x"26",x"4d",x"26",x"86"),
   134 => (x"26",x"4b",x"26",x"4c"),
   135 => (x"00",x"4f",x"26",x"4a"),
   136 => (x"1e",x"00",x"00",x"00"),
   137 => (x"d4",x"ff",x"1e",x"75"),
   138 => (x"49",x"ff",x"c3",x"4d"),
   139 => (x"c8",x"48",x"6d",x"7d"),
   140 => (x"6d",x"7d",x"71",x"38"),
   141 => (x"71",x"38",x"c8",x"b0"),
   142 => (x"c8",x"b0",x"6d",x"7d"),
   143 => (x"6d",x"7d",x"71",x"38"),
   144 => (x"26",x"38",x"c8",x"b0"),
   145 => (x"1e",x"4f",x"26",x"4d"),
   146 => (x"d4",x"ff",x"1e",x"75"),
   147 => (x"49",x"ff",x"c3",x"4d"),
   148 => (x"c8",x"48",x"6d",x"7d"),
   149 => (x"6d",x"7d",x"71",x"30"),
   150 => (x"71",x"30",x"c8",x"b0"),
   151 => (x"c8",x"b0",x"6d",x"7d"),
   152 => (x"6d",x"7d",x"71",x"30"),
   153 => (x"26",x"4d",x"26",x"b0"),
   154 => (x"1e",x"75",x"1e",x"4f"),
   155 => (x"cc",x"4d",x"d4",x"ff"),
   156 => (x"66",x"c8",x"49",x"66"),
   157 => (x"e6",x"fe",x"7d",x"48"),
   158 => (x"31",x"c9",x"02",x"67"),
   159 => (x"09",x"39",x"d8",x"07"),
   160 => (x"09",x"39",x"09",x"7d"),
   161 => (x"09",x"39",x"09",x"7d"),
   162 => (x"09",x"39",x"09",x"7d"),
   163 => (x"70",x"38",x"d0",x"7d"),
   164 => (x"c0",x"f1",x"c9",x"7d"),
   165 => (x"48",x"ff",x"c3",x"49"),
   166 => (x"05",x"a8",x"08",x"6d"),
   167 => (x"7d",x"08",x"87",x"c7"),
   168 => (x"f3",x"05",x"89",x"c1"),
   169 => (x"26",x"4d",x"26",x"87"),
   170 => (x"d4",x"ff",x"1e",x"4f"),
   171 => (x"48",x"c8",x"c3",x"49"),
   172 => (x"05",x"80",x"79",x"ff"),
   173 => (x"4f",x"26",x"87",x"fa"),
   174 => (x"5b",x"5a",x"5e",x"0e"),
   175 => (x"c0",x"0e",x"5d",x"5c"),
   176 => (x"f7",x"c1",x"f0",x"ff"),
   177 => (x"c0",x"c0",x"c1",x"4d"),
   178 => (x"4b",x"c0",x"c0",x"c0"),
   179 => (x"00",x"02",x"a9",x"27"),
   180 => (x"f8",x"c4",x"0f",x"00"),
   181 => (x"1e",x"c0",x"4c",x"df"),
   182 => (x"69",x"27",x"1e",x"75"),
   183 => (x"0f",x"00",x"00",x"02"),
   184 => (x"4a",x"70",x"86",x"c8"),
   185 => (x"05",x"aa",x"b7",x"c1"),
   186 => (x"ff",x"87",x"ef",x"c0"),
   187 => (x"ff",x"c3",x"49",x"d4"),
   188 => (x"c0",x"1e",x"73",x"79"),
   189 => (x"e9",x"c1",x"f0",x"e1"),
   190 => (x"02",x"69",x"27",x"1e"),
   191 => (x"c8",x"0f",x"00",x"00"),
   192 => (x"72",x"4a",x"70",x"86"),
   193 => (x"cb",x"c0",x"05",x"9a"),
   194 => (x"49",x"d4",x"ff",x"87"),
   195 => (x"c1",x"79",x"ff",x"c3"),
   196 => (x"87",x"d0",x"c0",x"48"),
   197 => (x"00",x"02",x"a9",x"27"),
   198 => (x"8c",x"c1",x"0f",x"00"),
   199 => (x"fe",x"05",x"9c",x"74"),
   200 => (x"48",x"c0",x"87",x"f4"),
   201 => (x"4c",x"26",x"4d",x"26"),
   202 => (x"4a",x"26",x"4b",x"26"),
   203 => (x"5e",x"0e",x"4f",x"26"),
   204 => (x"0e",x"5c",x"5b",x"5a"),
   205 => (x"c1",x"f0",x"ff",x"c0"),
   206 => (x"d4",x"ff",x"4c",x"c1"),
   207 => (x"79",x"ff",x"c3",x"49"),
   208 => (x"00",x"17",x"7d",x"27"),
   209 => (x"61",x"27",x"1e",x"00"),
   210 => (x"0f",x"00",x"00",x"00"),
   211 => (x"4b",x"d3",x"86",x"c4"),
   212 => (x"1e",x"74",x"1e",x"c0"),
   213 => (x"00",x"02",x"69",x"27"),
   214 => (x"86",x"c8",x"0f",x"00"),
   215 => (x"9a",x"72",x"4a",x"70"),
   216 => (x"87",x"cb",x"c0",x"05"),
   217 => (x"c3",x"49",x"d4",x"ff"),
   218 => (x"48",x"c1",x"79",x"ff"),
   219 => (x"27",x"87",x"d0",x"c0"),
   220 => (x"00",x"00",x"02",x"a9"),
   221 => (x"73",x"8b",x"c1",x"0f"),
   222 => (x"d3",x"ff",x"05",x"9b"),
   223 => (x"26",x"48",x"c0",x"87"),
   224 => (x"26",x"4b",x"26",x"4c"),
   225 => (x"0e",x"4f",x"26",x"4a"),
   226 => (x"5c",x"5b",x"5a",x"5e"),
   227 => (x"c3",x"1e",x"0e",x"5d"),
   228 => (x"d4",x"ff",x"4d",x"ff"),
   229 => (x"02",x"a9",x"27",x"4c"),
   230 => (x"c6",x"0f",x"00",x"00"),
   231 => (x"e1",x"c0",x"1e",x"ea"),
   232 => (x"1e",x"c8",x"c1",x"f0"),
   233 => (x"00",x"02",x"69",x"27"),
   234 => (x"86",x"c8",x"0f",x"00"),
   235 => (x"1e",x"72",x"4a",x"70"),
   236 => (x"00",x"04",x"e6",x"27"),
   237 => (x"9a",x"27",x"1e",x"00"),
   238 => (x"0f",x"00",x"00",x"00"),
   239 => (x"b7",x"c1",x"86",x"c8"),
   240 => (x"cb",x"c0",x"02",x"aa"),
   241 => (x"03",x"2e",x"27",x"87"),
   242 => (x"c0",x"0f",x"00",x"00"),
   243 => (x"87",x"c9",x"c3",x"48"),
   244 => (x"00",x"02",x"47",x"27"),
   245 => (x"4a",x"70",x"0f",x"00"),
   246 => (x"9a",x"ff",x"ff",x"cf"),
   247 => (x"aa",x"b7",x"ea",x"c6"),
   248 => (x"87",x"cb",x"c0",x"02"),
   249 => (x"00",x"03",x"2e",x"27"),
   250 => (x"48",x"c0",x"0f",x"00"),
   251 => (x"75",x"87",x"ea",x"c2"),
   252 => (x"c0",x"49",x"76",x"7c"),
   253 => (x"b8",x"27",x"79",x"f1"),
   254 => (x"0f",x"00",x"00",x"02"),
   255 => (x"9a",x"72",x"4a",x"70"),
   256 => (x"87",x"eb",x"c1",x"02"),
   257 => (x"ff",x"c0",x"1e",x"c0"),
   258 => (x"1e",x"fa",x"c1",x"f0"),
   259 => (x"00",x"02",x"69",x"27"),
   260 => (x"86",x"c8",x"0f",x"00"),
   261 => (x"9b",x"73",x"4b",x"70"),
   262 => (x"87",x"c3",x"c1",x"05"),
   263 => (x"a4",x"27",x"1e",x"73"),
   264 => (x"1e",x"00",x"00",x"04"),
   265 => (x"00",x"00",x"9a",x"27"),
   266 => (x"86",x"c8",x"0f",x"00"),
   267 => (x"4b",x"6c",x"7c",x"75"),
   268 => (x"1e",x"73",x"9b",x"75"),
   269 => (x"00",x"04",x"b0",x"27"),
   270 => (x"9a",x"27",x"1e",x"00"),
   271 => (x"0f",x"00",x"00",x"00"),
   272 => (x"7c",x"75",x"86",x"c8"),
   273 => (x"7c",x"75",x"7c",x"75"),
   274 => (x"4a",x"73",x"7c",x"75"),
   275 => (x"72",x"9a",x"c0",x"c1"),
   276 => (x"c5",x"c0",x"02",x"9a"),
   277 => (x"c0",x"48",x"c1",x"87"),
   278 => (x"48",x"c0",x"87",x"ff"),
   279 => (x"73",x"87",x"fa",x"c0"),
   280 => (x"04",x"be",x"27",x"1e"),
   281 => (x"27",x"1e",x"00",x"00"),
   282 => (x"00",x"00",x"00",x"9a"),
   283 => (x"6e",x"86",x"c8",x"0f"),
   284 => (x"a9",x"b7",x"c2",x"49"),
   285 => (x"87",x"d3",x"c0",x"05"),
   286 => (x"00",x"04",x"ca",x"27"),
   287 => (x"9a",x"27",x"1e",x"00"),
   288 => (x"0f",x"00",x"00",x"00"),
   289 => (x"48",x"c0",x"86",x"c4"),
   290 => (x"6e",x"87",x"ce",x"c0"),
   291 => (x"c4",x"88",x"c1",x"48"),
   292 => (x"05",x"6e",x"58",x"a6"),
   293 => (x"c0",x"87",x"df",x"fd"),
   294 => (x"4d",x"26",x"26",x"48"),
   295 => (x"4b",x"26",x"4c",x"26"),
   296 => (x"4f",x"26",x"4a",x"26"),
   297 => (x"35",x"44",x"4d",x"43"),
   298 => (x"64",x"25",x"20",x"38"),
   299 => (x"00",x"20",x"20",x"0a"),
   300 => (x"35",x"44",x"4d",x"43"),
   301 => (x"20",x"32",x"5f",x"38"),
   302 => (x"20",x"0a",x"64",x"25"),
   303 => (x"4d",x"43",x"00",x"20"),
   304 => (x"20",x"38",x"35",x"44"),
   305 => (x"20",x"0a",x"64",x"25"),
   306 => (x"44",x"53",x"00",x"20"),
   307 => (x"49",x"20",x"43",x"48"),
   308 => (x"69",x"74",x"69",x"6e"),
   309 => (x"7a",x"69",x"6c",x"61"),
   310 => (x"6f",x"69",x"74",x"61"),
   311 => (x"72",x"65",x"20",x"6e"),
   312 => (x"21",x"72",x"6f",x"72"),
   313 => (x"6d",x"63",x"00",x"0a"),
   314 => (x"4d",x"43",x"5f",x"64"),
   315 => (x"72",x"20",x"38",x"44"),
   316 => (x"6f",x"70",x"73",x"65"),
   317 => (x"3a",x"65",x"73",x"6e"),
   318 => (x"0a",x"64",x"25",x"20"),
   319 => (x"5a",x"5e",x"0e",x"00"),
   320 => (x"0e",x"5d",x"5c",x"5b"),
   321 => (x"4c",x"d0",x"ff",x"1e"),
   322 => (x"4b",x"c0",x"c0",x"c8"),
   323 => (x"00",x"02",x"1f",x"27"),
   324 => (x"79",x"c1",x"49",x"00"),
   325 => (x"00",x"06",x"1a",x"27"),
   326 => (x"61",x"27",x"1e",x"00"),
   327 => (x"0f",x"00",x"00",x"00"),
   328 => (x"4d",x"c7",x"86",x"c4"),
   329 => (x"98",x"73",x"48",x"6c"),
   330 => (x"6e",x"58",x"a6",x"c4"),
   331 => (x"87",x"cc",x"c0",x"02"),
   332 => (x"98",x"73",x"48",x"6c"),
   333 => (x"6e",x"58",x"a6",x"c4"),
   334 => (x"87",x"f4",x"ff",x"05"),
   335 => (x"a9",x"27",x"7c",x"c0"),
   336 => (x"0f",x"00",x"00",x"02"),
   337 => (x"98",x"73",x"48",x"6c"),
   338 => (x"6e",x"58",x"a6",x"c4"),
   339 => (x"87",x"cc",x"c0",x"02"),
   340 => (x"98",x"73",x"48",x"6c"),
   341 => (x"6e",x"58",x"a6",x"c4"),
   342 => (x"87",x"f4",x"ff",x"05"),
   343 => (x"1e",x"c0",x"7c",x"c1"),
   344 => (x"c1",x"d0",x"e5",x"c0"),
   345 => (x"69",x"27",x"1e",x"c0"),
   346 => (x"0f",x"00",x"00",x"02"),
   347 => (x"4a",x"70",x"86",x"c8"),
   348 => (x"05",x"aa",x"b7",x"c1"),
   349 => (x"c1",x"87",x"c2",x"c0"),
   350 => (x"ad",x"b7",x"c2",x"4d"),
   351 => (x"87",x"d3",x"c0",x"05"),
   352 => (x"00",x"06",x"15",x"27"),
   353 => (x"61",x"27",x"1e",x"00"),
   354 => (x"0f",x"00",x"00",x"00"),
   355 => (x"48",x"c0",x"86",x"c4"),
   356 => (x"c1",x"87",x"f7",x"c1"),
   357 => (x"05",x"9d",x"75",x"8d"),
   358 => (x"27",x"87",x"c9",x"fe"),
   359 => (x"00",x"00",x"03",x"87"),
   360 => (x"02",x"23",x"27",x"0f"),
   361 => (x"27",x"58",x"00",x"00"),
   362 => (x"00",x"00",x"02",x"1f"),
   363 => (x"d0",x"c0",x"05",x"bf"),
   364 => (x"c0",x"1e",x"c1",x"87"),
   365 => (x"d0",x"c1",x"f0",x"ff"),
   366 => (x"02",x"69",x"27",x"1e"),
   367 => (x"c8",x"0f",x"00",x"00"),
   368 => (x"49",x"d4",x"ff",x"86"),
   369 => (x"27",x"79",x"ff",x"c3"),
   370 => (x"00",x"00",x"08",x"b0"),
   371 => (x"19",x"18",x"27",x"0f"),
   372 => (x"27",x"58",x"00",x"00"),
   373 => (x"00",x"00",x"19",x"14"),
   374 => (x"1e",x"27",x"1e",x"bf"),
   375 => (x"1e",x"00",x"00",x"06"),
   376 => (x"00",x"00",x"9a",x"27"),
   377 => (x"86",x"c8",x"0f",x"00"),
   378 => (x"98",x"73",x"48",x"6c"),
   379 => (x"6e",x"58",x"a6",x"c4"),
   380 => (x"87",x"cc",x"c0",x"02"),
   381 => (x"98",x"73",x"48",x"6c"),
   382 => (x"6e",x"58",x"a6",x"c4"),
   383 => (x"87",x"f4",x"ff",x"05"),
   384 => (x"d4",x"ff",x"7c",x"c0"),
   385 => (x"79",x"ff",x"c3",x"49"),
   386 => (x"26",x"26",x"48",x"c1"),
   387 => (x"26",x"4c",x"26",x"4d"),
   388 => (x"26",x"4a",x"26",x"4b"),
   389 => (x"52",x"45",x"49",x"4f"),
   390 => (x"50",x"53",x"00",x"52"),
   391 => (x"44",x"53",x"00",x"49"),
   392 => (x"72",x"61",x"63",x"20"),
   393 => (x"69",x"73",x"20",x"64"),
   394 => (x"69",x"20",x"65",x"7a"),
   395 => (x"64",x"25",x"20",x"73"),
   396 => (x"5e",x"0e",x"00",x"0a"),
   397 => (x"5d",x"5c",x"5b",x"5a"),
   398 => (x"ff",x"c3",x"1e",x"0e"),
   399 => (x"4c",x"d4",x"ff",x"4d"),
   400 => (x"d0",x"ff",x"7c",x"75"),
   401 => (x"c0",x"c8",x"48",x"bf"),
   402 => (x"a6",x"c4",x"98",x"c0"),
   403 => (x"c0",x"02",x"6e",x"58"),
   404 => (x"c0",x"c8",x"87",x"d2"),
   405 => (x"d0",x"ff",x"4a",x"c0"),
   406 => (x"98",x"72",x"48",x"bf"),
   407 => (x"6e",x"58",x"a6",x"c4"),
   408 => (x"87",x"f2",x"ff",x"05"),
   409 => (x"c4",x"49",x"d0",x"ff"),
   410 => (x"7c",x"75",x"79",x"c1"),
   411 => (x"c0",x"1e",x"66",x"d8"),
   412 => (x"d8",x"c1",x"f0",x"ff"),
   413 => (x"02",x"69",x"27",x"1e"),
   414 => (x"c8",x"0f",x"00",x"00"),
   415 => (x"72",x"4a",x"70",x"86"),
   416 => (x"d3",x"c0",x"02",x"9a"),
   417 => (x"07",x"3a",x"27",x"87"),
   418 => (x"27",x"1e",x"00",x"00"),
   419 => (x"00",x"00",x"00",x"61"),
   420 => (x"c1",x"86",x"c4",x"0f"),
   421 => (x"87",x"d7",x"c2",x"48"),
   422 => (x"fe",x"c3",x"7c",x"75"),
   423 => (x"c0",x"49",x"76",x"7c"),
   424 => (x"bf",x"66",x"dc",x"79"),
   425 => (x"d8",x"4b",x"72",x"4a"),
   426 => (x"48",x"73",x"2b",x"b7"),
   427 => (x"7c",x"70",x"98",x"75"),
   428 => (x"b7",x"d0",x"4b",x"72"),
   429 => (x"75",x"48",x"73",x"2b"),
   430 => (x"72",x"7c",x"70",x"98"),
   431 => (x"2b",x"b7",x"c8",x"4b"),
   432 => (x"98",x"75",x"48",x"73"),
   433 => (x"48",x"72",x"7c",x"70"),
   434 => (x"7c",x"70",x"98",x"75"),
   435 => (x"c4",x"48",x"66",x"dc"),
   436 => (x"a6",x"e0",x"c0",x"80"),
   437 => (x"c1",x"48",x"6e",x"58"),
   438 => (x"58",x"a6",x"c4",x"80"),
   439 => (x"c0",x"c2",x"49",x"6e"),
   440 => (x"fe",x"04",x"a9",x"b7"),
   441 => (x"7c",x"75",x"87",x"fb"),
   442 => (x"7c",x"75",x"7c",x"75"),
   443 => (x"4b",x"e0",x"da",x"d8"),
   444 => (x"4a",x"6c",x"7c",x"75"),
   445 => (x"9a",x"72",x"9a",x"75"),
   446 => (x"87",x"c8",x"c0",x"05"),
   447 => (x"9b",x"73",x"8b",x"c1"),
   448 => (x"87",x"ec",x"ff",x"05"),
   449 => (x"d0",x"ff",x"7c",x"75"),
   450 => (x"c0",x"c8",x"48",x"bf"),
   451 => (x"a6",x"c4",x"98",x"c0"),
   452 => (x"c0",x"02",x"6e",x"58"),
   453 => (x"c0",x"c8",x"87",x"d2"),
   454 => (x"d0",x"ff",x"4a",x"c0"),
   455 => (x"98",x"72",x"48",x"bf"),
   456 => (x"6e",x"58",x"a6",x"c4"),
   457 => (x"87",x"f2",x"ff",x"05"),
   458 => (x"c0",x"49",x"d0",x"ff"),
   459 => (x"26",x"48",x"c0",x"79"),
   460 => (x"4c",x"26",x"4d",x"26"),
   461 => (x"4a",x"26",x"4b",x"26"),
   462 => (x"72",x"57",x"4f",x"26"),
   463 => (x"20",x"65",x"74",x"69"),
   464 => (x"6c",x"69",x"61",x"66"),
   465 => (x"00",x"0a",x"64",x"65"),
   466 => (x"5b",x"5a",x"5e",x"0e"),
   467 => (x"1e",x"0e",x"5d",x"5c"),
   468 => (x"dc",x"4c",x"66",x"d8"),
   469 => (x"49",x"76",x"4b",x"66"),
   470 => (x"ee",x"c5",x"79",x"c0"),
   471 => (x"ff",x"4d",x"df",x"cd"),
   472 => (x"ff",x"c3",x"49",x"d4"),
   473 => (x"bf",x"d4",x"ff",x"79"),
   474 => (x"9a",x"ff",x"c3",x"4a"),
   475 => (x"aa",x"b7",x"fe",x"c3"),
   476 => (x"87",x"e5",x"c1",x"05"),
   477 => (x"00",x"19",x"10",x"27"),
   478 => (x"79",x"c0",x"49",x"00"),
   479 => (x"04",x"ab",x"b7",x"c4"),
   480 => (x"27",x"87",x"e4",x"c0"),
   481 => (x"00",x"00",x"02",x"23"),
   482 => (x"72",x"4a",x"70",x"0f"),
   483 => (x"27",x"84",x"c4",x"7c"),
   484 => (x"00",x"00",x"19",x"10"),
   485 => (x"80",x"72",x"48",x"bf"),
   486 => (x"00",x"19",x"14",x"27"),
   487 => (x"8b",x"c4",x"58",x"00"),
   488 => (x"03",x"ab",x"b7",x"c4"),
   489 => (x"c0",x"87",x"dc",x"ff"),
   490 => (x"c0",x"06",x"ab",x"b7"),
   491 => (x"d4",x"ff",x"87",x"e5"),
   492 => (x"7d",x"ff",x"c3",x"4d"),
   493 => (x"97",x"72",x"4a",x"6d"),
   494 => (x"27",x"84",x"c1",x"7c"),
   495 => (x"00",x"00",x"19",x"10"),
   496 => (x"80",x"72",x"48",x"bf"),
   497 => (x"00",x"19",x"14",x"27"),
   498 => (x"8b",x"c1",x"58",x"00"),
   499 => (x"01",x"ab",x"b7",x"c0"),
   500 => (x"c1",x"87",x"de",x"ff"),
   501 => (x"c1",x"49",x"76",x"4d"),
   502 => (x"75",x"8d",x"c1",x"79"),
   503 => (x"fe",x"fd",x"05",x"9d"),
   504 => (x"49",x"d4",x"ff",x"87"),
   505 => (x"6e",x"79",x"ff",x"c3"),
   506 => (x"4d",x"26",x"26",x"48"),
   507 => (x"4b",x"26",x"4c",x"26"),
   508 => (x"4f",x"26",x"4a",x"26"),
   509 => (x"5b",x"5a",x"5e",x"0e"),
   510 => (x"1e",x"0e",x"5d",x"5c"),
   511 => (x"c8",x"4b",x"d0",x"ff"),
   512 => (x"c0",x"4a",x"c0",x"c0"),
   513 => (x"49",x"d4",x"ff",x"4c"),
   514 => (x"6b",x"79",x"ff",x"c3"),
   515 => (x"c4",x"98",x"72",x"48"),
   516 => (x"02",x"6e",x"58",x"a6"),
   517 => (x"6b",x"87",x"cc",x"c0"),
   518 => (x"c4",x"98",x"72",x"48"),
   519 => (x"05",x"6e",x"58",x"a6"),
   520 => (x"c4",x"87",x"f4",x"ff"),
   521 => (x"d4",x"ff",x"7b",x"c1"),
   522 => (x"79",x"ff",x"c3",x"49"),
   523 => (x"c0",x"1e",x"66",x"d8"),
   524 => (x"d1",x"c1",x"f0",x"ff"),
   525 => (x"02",x"69",x"27",x"1e"),
   526 => (x"c8",x"0f",x"00",x"00"),
   527 => (x"75",x"4d",x"70",x"86"),
   528 => (x"d6",x"c0",x"02",x"9d"),
   529 => (x"dc",x"1e",x"75",x"87"),
   530 => (x"90",x"27",x"1e",x"66"),
   531 => (x"1e",x"00",x"00",x"08"),
   532 => (x"00",x"00",x"9a",x"27"),
   533 => (x"86",x"cc",x"0f",x"00"),
   534 => (x"c8",x"87",x"e8",x"c0"),
   535 => (x"e0",x"c0",x"1e",x"c0"),
   536 => (x"e3",x"fb",x"1e",x"66"),
   537 => (x"70",x"86",x"c8",x"87"),
   538 => (x"72",x"48",x"6b",x"4c"),
   539 => (x"58",x"a6",x"c4",x"98"),
   540 => (x"cc",x"c0",x"02",x"6e"),
   541 => (x"72",x"48",x"6b",x"87"),
   542 => (x"58",x"a6",x"c4",x"98"),
   543 => (x"f4",x"ff",x"05",x"6e"),
   544 => (x"74",x"7b",x"c0",x"87"),
   545 => (x"4d",x"26",x"26",x"48"),
   546 => (x"4b",x"26",x"4c",x"26"),
   547 => (x"4f",x"26",x"4a",x"26"),
   548 => (x"64",x"61",x"65",x"52"),
   549 => (x"6d",x"6f",x"63",x"20"),
   550 => (x"64",x"6e",x"61",x"6d"),
   551 => (x"69",x"61",x"66",x"20"),
   552 => (x"20",x"64",x"65",x"6c"),
   553 => (x"25",x"20",x"74",x"61"),
   554 => (x"25",x"28",x"20",x"64"),
   555 => (x"00",x"0a",x"29",x"64"),
   556 => (x"5b",x"5a",x"5e",x"0e"),
   557 => (x"1e",x"0e",x"5d",x"5c"),
   558 => (x"ff",x"c0",x"1e",x"c0"),
   559 => (x"1e",x"c9",x"c1",x"f0"),
   560 => (x"00",x"02",x"69",x"27"),
   561 => (x"86",x"c8",x"0f",x"00"),
   562 => (x"20",x"27",x"1e",x"d2"),
   563 => (x"1e",x"00",x"00",x"19"),
   564 => (x"c8",x"87",x"f5",x"f9"),
   565 => (x"c1",x"4d",x"c0",x"86"),
   566 => (x"ad",x"b7",x"d2",x"85"),
   567 => (x"87",x"f7",x"ff",x"04"),
   568 => (x"00",x"19",x"20",x"27"),
   569 => (x"4a",x"bf",x"97",x"00"),
   570 => (x"c1",x"9a",x"c0",x"c3"),
   571 => (x"05",x"aa",x"b7",x"c0"),
   572 => (x"27",x"87",x"f2",x"c0"),
   573 => (x"00",x"00",x"19",x"27"),
   574 => (x"d0",x"4a",x"bf",x"97"),
   575 => (x"19",x"28",x"27",x"32"),
   576 => (x"bf",x"97",x"00",x"00"),
   577 => (x"72",x"33",x"c8",x"4b"),
   578 => (x"27",x"b2",x"73",x"4a"),
   579 => (x"00",x"00",x"19",x"29"),
   580 => (x"72",x"4b",x"bf",x"97"),
   581 => (x"cf",x"b2",x"73",x"4a"),
   582 => (x"9a",x"ff",x"ff",x"ff"),
   583 => (x"85",x"c1",x"4d",x"72"),
   584 => (x"cb",x"c3",x"35",x"ca"),
   585 => (x"19",x"29",x"27",x"87"),
   586 => (x"bf",x"97",x"00",x"00"),
   587 => (x"c6",x"32",x"c1",x"4a"),
   588 => (x"19",x"2a",x"27",x"9a"),
   589 => (x"bf",x"97",x"00",x"00"),
   590 => (x"2b",x"b7",x"c7",x"4b"),
   591 => (x"b2",x"73",x"4a",x"72"),
   592 => (x"00",x"19",x"25",x"27"),
   593 => (x"4b",x"bf",x"97",x"00"),
   594 => (x"98",x"cf",x"48",x"73"),
   595 => (x"27",x"58",x"a6",x"c4"),
   596 => (x"00",x"00",x"19",x"26"),
   597 => (x"c3",x"4b",x"bf",x"97"),
   598 => (x"27",x"33",x"ca",x"9b"),
   599 => (x"00",x"00",x"19",x"27"),
   600 => (x"c2",x"4c",x"bf",x"97"),
   601 => (x"74",x"4b",x"73",x"34"),
   602 => (x"19",x"28",x"27",x"b3"),
   603 => (x"bf",x"97",x"00",x"00"),
   604 => (x"9c",x"c0",x"c3",x"4c"),
   605 => (x"73",x"2c",x"b7",x"c6"),
   606 => (x"73",x"b3",x"74",x"4b"),
   607 => (x"1e",x"66",x"c4",x"1e"),
   608 => (x"fd",x"27",x"1e",x"72"),
   609 => (x"1e",x"00",x"00",x"09"),
   610 => (x"00",x"00",x"9a",x"27"),
   611 => (x"86",x"d0",x"0f",x"00"),
   612 => (x"48",x"c1",x"82",x"c2"),
   613 => (x"4a",x"70",x"30",x"72"),
   614 => (x"2a",x"27",x"1e",x"72"),
   615 => (x"1e",x"00",x"00",x"0a"),
   616 => (x"00",x"00",x"9a",x"27"),
   617 => (x"86",x"c8",x"0f",x"00"),
   618 => (x"30",x"6e",x"48",x"c1"),
   619 => (x"c1",x"58",x"a6",x"c4"),
   620 => (x"72",x"4d",x"73",x"83"),
   621 => (x"75",x"1e",x"6e",x"95"),
   622 => (x"0a",x"33",x"27",x"1e"),
   623 => (x"27",x"1e",x"00",x"00"),
   624 => (x"00",x"00",x"00",x"9a"),
   625 => (x"6e",x"86",x"cc",x"0f"),
   626 => (x"b7",x"c0",x"c8",x"49"),
   627 => (x"cf",x"c0",x"06",x"a9"),
   628 => (x"c1",x"4a",x"6e",x"87"),
   629 => (x"2a",x"b7",x"c1",x"35"),
   630 => (x"aa",x"b7",x"c0",x"c8"),
   631 => (x"87",x"f3",x"ff",x"01"),
   632 => (x"49",x"27",x"1e",x"75"),
   633 => (x"1e",x"00",x"00",x"0a"),
   634 => (x"00",x"00",x"9a",x"27"),
   635 => (x"86",x"c8",x"0f",x"00"),
   636 => (x"26",x"26",x"48",x"75"),
   637 => (x"26",x"4c",x"26",x"4d"),
   638 => (x"26",x"4a",x"26",x"4b"),
   639 => (x"73",x"5f",x"63",x"4f"),
   640 => (x"5f",x"65",x"7a",x"69"),
   641 => (x"74",x"6c",x"75",x"6d"),
   642 => (x"64",x"25",x"20",x"3a"),
   643 => (x"65",x"72",x"20",x"2c"),
   644 => (x"62",x"5f",x"64",x"61"),
   645 => (x"65",x"6c",x"5f",x"6c"),
   646 => (x"25",x"20",x"3a",x"6e"),
   647 => (x"63",x"20",x"2c",x"64"),
   648 => (x"65",x"7a",x"69",x"73"),
   649 => (x"64",x"25",x"20",x"3a"),
   650 => (x"75",x"4d",x"00",x"0a"),
   651 => (x"25",x"20",x"74",x"6c"),
   652 => (x"25",x"00",x"0a",x"64"),
   653 => (x"6c",x"62",x"20",x"64"),
   654 => (x"73",x"6b",x"63",x"6f"),
   655 => (x"20",x"66",x"6f",x"20"),
   656 => (x"65",x"7a",x"69",x"73"),
   657 => (x"0a",x"64",x"25",x"20"),
   658 => (x"20",x"64",x"25",x"00"),
   659 => (x"63",x"6f",x"6c",x"62"),
   660 => (x"6f",x"20",x"73",x"6b"),
   661 => (x"31",x"35",x"20",x"66"),
   662 => (x"79",x"62",x"20",x"32"),
   663 => (x"0a",x"73",x"65",x"74"),
   664 => (x"5a",x"5e",x"0e",x"00"),
   665 => (x"0e",x"5d",x"5c",x"5b"),
   666 => (x"c0",x"4d",x"66",x"d4"),
   667 => (x"49",x"66",x"dc",x"4c"),
   668 => (x"06",x"a9",x"b7",x"c0"),
   669 => (x"15",x"87",x"fb",x"c0"),
   670 => (x"c0",x"c0",x"c1",x"4b"),
   671 => (x"c4",x"93",x"c0",x"c0"),
   672 => (x"4b",x"93",x"b7",x"c0"),
   673 => (x"bf",x"97",x"66",x"d8"),
   674 => (x"c0",x"c0",x"c1",x"4a"),
   675 => (x"c4",x"92",x"c0",x"c0"),
   676 => (x"4a",x"92",x"b7",x"c0"),
   677 => (x"c1",x"48",x"66",x"d8"),
   678 => (x"58",x"a6",x"dc",x"80"),
   679 => (x"02",x"ab",x"b7",x"72"),
   680 => (x"c1",x"87",x"c5",x"c0"),
   681 => (x"87",x"cc",x"c0",x"48"),
   682 => (x"66",x"dc",x"84",x"c1"),
   683 => (x"ff",x"04",x"ac",x"b7"),
   684 => (x"48",x"c0",x"87",x"c5"),
   685 => (x"4c",x"26",x"4d",x"26"),
   686 => (x"4a",x"26",x"4b",x"26"),
   687 => (x"5e",x"0e",x"4f",x"26"),
   688 => (x"5d",x"5c",x"5b",x"5a"),
   689 => (x"1b",x"40",x"27",x"0e"),
   690 => (x"c0",x"49",x"00",x"00"),
   691 => (x"18",x"55",x"27",x"79"),
   692 => (x"27",x"1e",x"00",x"00"),
   693 => (x"00",x"00",x"00",x"61"),
   694 => (x"27",x"86",x"c4",x"0f"),
   695 => (x"00",x"00",x"19",x"38"),
   696 => (x"27",x"1e",x"c0",x"1e"),
   697 => (x"00",x"00",x"07",x"f4"),
   698 => (x"70",x"86",x"c8",x"0f"),
   699 => (x"05",x"9a",x"72",x"4a"),
   700 => (x"27",x"87",x"d3",x"c0"),
   701 => (x"00",x"00",x"17",x"81"),
   702 => (x"00",x"61",x"27",x"1e"),
   703 => (x"c4",x"0f",x"00",x"00"),
   704 => (x"d0",x"48",x"c0",x"86"),
   705 => (x"62",x"27",x"87",x"c5"),
   706 => (x"1e",x"00",x"00",x"18"),
   707 => (x"00",x"00",x"61",x"27"),
   708 => (x"86",x"c4",x"0f",x"00"),
   709 => (x"6c",x"27",x"4c",x"c0"),
   710 => (x"49",x"00",x"00",x"1b"),
   711 => (x"1e",x"c8",x"79",x"c1"),
   712 => (x"00",x"18",x"79",x"27"),
   713 => (x"6e",x"27",x"1e",x"00"),
   714 => (x"1e",x"00",x"00",x"19"),
   715 => (x"00",x"0a",x"61",x"27"),
   716 => (x"86",x"cc",x"0f",x"00"),
   717 => (x"9a",x"72",x"4a",x"70"),
   718 => (x"87",x"c8",x"c0",x"05"),
   719 => (x"00",x"1b",x"6c",x"27"),
   720 => (x"79",x"c0",x"49",x"00"),
   721 => (x"82",x"27",x"1e",x"c8"),
   722 => (x"1e",x"00",x"00",x"18"),
   723 => (x"00",x"19",x"8a",x"27"),
   724 => (x"61",x"27",x"1e",x"00"),
   725 => (x"0f",x"00",x"00",x"0a"),
   726 => (x"4a",x"70",x"86",x"cc"),
   727 => (x"c0",x"05",x"9a",x"72"),
   728 => (x"6c",x"27",x"87",x"c8"),
   729 => (x"49",x"00",x"00",x"1b"),
   730 => (x"6c",x"27",x"79",x"c0"),
   731 => (x"bf",x"00",x"00",x"1b"),
   732 => (x"18",x"8b",x"27",x"1e"),
   733 => (x"27",x"1e",x"00",x"00"),
   734 => (x"00",x"00",x"00",x"9a"),
   735 => (x"27",x"86",x"c8",x"0f"),
   736 => (x"00",x"00",x"1b",x"6c"),
   737 => (x"ca",x"c3",x"02",x"bf"),
   738 => (x"19",x"38",x"27",x"87"),
   739 => (x"27",x"4d",x"00",x"00"),
   740 => (x"00",x"00",x"1a",x"f6"),
   741 => (x"1b",x"36",x"27",x"4b"),
   742 => (x"bf",x"9f",x"00",x"00"),
   743 => (x"ff",x"ff",x"cf",x"4a"),
   744 => (x"27",x"1e",x"72",x"9a"),
   745 => (x"00",x"00",x"1b",x"36"),
   746 => (x"19",x"38",x"27",x"4a"),
   747 => (x"72",x"8a",x"00",x"00"),
   748 => (x"c8",x"1e",x"d0",x"1e"),
   749 => (x"b3",x"27",x"1e",x"c0"),
   750 => (x"1e",x"00",x"00",x"17"),
   751 => (x"00",x"00",x"9a",x"27"),
   752 => (x"86",x"d4",x"0f",x"00"),
   753 => (x"82",x"c8",x"4a",x"73"),
   754 => (x"36",x"27",x"4c",x"6a"),
   755 => (x"9f",x"00",x"00",x"1b"),
   756 => (x"ff",x"cf",x"4a",x"bf"),
   757 => (x"d6",x"c5",x"9a",x"ff"),
   758 => (x"c0",x"05",x"aa",x"ea"),
   759 => (x"4a",x"73",x"87",x"d3"),
   760 => (x"1e",x"6a",x"82",x"c8"),
   761 => (x"00",x"12",x"7c",x"27"),
   762 => (x"86",x"c4",x"0f",x"00"),
   763 => (x"e7",x"c0",x"4c",x"70"),
   764 => (x"c7",x"4a",x"75",x"87"),
   765 => (x"6a",x"9f",x"82",x"fe"),
   766 => (x"ff",x"ff",x"cf",x"4a"),
   767 => (x"d5",x"e9",x"ca",x"9a"),
   768 => (x"d3",x"c0",x"02",x"aa"),
   769 => (x"17",x"95",x"27",x"87"),
   770 => (x"27",x"1e",x"00",x"00"),
   771 => (x"00",x"00",x"00",x"61"),
   772 => (x"c0",x"86",x"c4",x"0f"),
   773 => (x"87",x"f3",x"cb",x"48"),
   774 => (x"f0",x"27",x"1e",x"74"),
   775 => (x"1e",x"00",x"00",x"17"),
   776 => (x"00",x"00",x"9a",x"27"),
   777 => (x"86",x"c8",x"0f",x"00"),
   778 => (x"00",x"19",x"38",x"27"),
   779 => (x"1e",x"74",x"1e",x"00"),
   780 => (x"00",x"07",x"f4",x"27"),
   781 => (x"86",x"c8",x"0f",x"00"),
   782 => (x"9a",x"72",x"4a",x"70"),
   783 => (x"87",x"c5",x"c0",x"05"),
   784 => (x"c6",x"cb",x"48",x"c0"),
   785 => (x"18",x"08",x"27",x"87"),
   786 => (x"27",x"1e",x"00",x"00"),
   787 => (x"00",x"00",x"00",x"61"),
   788 => (x"27",x"86",x"c4",x"0f"),
   789 => (x"00",x"00",x"18",x"9e"),
   790 => (x"00",x"9a",x"27",x"1e"),
   791 => (x"c4",x"0f",x"00",x"00"),
   792 => (x"27",x"1e",x"c8",x"86"),
   793 => (x"00",x"00",x"18",x"b6"),
   794 => (x"19",x"8a",x"27",x"1e"),
   795 => (x"27",x"1e",x"00",x"00"),
   796 => (x"00",x"00",x"0a",x"61"),
   797 => (x"70",x"86",x"cc",x"0f"),
   798 => (x"05",x"9a",x"72",x"4a"),
   799 => (x"27",x"87",x"cb",x"c0"),
   800 => (x"00",x"00",x"1b",x"40"),
   801 => (x"c0",x"79",x"c1",x"49"),
   802 => (x"1e",x"c8",x"87",x"f1"),
   803 => (x"00",x"18",x"bf",x"27"),
   804 => (x"6e",x"27",x"1e",x"00"),
   805 => (x"1e",x"00",x"00",x"19"),
   806 => (x"00",x"0a",x"61",x"27"),
   807 => (x"86",x"cc",x"0f",x"00"),
   808 => (x"9a",x"72",x"4a",x"70"),
   809 => (x"87",x"d3",x"c0",x"02"),
   810 => (x"00",x"18",x"2f",x"27"),
   811 => (x"9a",x"27",x"1e",x"00"),
   812 => (x"0f",x"00",x"00",x"00"),
   813 => (x"48",x"c0",x"86",x"c4"),
   814 => (x"27",x"87",x"d0",x"c9"),
   815 => (x"00",x"00",x"1b",x"36"),
   816 => (x"c3",x"4a",x"bf",x"97"),
   817 => (x"d5",x"c1",x"9a",x"ff"),
   818 => (x"d2",x"c0",x"05",x"aa"),
   819 => (x"1b",x"37",x"27",x"87"),
   820 => (x"bf",x"97",x"00",x"00"),
   821 => (x"9a",x"ff",x"c3",x"4a"),
   822 => (x"02",x"aa",x"ea",x"c2"),
   823 => (x"c0",x"87",x"c5",x"c0"),
   824 => (x"87",x"e7",x"c8",x"48"),
   825 => (x"00",x"19",x"38",x"27"),
   826 => (x"4a",x"bf",x"97",x"00"),
   827 => (x"c3",x"9a",x"ff",x"c3"),
   828 => (x"c0",x"02",x"aa",x"e9"),
   829 => (x"38",x"27",x"87",x"d7"),
   830 => (x"97",x"00",x"00",x"19"),
   831 => (x"ff",x"c3",x"4a",x"bf"),
   832 => (x"aa",x"eb",x"c3",x"9a"),
   833 => (x"87",x"c5",x"c0",x"02"),
   834 => (x"fe",x"c7",x"48",x"c0"),
   835 => (x"19",x"43",x"27",x"87"),
   836 => (x"bf",x"97",x"00",x"00"),
   837 => (x"9a",x"ff",x"c3",x"4a"),
   838 => (x"c0",x"05",x"9a",x"72"),
   839 => (x"44",x"27",x"87",x"d1"),
   840 => (x"97",x"00",x"00",x"19"),
   841 => (x"ff",x"c3",x"4a",x"bf"),
   842 => (x"02",x"aa",x"c2",x"9a"),
   843 => (x"c0",x"87",x"c5",x"c0"),
   844 => (x"87",x"d7",x"c7",x"48"),
   845 => (x"00",x"19",x"45",x"27"),
   846 => (x"48",x"bf",x"97",x"00"),
   847 => (x"27",x"98",x"ff",x"c3"),
   848 => (x"00",x"00",x"1b",x"3c"),
   849 => (x"1b",x"38",x"27",x"58"),
   850 => (x"4a",x"bf",x"00",x"00"),
   851 => (x"8b",x"c1",x"4b",x"72"),
   852 => (x"00",x"1b",x"3c",x"27"),
   853 => (x"79",x"73",x"49",x"00"),
   854 => (x"1e",x"72",x"1e",x"73"),
   855 => (x"00",x"18",x"c8",x"27"),
   856 => (x"9a",x"27",x"1e",x"00"),
   857 => (x"0f",x"00",x"00",x"00"),
   858 => (x"46",x"27",x"86",x"cc"),
   859 => (x"97",x"00",x"00",x"19"),
   860 => (x"ff",x"c3",x"4a",x"bf"),
   861 => (x"27",x"82",x"74",x"9a"),
   862 => (x"00",x"00",x"19",x"47"),
   863 => (x"c3",x"4b",x"bf",x"97"),
   864 => (x"33",x"c8",x"9b",x"ff"),
   865 => (x"80",x"72",x"48",x"73"),
   866 => (x"00",x"1b",x"50",x"27"),
   867 => (x"48",x"27",x"58",x"00"),
   868 => (x"97",x"00",x"00",x"19"),
   869 => (x"ff",x"c3",x"48",x"bf"),
   870 => (x"1b",x"64",x"27",x"98"),
   871 => (x"27",x"58",x"00",x"00"),
   872 => (x"00",x"00",x"1b",x"40"),
   873 => (x"e5",x"c3",x"02",x"bf"),
   874 => (x"27",x"1e",x"c8",x"87"),
   875 => (x"00",x"00",x"18",x"4c"),
   876 => (x"19",x"8a",x"27",x"1e"),
   877 => (x"27",x"1e",x"00",x"00"),
   878 => (x"00",x"00",x"0a",x"61"),
   879 => (x"70",x"86",x"cc",x"0f"),
   880 => (x"02",x"9a",x"72",x"4a"),
   881 => (x"c0",x"87",x"c5",x"c0"),
   882 => (x"87",x"ff",x"c4",x"48"),
   883 => (x"00",x"1b",x"38",x"27"),
   884 => (x"73",x"4b",x"bf",x"00"),
   885 => (x"27",x"30",x"c4",x"48"),
   886 => (x"00",x"00",x"1b",x"68"),
   887 => (x"1b",x"5c",x"27",x"58"),
   888 => (x"73",x"49",x"00",x"00"),
   889 => (x"19",x"5d",x"27",x"79"),
   890 => (x"bf",x"97",x"00",x"00"),
   891 => (x"9a",x"ff",x"c3",x"4a"),
   892 => (x"5c",x"27",x"32",x"c8"),
   893 => (x"97",x"00",x"00",x"19"),
   894 => (x"ff",x"c3",x"4c",x"bf"),
   895 => (x"27",x"82",x"74",x"9c"),
   896 => (x"00",x"00",x"19",x"5e"),
   897 => (x"c3",x"4c",x"bf",x"97"),
   898 => (x"34",x"d0",x"9c",x"ff"),
   899 => (x"5f",x"27",x"82",x"74"),
   900 => (x"97",x"00",x"00",x"19"),
   901 => (x"ff",x"c3",x"4c",x"bf"),
   902 => (x"74",x"34",x"d8",x"9c"),
   903 => (x"1b",x"68",x"27",x"82"),
   904 => (x"72",x"49",x"00",x"00"),
   905 => (x"1b",x"60",x"27",x"79"),
   906 => (x"92",x"bf",x"00",x"00"),
   907 => (x"00",x"1b",x"4c",x"27"),
   908 => (x"27",x"82",x"bf",x"00"),
   909 => (x"00",x"00",x"1b",x"50"),
   910 => (x"27",x"79",x"72",x"49"),
   911 => (x"00",x"00",x"19",x"65"),
   912 => (x"c3",x"4c",x"bf",x"97"),
   913 => (x"34",x"c8",x"9c",x"ff"),
   914 => (x"00",x"19",x"64",x"27"),
   915 => (x"4d",x"bf",x"97",x"00"),
   916 => (x"75",x"9d",x"ff",x"c3"),
   917 => (x"19",x"66",x"27",x"84"),
   918 => (x"bf",x"97",x"00",x"00"),
   919 => (x"9d",x"ff",x"c3",x"4d"),
   920 => (x"84",x"75",x"35",x"d0"),
   921 => (x"00",x"19",x"67",x"27"),
   922 => (x"4d",x"bf",x"97",x"00"),
   923 => (x"cf",x"9d",x"ff",x"c3"),
   924 => (x"75",x"35",x"d8",x"9d"),
   925 => (x"1b",x"54",x"27",x"84"),
   926 => (x"74",x"49",x"00",x"00"),
   927 => (x"74",x"8c",x"c2",x"79"),
   928 => (x"72",x"48",x"73",x"93"),
   929 => (x"1b",x"5c",x"27",x"80"),
   930 => (x"c1",x"58",x"00",x"00"),
   931 => (x"4a",x"27",x"87",x"fb"),
   932 => (x"97",x"00",x"00",x"19"),
   933 => (x"ff",x"c3",x"4a",x"bf"),
   934 => (x"27",x"32",x"c8",x"9a"),
   935 => (x"00",x"00",x"19",x"49"),
   936 => (x"c3",x"4b",x"bf",x"97"),
   937 => (x"82",x"73",x"9b",x"ff"),
   938 => (x"00",x"1b",x"64",x"27"),
   939 => (x"79",x"72",x"49",x"00"),
   940 => (x"ff",x"c7",x"32",x"c5"),
   941 => (x"27",x"2a",x"c9",x"82"),
   942 => (x"00",x"00",x"1b",x"5c"),
   943 => (x"27",x"79",x"72",x"49"),
   944 => (x"00",x"00",x"19",x"4f"),
   945 => (x"c3",x"4b",x"bf",x"97"),
   946 => (x"33",x"c8",x"9b",x"ff"),
   947 => (x"00",x"19",x"4e",x"27"),
   948 => (x"4c",x"bf",x"97",x"00"),
   949 => (x"74",x"9c",x"ff",x"c3"),
   950 => (x"1b",x"68",x"27",x"83"),
   951 => (x"73",x"49",x"00",x"00"),
   952 => (x"1b",x"60",x"27",x"79"),
   953 => (x"93",x"bf",x"00",x"00"),
   954 => (x"00",x"1b",x"4c",x"27"),
   955 => (x"27",x"83",x"bf",x"00"),
   956 => (x"00",x"00",x"1b",x"58"),
   957 => (x"27",x"79",x"73",x"49"),
   958 => (x"00",x"00",x"1b",x"54"),
   959 => (x"73",x"79",x"c0",x"49"),
   960 => (x"27",x"80",x"72",x"48"),
   961 => (x"00",x"00",x"1b",x"54"),
   962 => (x"26",x"48",x"c1",x"58"),
   963 => (x"26",x"4c",x"26",x"4d"),
   964 => (x"26",x"4a",x"26",x"4b"),
   965 => (x"5a",x"5e",x"0e",x"4f"),
   966 => (x"0e",x"5d",x"5c",x"5b"),
   967 => (x"00",x"1b",x"40",x"27"),
   968 => (x"c0",x"02",x"bf",x"00"),
   969 => (x"66",x"d4",x"87",x"cf"),
   970 => (x"2d",x"b7",x"c7",x"4d"),
   971 => (x"c1",x"4b",x"66",x"d4"),
   972 => (x"cc",x"c0",x"9b",x"ff"),
   973 => (x"4d",x"66",x"d4",x"87"),
   974 => (x"d4",x"2d",x"b7",x"c8"),
   975 => (x"ff",x"c3",x"4b",x"66"),
   976 => (x"19",x"38",x"27",x"9b"),
   977 => (x"27",x"1e",x"00",x"00"),
   978 => (x"00",x"00",x"1b",x"4c"),
   979 => (x"82",x"75",x"4a",x"bf"),
   980 => (x"f4",x"27",x"1e",x"72"),
   981 => (x"0f",x"00",x"00",x"07"),
   982 => (x"4a",x"70",x"86",x"c8"),
   983 => (x"c0",x"05",x"9a",x"72"),
   984 => (x"48",x"c0",x"87",x"c5"),
   985 => (x"27",x"87",x"f2",x"c0"),
   986 => (x"00",x"00",x"1b",x"40"),
   987 => (x"d5",x"c0",x"02",x"bf"),
   988 => (x"c4",x"4a",x"73",x"87"),
   989 => (x"19",x"38",x"27",x"92"),
   990 => (x"6a",x"82",x"00",x"00"),
   991 => (x"ff",x"ff",x"cf",x"4c"),
   992 => (x"c0",x"9c",x"ff",x"ff"),
   993 => (x"4a",x"73",x"87",x"d1"),
   994 => (x"38",x"27",x"92",x"c2"),
   995 => (x"82",x"00",x"00",x"19"),
   996 => (x"cf",x"4c",x"6a",x"9f"),
   997 => (x"74",x"9c",x"ff",x"ff"),
   998 => (x"26",x"4d",x"26",x"48"),
   999 => (x"26",x"4b",x"26",x"4c"),
  1000 => (x"0e",x"4f",x"26",x"4a"),
  1001 => (x"5c",x"5b",x"5a",x"5e"),
  1002 => (x"8e",x"cc",x"0e",x"5d"),
  1003 => (x"ff",x"ff",x"ff",x"cf"),
  1004 => (x"4c",x"c0",x"4d",x"f8"),
  1005 => (x"54",x"27",x"49",x"76"),
  1006 => (x"bf",x"00",x"00",x"1b"),
  1007 => (x"49",x"a6",x"c4",x"79"),
  1008 => (x"00",x"1b",x"58",x"27"),
  1009 => (x"27",x"79",x"bf",x"00"),
  1010 => (x"00",x"00",x"1b",x"40"),
  1011 => (x"cc",x"c0",x"02",x"bf"),
  1012 => (x"1b",x"38",x"27",x"87"),
  1013 => (x"4a",x"bf",x"00",x"00"),
  1014 => (x"c9",x"c0",x"32",x"c4"),
  1015 => (x"1b",x"5c",x"27",x"87"),
  1016 => (x"4a",x"bf",x"00",x"00"),
  1017 => (x"a6",x"c8",x"32",x"c4"),
  1018 => (x"c0",x"79",x"72",x"49"),
  1019 => (x"49",x"66",x"c8",x"4b"),
  1020 => (x"c3",x"06",x"a9",x"c0"),
  1021 => (x"4a",x"73",x"87",x"e0"),
  1022 => (x"9a",x"72",x"9a",x"cf"),
  1023 => (x"87",x"e4",x"c0",x"05"),
  1024 => (x"00",x"19",x"38",x"27"),
  1025 => (x"66",x"c8",x"1e",x"00"),
  1026 => (x"48",x"66",x"c8",x"4a"),
  1027 => (x"a6",x"cc",x"80",x"c1"),
  1028 => (x"27",x"1e",x"72",x"58"),
  1029 => (x"00",x"00",x"07",x"f4"),
  1030 => (x"27",x"86",x"c8",x"0f"),
  1031 => (x"00",x"00",x"19",x"38"),
  1032 => (x"87",x"c3",x"c0",x"4c"),
  1033 => (x"97",x"84",x"e0",x"c0"),
  1034 => (x"ff",x"c3",x"4a",x"6c"),
  1035 => (x"02",x"9a",x"72",x"9a"),
  1036 => (x"97",x"87",x"da",x"c2"),
  1037 => (x"ff",x"c3",x"4a",x"6c"),
  1038 => (x"aa",x"e5",x"c3",x"9a"),
  1039 => (x"87",x"cd",x"c2",x"02"),
  1040 => (x"82",x"cb",x"4a",x"74"),
  1041 => (x"c3",x"4a",x"6a",x"97"),
  1042 => (x"9a",x"d8",x"9a",x"ff"),
  1043 => (x"c1",x"05",x"9a",x"72"),
  1044 => (x"1e",x"74",x"87",x"fb"),
  1045 => (x"00",x"00",x"61",x"27"),
  1046 => (x"86",x"c4",x"0f",x"00"),
  1047 => (x"e8",x"c0",x"1e",x"cb"),
  1048 => (x"1e",x"74",x"1e",x"66"),
  1049 => (x"00",x"0a",x"61",x"27"),
  1050 => (x"86",x"cc",x"0f",x"00"),
  1051 => (x"9a",x"72",x"4a",x"70"),
  1052 => (x"87",x"d9",x"c1",x"05"),
  1053 => (x"83",x"dc",x"4b",x"74"),
  1054 => (x"4a",x"66",x"e0",x"c0"),
  1055 => (x"7a",x"6b",x"82",x"c4"),
  1056 => (x"83",x"da",x"4b",x"74"),
  1057 => (x"4a",x"66",x"e0",x"c0"),
  1058 => (x"6b",x"9f",x"82",x"c8"),
  1059 => (x"ff",x"ff",x"cf",x"48"),
  1060 => (x"72",x"7a",x"70",x"98"),
  1061 => (x"1b",x"40",x"27",x"4d"),
  1062 => (x"02",x"bf",x"00",x"00"),
  1063 => (x"74",x"87",x"d9",x"c0"),
  1064 => (x"9f",x"82",x"d4",x"4a"),
  1065 => (x"ff",x"cf",x"4a",x"6a"),
  1066 => (x"ff",x"c0",x"9a",x"ff"),
  1067 => (x"48",x"72",x"9a",x"ff"),
  1068 => (x"a6",x"c4",x"30",x"d0"),
  1069 => (x"87",x"c4",x"c0",x"58"),
  1070 => (x"79",x"c0",x"49",x"76"),
  1071 => (x"80",x"6d",x"48",x"6e"),
  1072 => (x"e0",x"c0",x"7d",x"70"),
  1073 => (x"79",x"c0",x"49",x"66"),
  1074 => (x"cc",x"c1",x"48",x"c1"),
  1075 => (x"c8",x"83",x"c1",x"87"),
  1076 => (x"fc",x"04",x"ab",x"66"),
  1077 => (x"ff",x"cf",x"87",x"e0"),
  1078 => (x"4d",x"f8",x"ff",x"ff"),
  1079 => (x"00",x"1b",x"40",x"27"),
  1080 => (x"c0",x"02",x"bf",x"00"),
  1081 => (x"1e",x"6e",x"87",x"f1"),
  1082 => (x"00",x"0f",x"15",x"27"),
  1083 => (x"86",x"c4",x"0f",x"00"),
  1084 => (x"6e",x"58",x"a6",x"c4"),
  1085 => (x"75",x"9a",x"75",x"4a"),
  1086 => (x"da",x"c0",x"02",x"aa"),
  1087 => (x"c2",x"4a",x"6e",x"87"),
  1088 => (x"1b",x"38",x"27",x"8a"),
  1089 => (x"92",x"bf",x"00",x"00"),
  1090 => (x"00",x"1b",x"50",x"27"),
  1091 => (x"72",x"48",x"bf",x"00"),
  1092 => (x"58",x"a6",x"c8",x"80"),
  1093 => (x"c0",x"87",x"d4",x"fb"),
  1094 => (x"ff",x"ff",x"cf",x"48"),
  1095 => (x"cc",x"4d",x"f8",x"ff"),
  1096 => (x"26",x"4d",x"26",x"86"),
  1097 => (x"26",x"4b",x"26",x"4c"),
  1098 => (x"0e",x"4f",x"26",x"4a"),
  1099 => (x"0e",x"5b",x"5a",x"5e"),
  1100 => (x"4a",x"bf",x"66",x"cc"),
  1101 => (x"66",x"cc",x"82",x"c1"),
  1102 => (x"27",x"79",x"72",x"49"),
  1103 => (x"00",x"00",x"1b",x"3c"),
  1104 => (x"9a",x"72",x"9a",x"bf"),
  1105 => (x"87",x"d3",x"c0",x"05"),
  1106 => (x"c8",x"4a",x"66",x"cc"),
  1107 => (x"27",x"1e",x"6a",x"82"),
  1108 => (x"00",x"00",x"0f",x"15"),
  1109 => (x"70",x"86",x"c4",x"0f"),
  1110 => (x"c1",x"7a",x"73",x"4b"),
  1111 => (x"26",x"4b",x"26",x"48"),
  1112 => (x"0e",x"4f",x"26",x"4a"),
  1113 => (x"0e",x"5b",x"5a",x"5e"),
  1114 => (x"00",x"1b",x"50",x"27"),
  1115 => (x"cc",x"4a",x"bf",x"00"),
  1116 => (x"83",x"c8",x"4b",x"66"),
  1117 => (x"8b",x"c2",x"4b",x"6b"),
  1118 => (x"00",x"1b",x"38",x"27"),
  1119 => (x"73",x"93",x"bf",x"00"),
  1120 => (x"1b",x"3c",x"27",x"82"),
  1121 => (x"4b",x"bf",x"00",x"00"),
  1122 => (x"9b",x"bf",x"66",x"cc"),
  1123 => (x"66",x"d0",x"82",x"73"),
  1124 => (x"27",x"1e",x"72",x"1e"),
  1125 => (x"00",x"00",x"07",x"f4"),
  1126 => (x"70",x"86",x"c8",x"0f"),
  1127 => (x"05",x"9a",x"72",x"4a"),
  1128 => (x"c0",x"87",x"c5",x"c0"),
  1129 => (x"87",x"c2",x"c0",x"48"),
  1130 => (x"4b",x"26",x"48",x"c1"),
  1131 => (x"4f",x"26",x"4a",x"26"),
  1132 => (x"5b",x"5a",x"5e",x"0e"),
  1133 => (x"d8",x"0e",x"5d",x"5c"),
  1134 => (x"66",x"d4",x"4c",x"66"),
  1135 => (x"1b",x"70",x"27",x"1e"),
  1136 => (x"27",x"1e",x"00",x"00"),
  1137 => (x"00",x"00",x"0f",x"a3"),
  1138 => (x"70",x"86",x"c8",x"0f"),
  1139 => (x"02",x"9a",x"72",x"4a"),
  1140 => (x"27",x"87",x"df",x"c1"),
  1141 => (x"00",x"00",x"1b",x"74"),
  1142 => (x"ff",x"c7",x"4a",x"bf"),
  1143 => (x"72",x"2a",x"c9",x"82"),
  1144 => (x"27",x"4b",x"c0",x"4d"),
  1145 => (x"00",x"00",x"12",x"54"),
  1146 => (x"00",x"61",x"27",x"1e"),
  1147 => (x"c4",x"0f",x"00",x"00"),
  1148 => (x"ad",x"b7",x"c0",x"86"),
  1149 => (x"87",x"d0",x"c1",x"06"),
  1150 => (x"70",x"27",x"1e",x"74"),
  1151 => (x"1e",x"00",x"00",x"1b"),
  1152 => (x"00",x"11",x"63",x"27"),
  1153 => (x"86",x"c8",x"0f",x"00"),
  1154 => (x"9a",x"72",x"4a",x"70"),
  1155 => (x"87",x"c5",x"c0",x"05"),
  1156 => (x"f5",x"c0",x"48",x"c0"),
  1157 => (x"1b",x"70",x"27",x"87"),
  1158 => (x"27",x"1e",x"00",x"00"),
  1159 => (x"00",x"00",x"11",x"2b"),
  1160 => (x"c8",x"86",x"c4",x"0f"),
  1161 => (x"83",x"c1",x"84",x"c0"),
  1162 => (x"04",x"ab",x"b7",x"75"),
  1163 => (x"c0",x"87",x"c9",x"ff"),
  1164 => (x"66",x"d4",x"87",x"d6"),
  1165 => (x"12",x"6d",x"27",x"1e"),
  1166 => (x"27",x"1e",x"00",x"00"),
  1167 => (x"00",x"00",x"00",x"9a"),
  1168 => (x"c0",x"86",x"c8",x"0f"),
  1169 => (x"87",x"c2",x"c0",x"48"),
  1170 => (x"4d",x"26",x"48",x"c1"),
  1171 => (x"4b",x"26",x"4c",x"26"),
  1172 => (x"4f",x"26",x"4a",x"26"),
  1173 => (x"6e",x"65",x"70",x"4f"),
  1174 => (x"66",x"20",x"64",x"65"),
  1175 => (x"2c",x"65",x"6c",x"69"),
  1176 => (x"61",x"6f",x"6c",x"20"),
  1177 => (x"67",x"6e",x"69",x"64"),
  1178 => (x"0a",x"2e",x"2e",x"2e"),
  1179 => (x"6e",x"61",x"43",x"00"),
  1180 => (x"6f",x"20",x"74",x"27"),
  1181 => (x"20",x"6e",x"65",x"70"),
  1182 => (x"00",x"0a",x"73",x"25"),
  1183 => (x"5b",x"5a",x"5e",x"0e"),
  1184 => (x"4a",x"66",x"cc",x"0e"),
  1185 => (x"ff",x"c3",x"2a",x"d8"),
  1186 => (x"4b",x"66",x"cc",x"9a"),
  1187 => (x"fc",x"cf",x"2b",x"c8"),
  1188 => (x"b2",x"73",x"9b",x"c0"),
  1189 => (x"c8",x"4b",x"66",x"cc"),
  1190 => (x"f0",x"ff",x"c0",x"33"),
  1191 => (x"73",x"9b",x"c0",x"c0"),
  1192 => (x"4b",x"66",x"cc",x"b2"),
  1193 => (x"c0",x"ff",x"33",x"d8"),
  1194 => (x"9b",x"c0",x"c0",x"c0"),
  1195 => (x"48",x"72",x"b2",x"73"),
  1196 => (x"4a",x"26",x"4b",x"26"),
  1197 => (x"5e",x"0e",x"4f",x"26"),
  1198 => (x"cc",x"0e",x"5b",x"5a"),
  1199 => (x"2b",x"c8",x"4b",x"66"),
  1200 => (x"cc",x"9b",x"ff",x"c3"),
  1201 => (x"32",x"c8",x"4a",x"66"),
  1202 => (x"9a",x"c0",x"fc",x"cf"),
  1203 => (x"9b",x"ff",x"ff",x"cf"),
  1204 => (x"ff",x"cf",x"b2",x"73"),
  1205 => (x"48",x"72",x"9a",x"ff"),
  1206 => (x"4a",x"26",x"4b",x"26"),
  1207 => (x"5e",x"0e",x"4f",x"26"),
  1208 => (x"cc",x"0e",x"5b",x"5a"),
  1209 => (x"2a",x"d0",x"4a",x"66"),
  1210 => (x"9a",x"ff",x"ff",x"cf"),
  1211 => (x"d0",x"4b",x"66",x"cc"),
  1212 => (x"c0",x"c0",x"f0",x"33"),
  1213 => (x"72",x"b2",x"73",x"9b"),
  1214 => (x"26",x"4b",x"26",x"48"),
  1215 => (x"1e",x"4f",x"26",x"4a"),
  1216 => (x"c0",x"d0",x"1e",x"72"),
  1217 => (x"4a",x"c0",x"c0",x"c0"),
  1218 => (x"fd",x"ff",x"0f",x"72"),
  1219 => (x"26",x"4a",x"26",x"87"),
  1220 => (x"1e",x"72",x"1e",x"4f"),
  1221 => (x"c3",x"4a",x"66",x"cc"),
  1222 => (x"f7",x"c0",x"9a",x"df"),
  1223 => (x"aa",x"b7",x"c0",x"8a"),
  1224 => (x"87",x"c3",x"c0",x"03"),
  1225 => (x"c8",x"82",x"e7",x"c0"),
  1226 => (x"30",x"c4",x"48",x"66"),
  1227 => (x"c8",x"58",x"a6",x"cc"),
  1228 => (x"b0",x"72",x"48",x"66"),
  1229 => (x"c8",x"58",x"a6",x"cc"),
  1230 => (x"4a",x"26",x"48",x"66"),
  1231 => (x"5e",x"0e",x"4f",x"26"),
  1232 => (x"5d",x"5c",x"5b",x"5a"),
  1233 => (x"c0",x"c0",x"d0",x"0e"),
  1234 => (x"27",x"4d",x"c0",x"c0"),
  1235 => (x"00",x"00",x"1b",x"7c"),
  1236 => (x"80",x"c1",x"48",x"bf"),
  1237 => (x"00",x"1b",x"80",x"27"),
  1238 => (x"d4",x"97",x"58",x"00"),
  1239 => (x"c0",x"c1",x"4a",x"66"),
  1240 => (x"92",x"c0",x"c0",x"c0"),
  1241 => (x"92",x"b7",x"c0",x"c4"),
  1242 => (x"aa",x"d3",x"c1",x"4a"),
  1243 => (x"87",x"e9",x"c0",x"05"),
  1244 => (x"00",x"1b",x"7c",x"27"),
  1245 => (x"79",x"c0",x"49",x"00"),
  1246 => (x"00",x"1b",x"80",x"27"),
  1247 => (x"79",x"c0",x"49",x"00"),
  1248 => (x"00",x"1b",x"88",x"27"),
  1249 => (x"79",x"c0",x"49",x"00"),
  1250 => (x"00",x"1b",x"8c",x"27"),
  1251 => (x"79",x"c0",x"49",x"00"),
  1252 => (x"c1",x"49",x"c0",x"ff"),
  1253 => (x"ca",x"ca",x"79",x"d3"),
  1254 => (x"1b",x"7c",x"27",x"87"),
  1255 => (x"49",x"bf",x"00",x"00"),
  1256 => (x"c1",x"05",x"a9",x"c1"),
  1257 => (x"c0",x"ff",x"87",x"db"),
  1258 => (x"79",x"f4",x"c1",x"49"),
  1259 => (x"4a",x"66",x"d4",x"97"),
  1260 => (x"c0",x"c0",x"c0",x"c1"),
  1261 => (x"c0",x"c4",x"92",x"c0"),
  1262 => (x"72",x"4a",x"92",x"b7"),
  1263 => (x"1b",x"8c",x"27",x"1e"),
  1264 => (x"1e",x"bf",x"00",x"00"),
  1265 => (x"00",x"13",x"11",x"27"),
  1266 => (x"86",x"c8",x"0f",x"00"),
  1267 => (x"00",x"1b",x"90",x"27"),
  1268 => (x"8c",x"27",x"58",x"00"),
  1269 => (x"bf",x"00",x"00",x"1b"),
  1270 => (x"ac",x"b7",x"c3",x"4c"),
  1271 => (x"87",x"c6",x"c0",x"06"),
  1272 => (x"88",x"74",x"48",x"ca"),
  1273 => (x"4a",x"74",x"4c",x"70"),
  1274 => (x"48",x"72",x"82",x"c1"),
  1275 => (x"88",x"27",x"30",x"c1"),
  1276 => (x"58",x"00",x"00",x"1b"),
  1277 => (x"f0",x"c0",x"48",x"74"),
  1278 => (x"49",x"c0",x"ff",x"80"),
  1279 => (x"e2",x"c8",x"79",x"70"),
  1280 => (x"1b",x"8c",x"27",x"87"),
  1281 => (x"49",x"bf",x"00",x"00"),
  1282 => (x"01",x"a9",x"b7",x"c9"),
  1283 => (x"27",x"87",x"d4",x"c8"),
  1284 => (x"00",x"00",x"1b",x"8c"),
  1285 => (x"b7",x"c0",x"49",x"bf"),
  1286 => (x"c6",x"c8",x"06",x"a9"),
  1287 => (x"1b",x"8c",x"27",x"87"),
  1288 => (x"48",x"bf",x"00",x"00"),
  1289 => (x"ff",x"80",x"f0",x"c0"),
  1290 => (x"79",x"70",x"49",x"c0"),
  1291 => (x"00",x"1b",x"7c",x"27"),
  1292 => (x"c3",x"49",x"bf",x"00"),
  1293 => (x"c0",x"01",x"a9",x"b7"),
  1294 => (x"d4",x"97",x"87",x"e9"),
  1295 => (x"c0",x"c1",x"4a",x"66"),
  1296 => (x"92",x"c0",x"c0",x"c0"),
  1297 => (x"92",x"b7",x"c0",x"c4"),
  1298 => (x"27",x"1e",x"72",x"4a"),
  1299 => (x"00",x"00",x"1b",x"88"),
  1300 => (x"11",x"27",x"1e",x"bf"),
  1301 => (x"0f",x"00",x"00",x"13"),
  1302 => (x"8c",x"27",x"86",x"c8"),
  1303 => (x"58",x"00",x"00",x"1b"),
  1304 => (x"27",x"87",x"c0",x"c7"),
  1305 => (x"00",x"00",x"1b",x"84"),
  1306 => (x"82",x"c3",x"4a",x"bf"),
  1307 => (x"00",x"1b",x"7c",x"27"),
  1308 => (x"72",x"49",x"bf",x"00"),
  1309 => (x"c0",x"01",x"a9",x"b7"),
  1310 => (x"d4",x"97",x"87",x"f1"),
  1311 => (x"c0",x"c1",x"4a",x"66"),
  1312 => (x"92",x"c0",x"c0",x"c0"),
  1313 => (x"92",x"b7",x"c0",x"c4"),
  1314 => (x"27",x"1e",x"72",x"4a"),
  1315 => (x"00",x"00",x"1b",x"80"),
  1316 => (x"11",x"27",x"1e",x"bf"),
  1317 => (x"0f",x"00",x"00",x"13"),
  1318 => (x"84",x"27",x"86",x"c8"),
  1319 => (x"58",x"00",x"00",x"1b"),
  1320 => (x"00",x"1b",x"90",x"27"),
  1321 => (x"79",x"c1",x"49",x"00"),
  1322 => (x"27",x"87",x"f8",x"c5"),
  1323 => (x"00",x"00",x"1b",x"8c"),
  1324 => (x"b7",x"c0",x"49",x"bf"),
  1325 => (x"d0",x"c3",x"06",x"a9"),
  1326 => (x"1b",x"8c",x"27",x"87"),
  1327 => (x"49",x"bf",x"00",x"00"),
  1328 => (x"01",x"a9",x"b7",x"c3"),
  1329 => (x"27",x"87",x"c2",x"c3"),
  1330 => (x"00",x"00",x"1b",x"88"),
  1331 => (x"32",x"c1",x"4a",x"bf"),
  1332 => (x"7c",x"27",x"82",x"c1"),
  1333 => (x"bf",x"00",x"00",x"1b"),
  1334 => (x"a9",x"b7",x"72",x"49"),
  1335 => (x"87",x"c2",x"c2",x"01"),
  1336 => (x"4a",x"66",x"d4",x"97"),
  1337 => (x"c0",x"c0",x"c0",x"c1"),
  1338 => (x"c0",x"c4",x"92",x"c0"),
  1339 => (x"72",x"4a",x"92",x"b7"),
  1340 => (x"1b",x"94",x"27",x"1e"),
  1341 => (x"1e",x"bf",x"00",x"00"),
  1342 => (x"00",x"13",x"11",x"27"),
  1343 => (x"86",x"c8",x"0f",x"00"),
  1344 => (x"00",x"1b",x"98",x"27"),
  1345 => (x"90",x"27",x"58",x"00"),
  1346 => (x"bf",x"00",x"00",x"1b"),
  1347 => (x"27",x"8a",x"c1",x"4a"),
  1348 => (x"00",x"00",x"1b",x"90"),
  1349 => (x"c0",x"79",x"72",x"49"),
  1350 => (x"c4",x"03",x"aa",x"b7"),
  1351 => (x"80",x"27",x"87",x"c5"),
  1352 => (x"bf",x"00",x"00",x"1b"),
  1353 => (x"1b",x"94",x"27",x"4a"),
  1354 => (x"bf",x"97",x"00",x"00"),
  1355 => (x"1b",x"80",x"27",x"52"),
  1356 => (x"4a",x"bf",x"00",x"00"),
  1357 => (x"80",x"27",x"82",x"c1"),
  1358 => (x"49",x"00",x"00",x"1b"),
  1359 => (x"98",x"27",x"79",x"72"),
  1360 => (x"bf",x"00",x"00",x"1b"),
  1361 => (x"c0",x"06",x"aa",x"b7"),
  1362 => (x"98",x"27",x"87",x"cd"),
  1363 => (x"49",x"00",x"00",x"1b"),
  1364 => (x"00",x"1b",x"80",x"27"),
  1365 => (x"27",x"79",x"bf",x"00"),
  1366 => (x"00",x"00",x"1b",x"90"),
  1367 => (x"c3",x"79",x"c1",x"49"),
  1368 => (x"90",x"27",x"87",x"c1"),
  1369 => (x"bf",x"00",x"00",x"1b"),
  1370 => (x"87",x"f7",x"c2",x"05"),
  1371 => (x"00",x"1b",x"94",x"27"),
  1372 => (x"c4",x"4a",x"bf",x"00"),
  1373 => (x"1b",x"94",x"27",x"32"),
  1374 => (x"72",x"49",x"00",x"00"),
  1375 => (x"1b",x"80",x"27",x"79"),
  1376 => (x"49",x"bf",x"00",x"00"),
  1377 => (x"da",x"c2",x"51",x"72"),
  1378 => (x"1b",x"8c",x"27",x"87"),
  1379 => (x"49",x"bf",x"00",x"00"),
  1380 => (x"04",x"a9",x"b7",x"c7"),
  1381 => (x"c0",x"87",x"fd",x"c1"),
  1382 => (x"49",x"f4",x"fe",x"4b"),
  1383 => (x"98",x"27",x"79",x"c1"),
  1384 => (x"bf",x"00",x"00",x"1b"),
  1385 => (x"27",x"1e",x"75",x"1e"),
  1386 => (x"00",x"00",x"18",x"ec"),
  1387 => (x"00",x"9a",x"27",x"1e"),
  1388 => (x"cc",x"0f",x"00",x"00"),
  1389 => (x"1b",x"80",x"27",x"86"),
  1390 => (x"75",x"49",x"00",x"00"),
  1391 => (x"1b",x"80",x"27",x"79"),
  1392 => (x"49",x"bf",x"00",x"00"),
  1393 => (x"00",x"1b",x"98",x"27"),
  1394 => (x"a9",x"b7",x"bf",x"00"),
  1395 => (x"87",x"e5",x"c0",x"03"),
  1396 => (x"00",x"1b",x"80",x"27"),
  1397 => (x"83",x"bf",x"bf",x"00"),
  1398 => (x"00",x"1b",x"80",x"27"),
  1399 => (x"c4",x"4a",x"bf",x"00"),
  1400 => (x"1b",x"80",x"27",x"82"),
  1401 => (x"72",x"49",x"00",x"00"),
  1402 => (x"1b",x"98",x"27",x"79"),
  1403 => (x"b7",x"bf",x"00",x"00"),
  1404 => (x"db",x"ff",x"04",x"aa"),
  1405 => (x"27",x"1e",x"73",x"87"),
  1406 => (x"00",x"00",x"19",x"0b"),
  1407 => (x"00",x"9a",x"27",x"1e"),
  1408 => (x"c8",x"0f",x"00",x"00"),
  1409 => (x"49",x"c0",x"ff",x"86"),
  1410 => (x"27",x"79",x"c2",x"c1"),
  1411 => (x"00",x"00",x"12",x"ff"),
  1412 => (x"87",x"cf",x"c0",x"0f"),
  1413 => (x"00",x"1b",x"8c",x"27"),
  1414 => (x"c0",x"48",x"bf",x"00"),
  1415 => (x"c0",x"ff",x"80",x"f0"),
  1416 => (x"26",x"79",x"70",x"49"),
  1417 => (x"26",x"4c",x"26",x"4d"),
  1418 => (x"26",x"4a",x"26",x"4b"),
  1419 => (x"5a",x"5e",x"0e",x"4f"),
  1420 => (x"0e",x"5d",x"5c",x"5b"),
  1421 => (x"17",x"3f",x"27",x"1e"),
  1422 => (x"27",x"1e",x"00",x"00"),
  1423 => (x"00",x"00",x"00",x"61"),
  1424 => (x"27",x"86",x"c4",x"0f"),
  1425 => (x"00",x"00",x"04",x"fd"),
  1426 => (x"72",x"4a",x"70",x"0f"),
  1427 => (x"d3",x"c0",x"02",x"9a"),
  1428 => (x"0a",x"be",x"27",x"87"),
  1429 => (x"70",x"0f",x"00",x"00"),
  1430 => (x"02",x"9a",x"72",x"4a"),
  1431 => (x"c1",x"87",x"c5",x"c0"),
  1432 => (x"87",x"c2",x"c0",x"4a"),
  1433 => (x"49",x"76",x"4a",x"c0"),
  1434 => (x"55",x"27",x"79",x"72"),
  1435 => (x"1e",x"00",x"00",x"17"),
  1436 => (x"00",x"00",x"61",x"27"),
  1437 => (x"86",x"c4",x"0f",x"00"),
  1438 => (x"00",x"1b",x"98",x"27"),
  1439 => (x"79",x"c0",x"49",x"00"),
  1440 => (x"27",x"1e",x"ee",x"c0"),
  1441 => (x"00",x"00",x"00",x"42"),
  1442 => (x"c3",x"86",x"c4",x"0f"),
  1443 => (x"4b",x"ff",x"c8",x"f4"),
  1444 => (x"4c",x"bf",x"c0",x"ff"),
  1445 => (x"c0",x"c8",x"4a",x"74"),
  1446 => (x"02",x"9a",x"72",x"9a"),
  1447 => (x"74",x"87",x"e0",x"c1"),
  1448 => (x"9d",x"ff",x"c3",x"4d"),
  1449 => (x"c1",x"05",x"ad",x"db"),
  1450 => (x"02",x"6e",x"87",x"c6"),
  1451 => (x"d0",x"87",x"f3",x"c0"),
  1452 => (x"c0",x"c0",x"c0",x"c0"),
  1453 => (x"17",x"23",x"27",x"1e"),
  1454 => (x"27",x"1e",x"00",x"00"),
  1455 => (x"00",x"00",x"11",x"b0"),
  1456 => (x"70",x"86",x"c8",x"0f"),
  1457 => (x"02",x"9a",x"72",x"4a"),
  1458 => (x"27",x"87",x"d7",x"c0"),
  1459 => (x"00",x"00",x"17",x"17"),
  1460 => (x"00",x"61",x"27",x"1e"),
  1461 => (x"c4",x"0f",x"00",x"00"),
  1462 => (x"12",x"ff",x"27",x"86"),
  1463 => (x"c0",x"0f",x"00",x"00"),
  1464 => (x"2f",x"27",x"87",x"ce"),
  1465 => (x"1e",x"00",x"00",x"17"),
  1466 => (x"00",x"00",x"61",x"27"),
  1467 => (x"86",x"c4",x"0f",x"00"),
  1468 => (x"3e",x"27",x"1e",x"75"),
  1469 => (x"0f",x"00",x"00",x"13"),
  1470 => (x"f4",x"c3",x"86",x"c4"),
  1471 => (x"73",x"4b",x"c0",x"c9"),
  1472 => (x"72",x"8b",x"c1",x"4a"),
  1473 => (x"c7",x"fe",x"05",x"9a"),
  1474 => (x"87",x"f4",x"fd",x"87"),
  1475 => (x"26",x"4d",x"26",x"26"),
  1476 => (x"26",x"4b",x"26",x"4c"),
  1477 => (x"42",x"4f",x"26",x"4a"),
  1478 => (x"69",x"74",x"6f",x"6f"),
  1479 => (x"2e",x"2e",x"67",x"6e"),
  1480 => (x"42",x"00",x"0a",x"2e"),
  1481 => (x"38",x"54",x"4f",x"4f"),
  1482 => (x"42",x"20",x"32",x"33"),
  1483 => (x"53",x"00",x"4e",x"49"),
  1484 => (x"6f",x"62",x"20",x"44"),
  1485 => (x"66",x"20",x"74",x"6f"),
  1486 => (x"65",x"6c",x"69",x"61"),
  1487 => (x"49",x"00",x"0a",x"64"),
  1488 => (x"69",x"74",x"69",x"6e"),
  1489 => (x"7a",x"69",x"6c",x"61"),
  1490 => (x"20",x"67",x"6e",x"69"),
  1491 => (x"63",x"20",x"44",x"53"),
  1492 => (x"0a",x"64",x"72",x"61"),
  1493 => (x"32",x"53",x"52",x"00"),
  1494 => (x"62",x"20",x"32",x"33"),
  1495 => (x"20",x"74",x"6f",x"6f"),
  1496 => (x"72",x"70",x"20",x"2d"),
  1497 => (x"20",x"73",x"73",x"65"),
  1498 => (x"20",x"43",x"53",x"45"),
  1499 => (x"62",x"20",x"6f",x"74"),
  1500 => (x"20",x"74",x"6f",x"6f"),
  1501 => (x"6d",x"6f",x"72",x"66"),
  1502 => (x"2e",x"44",x"53",x"20"),
  1503 => (x"44",x"4d",x"43",x"00"),
  1504 => (x"61",x"65",x"52",x"00"),
  1505 => (x"66",x"6f",x"20",x"64"),
  1506 => (x"52",x"42",x"4d",x"20"),
  1507 => (x"69",x"61",x"66",x"20"),
  1508 => (x"0a",x"64",x"65",x"6c"),
  1509 => (x"20",x"6f",x"4e",x"00"),
  1510 => (x"74",x"72",x"61",x"70"),
  1511 => (x"6f",x"69",x"74",x"69"),
  1512 => (x"69",x"73",x"20",x"6e"),
  1513 => (x"74",x"61",x"6e",x"67"),
  1514 => (x"20",x"65",x"72",x"75"),
  1515 => (x"6e",x"75",x"6f",x"66"),
  1516 => (x"4d",x"00",x"0a",x"64"),
  1517 => (x"69",x"73",x"52",x"42"),
  1518 => (x"20",x"3a",x"65",x"7a"),
  1519 => (x"20",x"2c",x"64",x"25"),
  1520 => (x"74",x"72",x"61",x"70"),
  1521 => (x"6f",x"69",x"74",x"69"),
  1522 => (x"7a",x"69",x"73",x"6e"),
  1523 => (x"25",x"20",x"3a",x"65"),
  1524 => (x"6f",x"20",x"2c",x"64"),
  1525 => (x"65",x"73",x"66",x"66"),
  1526 => (x"66",x"6f",x"20",x"74"),
  1527 => (x"67",x"69",x"73",x"20"),
  1528 => (x"64",x"25",x"20",x"3a"),
  1529 => (x"69",x"73",x"20",x"2c"),
  1530 => (x"78",x"30",x"20",x"67"),
  1531 => (x"00",x"0a",x"78",x"25"),
  1532 => (x"64",x"61",x"65",x"52"),
  1533 => (x"20",x"67",x"6e",x"69"),
  1534 => (x"74",x"6f",x"6f",x"62"),
  1535 => (x"63",x"65",x"73",x"20"),
  1536 => (x"20",x"72",x"6f",x"74"),
  1537 => (x"00",x"0a",x"64",x"25"),
  1538 => (x"64",x"61",x"65",x"52"),
  1539 => (x"6f",x"6f",x"62",x"20"),
  1540 => (x"65",x"73",x"20",x"74"),
  1541 => (x"72",x"6f",x"74",x"63"),
  1542 => (x"6f",x"72",x"66",x"20"),
  1543 => (x"69",x"66",x"20",x"6d"),
  1544 => (x"20",x"74",x"73",x"72"),
  1545 => (x"74",x"72",x"61",x"70"),
  1546 => (x"6f",x"69",x"74",x"69"),
  1547 => (x"55",x"00",x"0a",x"6e"),
  1548 => (x"70",x"75",x"73",x"6e"),
  1549 => (x"74",x"72",x"6f",x"70"),
  1550 => (x"70",x"20",x"64",x"65"),
  1551 => (x"69",x"74",x"72",x"61"),
  1552 => (x"6e",x"6f",x"69",x"74"),
  1553 => (x"70",x"79",x"74",x"20"),
  1554 => (x"00",x"0d",x"21",x"65"),
  1555 => (x"33",x"54",x"41",x"46"),
  1556 => (x"20",x"20",x"20",x"32"),
  1557 => (x"61",x"65",x"52",x"00"),
  1558 => (x"67",x"6e",x"69",x"64"),
  1559 => (x"52",x"42",x"4d",x"20"),
  1560 => (x"42",x"4d",x"00",x"0a"),
  1561 => (x"75",x"73",x"20",x"52"),
  1562 => (x"73",x"65",x"63",x"63"),
  1563 => (x"6c",x"75",x"66",x"73"),
  1564 => (x"72",x"20",x"79",x"6c"),
  1565 => (x"0a",x"64",x"61",x"65"),
  1566 => (x"54",x"41",x"46",x"00"),
  1567 => (x"20",x"20",x"36",x"31"),
  1568 => (x"41",x"46",x"00",x"20"),
  1569 => (x"20",x"32",x"33",x"54"),
  1570 => (x"50",x"00",x"20",x"20"),
  1571 => (x"69",x"74",x"72",x"61"),
  1572 => (x"6e",x"6f",x"69",x"74"),
  1573 => (x"6e",x"75",x"6f",x"63"),
  1574 => (x"64",x"25",x"20",x"74"),
  1575 => (x"75",x"48",x"00",x"0a"),
  1576 => (x"6e",x"69",x"74",x"6e"),
  1577 => (x"6f",x"66",x"20",x"67"),
  1578 => (x"69",x"66",x"20",x"72"),
  1579 => (x"79",x"73",x"65",x"6c"),
  1580 => (x"6d",x"65",x"74",x"73"),
  1581 => (x"41",x"46",x"00",x"0a"),
  1582 => (x"20",x"32",x"33",x"54"),
  1583 => (x"46",x"00",x"20",x"20"),
  1584 => (x"36",x"31",x"54",x"41"),
  1585 => (x"00",x"20",x"20",x"20"),
  1586 => (x"73",x"75",x"6c",x"43"),
  1587 => (x"20",x"72",x"65",x"74"),
  1588 => (x"65",x"7a",x"69",x"73"),
  1589 => (x"64",x"25",x"20",x"3a"),
  1590 => (x"6c",x"43",x"20",x"2c"),
  1591 => (x"65",x"74",x"73",x"75"),
  1592 => (x"61",x"6d",x"20",x"72"),
  1593 => (x"20",x"2c",x"6b",x"73"),
  1594 => (x"00",x"0a",x"64",x"25"),
  1595 => (x"63",x"65",x"68",x"43"),
  1596 => (x"6d",x"75",x"73",x"6b"),
  1597 => (x"67",x"6e",x"69",x"6d"),
  1598 => (x"6f",x"72",x"66",x"20"),
  1599 => (x"64",x"25",x"20",x"6d"),
  1600 => (x"20",x"6f",x"74",x"20"),
  1601 => (x"2e",x"2e",x"64",x"25"),
  1602 => (x"25",x"00",x"20",x"2e"),
  1603 => (x"25",x"00",x"0a",x"64"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
