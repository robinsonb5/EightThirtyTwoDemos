
package Toplevel_Config is
	constant Toplevel_UseSDRAM : boolean := true;
	constant Toplevel_UseUART : boolean := true;
	constant Toplevel_UseVGA : boolean := true;
	constant Toplevel_UseAudio : boolean := true;
end package;
