
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"d7",x"01"),
     1 => (x"58",x"0e",x"87",x"da"),
     2 => (x"27",x"0e",x"59",x"5e"),
     3 => (x"00",x"00",x"00",x"43"),
     4 => (x"26",x"49",x"26",x"0f"),
     5 => (x"26",x"80",x"ff",x"48"),
     6 => (x"26",x"27",x"4f",x"08"),
     7 => (x"4f",x"00",x"00",x"00"),
     8 => (x"00",x"00",x"35",x"27"),
     9 => (x"f8",x"27",x"4f",x"00"),
    10 => (x"4e",x"00",x"00",x"41"),
    11 => (x"00",x"06",x"6f",x"27"),
    12 => (x"fd",x"00",x"0f",x"00"),
    13 => (x"c0",x"f0",x"c1",x"87"),
    14 => (x"00",x"42",x"27",x"4e"),
    15 => (x"00",x"0f",x"00",x"00"),
    16 => (x"4f",x"4f",x"87",x"fd"),
    17 => (x"ff",x"86",x"fc",x"1e"),
    18 => (x"48",x"69",x"49",x"c0"),
    19 => (x"c4",x"98",x"c0",x"c4"),
    20 => (x"02",x"6e",x"58",x"a6"),
    21 => (x"c8",x"87",x"f3",x"ff"),
    22 => (x"66",x"c8",x"79",x"66"),
    23 => (x"26",x"8e",x"fc",x"48"),
    24 => (x"5b",x"5e",x"0e",x"4f"),
    25 => (x"66",x"cc",x"0e",x"5c"),
    26 => (x"13",x"4c",x"c0",x"4b"),
    27 => (x"02",x"9a",x"72",x"4a"),
    28 => (x"72",x"87",x"d9",x"c0"),
    29 => (x"99",x"ff",x"c3",x"49"),
    30 => (x"44",x"27",x"1e",x"71"),
    31 => (x"0f",x"00",x"00",x"00"),
    32 => (x"84",x"c1",x"86",x"c4"),
    33 => (x"9a",x"72",x"4a",x"13"),
    34 => (x"87",x"e7",x"ff",x"05"),
    35 => (x"4c",x"26",x"48",x"74"),
    36 => (x"4f",x"26",x"4b",x"26"),
    37 => (x"5c",x"5b",x"5e",x"0e"),
    38 => (x"66",x"d0",x"0e",x"5d"),
    39 => (x"17",x"40",x"27",x"4a"),
    40 => (x"27",x"4b",x"00",x"00"),
    41 => (x"00",x"00",x"0f",x"88"),
    42 => (x"72",x"4c",x"c0",x"4d"),
    43 => (x"c6",x"c0",x"05",x"9a"),
    44 => (x"53",x"f0",x"c0",x"87"),
    45 => (x"72",x"87",x"f0",x"c0"),
    46 => (x"ea",x"c0",x"02",x"9a"),
    47 => (x"72",x"1e",x"72",x"87"),
    48 => (x"4a",x"66",x"d8",x"49"),
    49 => (x"00",x"05",x"f3",x"27"),
    50 => (x"4a",x"26",x"0f",x"00"),
    51 => (x"53",x"11",x"81",x"75"),
    52 => (x"49",x"72",x"1e",x"71"),
    53 => (x"27",x"4a",x"66",x"d8"),
    54 => (x"00",x"00",x"05",x"f3"),
    55 => (x"26",x"4a",x"70",x"0f"),
    56 => (x"05",x"9a",x"72",x"49"),
    57 => (x"27",x"87",x"d6",x"ff"),
    58 => (x"00",x"00",x"17",x"40"),
    59 => (x"e8",x"c0",x"02",x"ab"),
    60 => (x"4d",x"66",x"d8",x"87"),
    61 => (x"c1",x"1e",x"66",x"dc"),
    62 => (x"49",x"6b",x"97",x"8b"),
    63 => (x"c0",x"c0",x"c0",x"c1"),
    64 => (x"c0",x"c4",x"91",x"c0"),
    65 => (x"71",x"49",x"91",x"b7"),
    66 => (x"c8",x"0f",x"75",x"1e"),
    67 => (x"27",x"84",x"c1",x"86"),
    68 => (x"00",x"00",x"17",x"40"),
    69 => (x"db",x"ff",x"05",x"ab"),
    70 => (x"26",x"48",x"74",x"87"),
    71 => (x"26",x"4c",x"26",x"4d"),
    72 => (x"0e",x"4f",x"26",x"4b"),
    73 => (x"5d",x"5c",x"5b",x"5e"),
    74 => (x"4c",x"66",x"d0",x"0e"),
    75 => (x"4b",x"14",x"4d",x"ff"),
    76 => (x"c0",x"c0",x"c0",x"c1"),
    77 => (x"c0",x"c4",x"93",x"c0"),
    78 => (x"73",x"4b",x"93",x"b7"),
    79 => (x"e5",x"c0",x"02",x"9b"),
    80 => (x"d8",x"85",x"c1",x"87"),
    81 => (x"1e",x"73",x"1e",x"66"),
    82 => (x"c8",x"0f",x"66",x"dc"),
    83 => (x"05",x"a8",x"73",x"86"),
    84 => (x"14",x"87",x"d3",x"c0"),
    85 => (x"c0",x"c0",x"c1",x"4b"),
    86 => (x"c4",x"93",x"c0",x"c0"),
    87 => (x"4b",x"93",x"b7",x"c0"),
    88 => (x"ff",x"05",x"9b",x"73"),
    89 => (x"48",x"75",x"87",x"db"),
    90 => (x"4c",x"26",x"4d",x"26"),
    91 => (x"4f",x"26",x"4b",x"26"),
    92 => (x"5c",x"5b",x"5e",x"0e"),
    93 => (x"86",x"f4",x"0e",x"5d"),
    94 => (x"4b",x"66",x"e4",x"c0"),
    95 => (x"a6",x"c4",x"4c",x"c0"),
    96 => (x"dc",x"78",x"c0",x"48"),
    97 => (x"4d",x"bf",x"97",x"66"),
    98 => (x"c0",x"c0",x"c0",x"c1"),
    99 => (x"c0",x"c4",x"95",x"c0"),
   100 => (x"dc",x"4d",x"95",x"b7"),
   101 => (x"80",x"c1",x"48",x"66"),
   102 => (x"58",x"a6",x"e0",x"c0"),
   103 => (x"c5",x"02",x"9d",x"75"),
   104 => (x"66",x"c4",x"87",x"cc"),
   105 => (x"87",x"ce",x"c4",x"02"),
   106 => (x"c0",x"48",x"a6",x"c8"),
   107 => (x"48",x"a6",x"c4",x"78"),
   108 => (x"49",x"75",x"78",x"c0"),
   109 => (x"02",x"ad",x"f0",x"c0"),
   110 => (x"c1",x"87",x"e8",x"c1"),
   111 => (x"c1",x"02",x"a9",x"e3"),
   112 => (x"e4",x"c1",x"87",x"e9"),
   113 => (x"e6",x"c0",x"02",x"a9"),
   114 => (x"a9",x"ec",x"c1",x"87"),
   115 => (x"87",x"d3",x"c1",x"02"),
   116 => (x"02",x"a9",x"f0",x"c1"),
   117 => (x"c1",x"87",x"e0",x"c0"),
   118 => (x"c0",x"02",x"a9",x"f3"),
   119 => (x"f5",x"c1",x"87",x"e1"),
   120 => (x"ca",x"c0",x"02",x"a9"),
   121 => (x"a9",x"f8",x"c1",x"87"),
   122 => (x"87",x"cb",x"c0",x"02"),
   123 => (x"c8",x"87",x"db",x"c1"),
   124 => (x"78",x"ca",x"48",x"a6"),
   125 => (x"c8",x"87",x"ea",x"c1"),
   126 => (x"78",x"d0",x"48",x"a6"),
   127 => (x"c0",x"87",x"e2",x"c1"),
   128 => (x"73",x"1e",x"66",x"e8"),
   129 => (x"66",x"e8",x"c0",x"1e"),
   130 => (x"c0",x"80",x"c4",x"48"),
   131 => (x"c0",x"58",x"a6",x"ec"),
   132 => (x"c4",x"49",x"66",x"e8"),
   133 => (x"fc",x"1e",x"69",x"89"),
   134 => (x"86",x"cc",x"87",x"c9"),
   135 => (x"84",x"71",x"49",x"70"),
   136 => (x"c4",x"87",x"fe",x"c0"),
   137 => (x"78",x"c1",x"48",x"a6"),
   138 => (x"c0",x"87",x"f6",x"c0"),
   139 => (x"c0",x"1e",x"66",x"e8"),
   140 => (x"c4",x"48",x"66",x"e4"),
   141 => (x"a6",x"e8",x"c0",x"80"),
   142 => (x"66",x"e4",x"c0",x"58"),
   143 => (x"69",x"89",x"c4",x"49"),
   144 => (x"c8",x"0f",x"73",x"1e"),
   145 => (x"c0",x"84",x"c1",x"86"),
   146 => (x"e8",x"c0",x"87",x"d7"),
   147 => (x"e5",x"c0",x"1e",x"66"),
   148 => (x"c8",x"0f",x"73",x"1e"),
   149 => (x"66",x"e8",x"c0",x"86"),
   150 => (x"73",x"1e",x"75",x"1e"),
   151 => (x"c1",x"86",x"c8",x"0f"),
   152 => (x"02",x"66",x"c8",x"84"),
   153 => (x"c0",x"87",x"e8",x"c1"),
   154 => (x"c4",x"48",x"66",x"e0"),
   155 => (x"a6",x"e4",x"c0",x"80"),
   156 => (x"66",x"e0",x"c0",x"58"),
   157 => (x"76",x"89",x"c4",x"49"),
   158 => (x"c1",x"78",x"69",x"48"),
   159 => (x"c0",x"05",x"ad",x"e4"),
   160 => (x"48",x"6e",x"87",x"dc"),
   161 => (x"03",x"a8",x"b7",x"c0"),
   162 => (x"c0",x"87",x"d3",x"c0"),
   163 => (x"44",x"27",x"1e",x"ed"),
   164 => (x"0f",x"00",x"00",x"00"),
   165 => (x"48",x"6e",x"86",x"c4"),
   166 => (x"c4",x"88",x"08",x"c0"),
   167 => (x"e8",x"c0",x"58",x"a6"),
   168 => (x"1e",x"73",x"1e",x"66"),
   169 => (x"cc",x"1e",x"66",x"d0"),
   170 => (x"e7",x"f7",x"1e",x"66"),
   171 => (x"70",x"86",x"d0",x"87"),
   172 => (x"c0",x"84",x"71",x"49"),
   173 => (x"e5",x"c0",x"87",x"d9"),
   174 => (x"c8",x"c0",x"05",x"ad"),
   175 => (x"48",x"a6",x"c4",x"87"),
   176 => (x"ca",x"c0",x"78",x"c1"),
   177 => (x"66",x"e8",x"c0",x"87"),
   178 => (x"73",x"1e",x"75",x"1e"),
   179 => (x"dc",x"86",x"c8",x"0f"),
   180 => (x"4d",x"bf",x"97",x"66"),
   181 => (x"c0",x"c0",x"c0",x"c1"),
   182 => (x"c0",x"c4",x"95",x"c0"),
   183 => (x"dc",x"4d",x"95",x"b7"),
   184 => (x"80",x"c1",x"48",x"66"),
   185 => (x"58",x"a6",x"e0",x"c0"),
   186 => (x"fa",x"05",x"9d",x"75"),
   187 => (x"48",x"74",x"87",x"f4"),
   188 => (x"4d",x"26",x"8e",x"f4"),
   189 => (x"4b",x"26",x"4c",x"26"),
   190 => (x"c0",x"1e",x"4f",x"26"),
   191 => (x"00",x"44",x"27",x"1e"),
   192 => (x"d0",x"1e",x"00",x"00"),
   193 => (x"66",x"d0",x"1e",x"66"),
   194 => (x"01",x"70",x"27",x"1e"),
   195 => (x"d0",x"0f",x"00",x"00"),
   196 => (x"1e",x"4f",x"26",x"86"),
   197 => (x"44",x"27",x"1e",x"c0"),
   198 => (x"1e",x"00",x"00",x"00"),
   199 => (x"d0",x"1e",x"a6",x"d0"),
   200 => (x"70",x"27",x"1e",x"66"),
   201 => (x"0f",x"00",x"00",x"01"),
   202 => (x"4f",x"26",x"86",x"d0"),
   203 => (x"4a",x"66",x"c8",x"1e"),
   204 => (x"c4",x"49",x"66",x"c8"),
   205 => (x"c0",x"02",x"69",x"81"),
   206 => (x"49",x"72",x"87",x"dc"),
   207 => (x"48",x"69",x"81",x"c4"),
   208 => (x"79",x"70",x"88",x"c1"),
   209 => (x"48",x"71",x"49",x"6a"),
   210 => (x"7a",x"70",x"80",x"c1"),
   211 => (x"51",x"66",x"c4",x"97"),
   212 => (x"c0",x"48",x"66",x"c4"),
   213 => (x"48",x"c0",x"87",x"c2"),
   214 => (x"f8",x"1e",x"4f",x"26"),
   215 => (x"cc",x"48",x"76",x"86"),
   216 => (x"a6",x"c4",x"78",x"66"),
   217 => (x"76",x"78",x"ff",x"48"),
   218 => (x"03",x"2c",x"27",x"1e"),
   219 => (x"dc",x"1e",x"00",x"00"),
   220 => (x"66",x"dc",x"1e",x"a6"),
   221 => (x"01",x"70",x"27",x"1e"),
   222 => (x"d0",x"0f",x"00",x"00"),
   223 => (x"26",x"8e",x"f8",x"86"),
   224 => (x"86",x"f8",x"1e",x"4f"),
   225 => (x"66",x"cc",x"48",x"76"),
   226 => (x"48",x"a6",x"c4",x"78"),
   227 => (x"76",x"78",x"66",x"d0"),
   228 => (x"03",x"2c",x"27",x"1e"),
   229 => (x"c0",x"1e",x"00",x"00"),
   230 => (x"c0",x"1e",x"a6",x"e0"),
   231 => (x"27",x"1e",x"66",x"e0"),
   232 => (x"00",x"00",x"01",x"70"),
   233 => (x"f8",x"86",x"d0",x"0f"),
   234 => (x"1e",x"4f",x"26",x"8e"),
   235 => (x"48",x"76",x"86",x"f8"),
   236 => (x"c4",x"78",x"66",x"cc"),
   237 => (x"78",x"ff",x"48",x"a6"),
   238 => (x"2c",x"27",x"1e",x"76"),
   239 => (x"1e",x"00",x"00",x"03"),
   240 => (x"dc",x"1e",x"66",x"dc"),
   241 => (x"70",x"27",x"1e",x"66"),
   242 => (x"0f",x"00",x"00",x"01"),
   243 => (x"8e",x"f8",x"86",x"d0"),
   244 => (x"73",x"1e",x"4f",x"26"),
   245 => (x"4b",x"66",x"cc",x"1e"),
   246 => (x"c8",x"7b",x"66",x"c8"),
   247 => (x"e0",x"27",x"1e",x"66"),
   248 => (x"0f",x"00",x"00",x"05"),
   249 => (x"98",x"70",x"86",x"c4"),
   250 => (x"87",x"c2",x"c0",x"05"),
   251 => (x"66",x"c8",x"7b",x"c3"),
   252 => (x"48",x"66",x"c8",x"49"),
   253 => (x"c0",x"02",x"a8",x"c0"),
   254 => (x"a9",x"c1",x"87",x"db"),
   255 => (x"87",x"da",x"c0",x"02"),
   256 => (x"c0",x"02",x"a9",x"c2"),
   257 => (x"a9",x"c3",x"87",x"ed"),
   258 => (x"87",x"ee",x"c0",x"02"),
   259 => (x"c0",x"02",x"a9",x"c4"),
   260 => (x"e5",x"c0",x"87",x"e6"),
   261 => (x"c0",x"7b",x"c0",x"87"),
   262 => (x"58",x"27",x"87",x"e0"),
   263 => (x"bf",x"00",x"00",x"17"),
   264 => (x"b7",x"e4",x"c1",x"48"),
   265 => (x"c5",x"c0",x"06",x"a8"),
   266 => (x"c0",x"7b",x"c0",x"87"),
   267 => (x"7b",x"c3",x"87",x"cc"),
   268 => (x"c1",x"87",x"c7",x"c0"),
   269 => (x"87",x"c2",x"c0",x"7b"),
   270 => (x"4b",x"26",x"7b",x"c2"),
   271 => (x"c4",x"1e",x"4f",x"26"),
   272 => (x"81",x"c2",x"49",x"66"),
   273 => (x"71",x"48",x"66",x"c8"),
   274 => (x"08",x"66",x"cc",x"80"),
   275 => (x"4f",x"26",x"08",x"78"),
   276 => (x"5c",x"5b",x"5e",x"0e"),
   277 => (x"66",x"d8",x"0e",x"5d"),
   278 => (x"74",x"84",x"c5",x"4c"),
   279 => (x"d0",x"93",x"c4",x"4b"),
   280 => (x"66",x"dc",x"83",x"66"),
   281 => (x"c1",x"49",x"74",x"7b"),
   282 => (x"c4",x"4a",x"71",x"81"),
   283 => (x"82",x"66",x"d0",x"92"),
   284 => (x"4a",x"74",x"7a",x"6b"),
   285 => (x"92",x"c4",x"82",x"de"),
   286 => (x"74",x"82",x"66",x"d0"),
   287 => (x"71",x"4d",x"74",x"7a"),
   288 => (x"c0",x"01",x"ac",x"b7"),
   289 => (x"4a",x"74",x"87",x"dd"),
   290 => (x"d4",x"92",x"c8",x"c3"),
   291 => (x"49",x"75",x"82",x"66"),
   292 => (x"81",x"72",x"91",x"c4"),
   293 => (x"85",x"c1",x"79",x"74"),
   294 => (x"81",x"c1",x"49",x"74"),
   295 => (x"06",x"ad",x"b7",x"71"),
   296 => (x"74",x"87",x"e3",x"ff"),
   297 => (x"92",x"c8",x"c3",x"4a"),
   298 => (x"74",x"82",x"66",x"d4"),
   299 => (x"c4",x"89",x"c1",x"49"),
   300 => (x"69",x"81",x"72",x"91"),
   301 => (x"70",x"80",x"c1",x"48"),
   302 => (x"c4",x"49",x"74",x"79"),
   303 => (x"4a",x"66",x"d0",x"91"),
   304 => (x"4b",x"74",x"82",x"71"),
   305 => (x"c8",x"c3",x"83",x"d4"),
   306 => (x"83",x"66",x"d4",x"93"),
   307 => (x"79",x"6a",x"81",x"73"),
   308 => (x"00",x"17",x"58",x"27"),
   309 => (x"78",x"c5",x"48",x"00"),
   310 => (x"4c",x"26",x"4d",x"26"),
   311 => (x"4f",x"26",x"4b",x"26"),
   312 => (x"0e",x"5b",x"5e",x"0e"),
   313 => (x"4b",x"66",x"c8",x"97"),
   314 => (x"c0",x"c1",x"4a",x"73"),
   315 => (x"92",x"c0",x"c0",x"c0"),
   316 => (x"92",x"b7",x"c0",x"c4"),
   317 => (x"66",x"cc",x"97",x"4a"),
   318 => (x"c0",x"c0",x"c1",x"49"),
   319 => (x"c4",x"91",x"c0",x"c0"),
   320 => (x"49",x"91",x"b7",x"c0"),
   321 => (x"02",x"aa",x"b7",x"71"),
   322 => (x"c0",x"87",x"c5",x"c0"),
   323 => (x"87",x"c9",x"c0",x"48"),
   324 => (x"00",x"17",x"64",x"27"),
   325 => (x"c1",x"5b",x"97",x"00"),
   326 => (x"26",x"4b",x"26",x"48"),
   327 => (x"5b",x"5e",x"0e",x"4f"),
   328 => (x"86",x"fc",x"0e",x"5c"),
   329 => (x"c2",x"4c",x"6e",x"97"),
   330 => (x"49",x"66",x"d4",x"4b"),
   331 => (x"81",x"73",x"81",x"c1"),
   332 => (x"c1",x"49",x"69",x"97"),
   333 => (x"c0",x"c0",x"c0",x"c0"),
   334 => (x"b7",x"c0",x"c4",x"91"),
   335 => (x"1e",x"71",x"49",x"91"),
   336 => (x"73",x"49",x"66",x"d4"),
   337 => (x"49",x"69",x"97",x"81"),
   338 => (x"c0",x"c0",x"c0",x"c1"),
   339 => (x"c0",x"c4",x"91",x"c0"),
   340 => (x"71",x"49",x"91",x"b7"),
   341 => (x"04",x"e0",x"27",x"1e"),
   342 => (x"c8",x"0f",x"00",x"00"),
   343 => (x"05",x"98",x"70",x"86"),
   344 => (x"c1",x"87",x"c5",x"c0"),
   345 => (x"83",x"c1",x"4c",x"c1"),
   346 => (x"06",x"ab",x"b7",x"c2"),
   347 => (x"74",x"87",x"fa",x"fe"),
   348 => (x"c0",x"c0",x"c1",x"49"),
   349 => (x"c4",x"91",x"c0",x"c0"),
   350 => (x"49",x"91",x"b7",x"c0"),
   351 => (x"a9",x"b7",x"d7",x"c1"),
   352 => (x"87",x"d7",x"c0",x"04"),
   353 => (x"c0",x"c1",x"49",x"74"),
   354 => (x"91",x"c0",x"c0",x"c0"),
   355 => (x"91",x"b7",x"c0",x"c4"),
   356 => (x"b7",x"da",x"c1",x"49"),
   357 => (x"c2",x"c0",x"03",x"a9"),
   358 => (x"74",x"4b",x"c7",x"87"),
   359 => (x"c0",x"c0",x"c1",x"49"),
   360 => (x"c4",x"91",x"c0",x"c0"),
   361 => (x"49",x"91",x"b7",x"c0"),
   362 => (x"05",x"a9",x"d2",x"c1"),
   363 => (x"c1",x"87",x"c5",x"c0"),
   364 => (x"87",x"e4",x"c0",x"48"),
   365 => (x"d4",x"4a",x"66",x"d0"),
   366 => (x"57",x"27",x"49",x"66"),
   367 => (x"0f",x"00",x"00",x"06"),
   368 => (x"06",x"a8",x"b7",x"c0"),
   369 => (x"73",x"87",x"cf",x"c0"),
   370 => (x"27",x"80",x"c7",x"48"),
   371 => (x"00",x"00",x"17",x"5c"),
   372 => (x"c0",x"48",x"c1",x"58"),
   373 => (x"48",x"c0",x"87",x"c2"),
   374 => (x"4c",x"26",x"8e",x"fc"),
   375 => (x"4f",x"26",x"4b",x"26"),
   376 => (x"48",x"66",x"c4",x"1e"),
   377 => (x"c0",x"05",x"a8",x"c2"),
   378 => (x"48",x"c1",x"87",x"c5"),
   379 => (x"c0",x"87",x"c2",x"c0"),
   380 => (x"1e",x"4f",x"26",x"48"),
   381 => (x"9a",x"72",x"1e",x"73"),
   382 => (x"c0",x"87",x"e7",x"02"),
   383 => (x"72",x"4b",x"c1",x"48"),
   384 => (x"87",x"d1",x"06",x"a9"),
   385 => (x"c9",x"06",x"82",x"72"),
   386 => (x"72",x"83",x"73",x"87"),
   387 => (x"87",x"f4",x"01",x"a9"),
   388 => (x"b2",x"c1",x"87",x"c3"),
   389 => (x"03",x"a9",x"72",x"3a"),
   390 => (x"07",x"80",x"73",x"89"),
   391 => (x"05",x"2b",x"2a",x"c1"),
   392 => (x"4b",x"26",x"87",x"f3"),
   393 => (x"75",x"1e",x"4f",x"26"),
   394 => (x"71",x"4d",x"c4",x"1e"),
   395 => (x"ff",x"04",x"a1",x"b7"),
   396 => (x"c3",x"81",x"c1",x"b9"),
   397 => (x"b7",x"72",x"07",x"bd"),
   398 => (x"ba",x"ff",x"04",x"a2"),
   399 => (x"bd",x"c1",x"82",x"c1"),
   400 => (x"87",x"ef",x"fe",x"07"),
   401 => (x"ff",x"04",x"2d",x"c1"),
   402 => (x"07",x"80",x"c1",x"b8"),
   403 => (x"b9",x"ff",x"04",x"2d"),
   404 => (x"26",x"07",x"81",x"c1"),
   405 => (x"1e",x"4f",x"26",x"4d"),
   406 => (x"48",x"12",x"1e",x"72"),
   407 => (x"87",x"c4",x"02",x"11"),
   408 => (x"87",x"f6",x"02",x"88"),
   409 => (x"4f",x"26",x"4a",x"26"),
   410 => (x"bf",x"c8",x"ff",x"1e"),
   411 => (x"0e",x"4f",x"26",x"48"),
   412 => (x"5d",x"5c",x"5b",x"5e"),
   413 => (x"c4",x"86",x"f0",x"0e"),
   414 => (x"54",x"27",x"4b",x"66"),
   415 => (x"48",x"00",x"00",x"17"),
   416 => (x"00",x"3f",x"58",x"27"),
   417 => (x"50",x"27",x"78",x"00"),
   418 => (x"48",x"00",x"00",x"17"),
   419 => (x"00",x"3f",x"88",x"27"),
   420 => (x"88",x"27",x"78",x"00"),
   421 => (x"48",x"00",x"00",x"3f"),
   422 => (x"00",x"3f",x"58",x"27"),
   423 => (x"8c",x"27",x"78",x"00"),
   424 => (x"48",x"00",x"00",x"3f"),
   425 => (x"90",x"27",x"78",x"c0"),
   426 => (x"48",x"00",x"00",x"3f"),
   427 => (x"94",x"27",x"78",x"c2"),
   428 => (x"48",x"00",x"00",x"3f"),
   429 => (x"27",x"78",x"e8",x"c0"),
   430 => (x"00",x"00",x"3f",x"98"),
   431 => (x"11",x"12",x"27",x"4a"),
   432 => (x"20",x"48",x"00",x"00"),
   433 => (x"20",x"42",x"20",x"42"),
   434 => (x"20",x"42",x"20",x"42"),
   435 => (x"20",x"42",x"20",x"42"),
   436 => (x"10",x"52",x"10",x"42"),
   437 => (x"27",x"52",x"10",x"52"),
   438 => (x"00",x"00",x"3f",x"b8"),
   439 => (x"11",x"31",x"27",x"4a"),
   440 => (x"20",x"48",x"00",x"00"),
   441 => (x"20",x"42",x"20",x"42"),
   442 => (x"20",x"42",x"20",x"42"),
   443 => (x"20",x"42",x"20",x"42"),
   444 => (x"10",x"52",x"10",x"42"),
   445 => (x"27",x"52",x"10",x"52"),
   446 => (x"00",x"00",x"1e",x"8c"),
   447 => (x"27",x"78",x"ca",x"48"),
   448 => (x"00",x"00",x"11",x"50"),
   449 => (x"03",x"13",x"27",x"1e"),
   450 => (x"c4",x"0f",x"00",x"00"),
   451 => (x"11",x"52",x"27",x"86"),
   452 => (x"27",x"1e",x"00",x"00"),
   453 => (x"00",x"00",x"03",x"13"),
   454 => (x"27",x"86",x"c4",x"0f"),
   455 => (x"00",x"00",x"11",x"82"),
   456 => (x"03",x"13",x"27",x"1e"),
   457 => (x"c4",x"0f",x"00",x"00"),
   458 => (x"17",x"38",x"27",x"86"),
   459 => (x"02",x"bf",x"00",x"00"),
   460 => (x"27",x"87",x"df",x"c0"),
   461 => (x"00",x"00",x"0f",x"99"),
   462 => (x"03",x"13",x"27",x"1e"),
   463 => (x"c4",x"0f",x"00",x"00"),
   464 => (x"0f",x"c5",x"27",x"86"),
   465 => (x"27",x"1e",x"00",x"00"),
   466 => (x"00",x"00",x"03",x"13"),
   467 => (x"c0",x"86",x"c4",x"0f"),
   468 => (x"c7",x"27",x"87",x"dc"),
   469 => (x"1e",x"00",x"00",x"0f"),
   470 => (x"00",x"03",x"13",x"27"),
   471 => (x"86",x"c4",x"0f",x"00"),
   472 => (x"00",x"0f",x"f6",x"27"),
   473 => (x"13",x"27",x"1e",x"00"),
   474 => (x"0f",x"00",x"00",x"03"),
   475 => (x"3c",x"27",x"86",x"c4"),
   476 => (x"bf",x"00",x"00",x"17"),
   477 => (x"11",x"84",x"27",x"1e"),
   478 => (x"27",x"1e",x"00",x"00"),
   479 => (x"00",x"00",x"03",x"13"),
   480 => (x"27",x"86",x"c8",x"0f"),
   481 => (x"00",x"00",x"06",x"68"),
   482 => (x"3f",x"44",x"27",x"0f"),
   483 => (x"c1",x"58",x"00",x"00"),
   484 => (x"17",x"3c",x"27",x"4c"),
   485 => (x"48",x"bf",x"00",x"00"),
   486 => (x"06",x"a8",x"b7",x"c0"),
   487 => (x"27",x"87",x"cf",x"c6"),
   488 => (x"00",x"00",x"0f",x"72"),
   489 => (x"0f",x"36",x"27",x"0f"),
   490 => (x"76",x"0f",x"00",x"00"),
   491 => (x"c3",x"78",x"c2",x"48"),
   492 => (x"3f",x"d8",x"27",x"4b"),
   493 => (x"27",x"4a",x"00",x"00"),
   494 => (x"00",x"00",x"10",x"17"),
   495 => (x"20",x"42",x"20",x"48"),
   496 => (x"20",x"42",x"20",x"42"),
   497 => (x"20",x"42",x"20",x"42"),
   498 => (x"10",x"42",x"20",x"42"),
   499 => (x"10",x"52",x"10",x"52"),
   500 => (x"48",x"a6",x"c8",x"52"),
   501 => (x"d8",x"27",x"78",x"c1"),
   502 => (x"1e",x"00",x"00",x"3f"),
   503 => (x"00",x"3f",x"b8",x"27"),
   504 => (x"1d",x"27",x"1e",x"00"),
   505 => (x"0f",x"00",x"00",x"05"),
   506 => (x"98",x"70",x"86",x"c8"),
   507 => (x"87",x"c5",x"c0",x"05"),
   508 => (x"c2",x"c0",x"49",x"c1"),
   509 => (x"27",x"49",x"c0",x"87"),
   510 => (x"00",x"00",x"17",x"60"),
   511 => (x"ab",x"b7",x"6e",x"59"),
   512 => (x"87",x"e9",x"c0",x"06"),
   513 => (x"91",x"c5",x"49",x"6e"),
   514 => (x"88",x"73",x"48",x"71"),
   515 => (x"cc",x"58",x"a6",x"d0"),
   516 => (x"1e",x"73",x"1e",x"a6"),
   517 => (x"27",x"1e",x"66",x"c8"),
   518 => (x"00",x"00",x"04",x"3e"),
   519 => (x"6e",x"86",x"cc",x"0f"),
   520 => (x"c4",x"80",x"c1",x"48"),
   521 => (x"b7",x"6e",x"58",x"a6"),
   522 => (x"d7",x"ff",x"01",x"ab"),
   523 => (x"1e",x"66",x"cc",x"87"),
   524 => (x"27",x"1e",x"66",x"c4"),
   525 => (x"00",x"00",x"18",x"30"),
   526 => (x"17",x"68",x"27",x"1e"),
   527 => (x"27",x"1e",x"00",x"00"),
   528 => (x"00",x"00",x"04",x"50"),
   529 => (x"27",x"86",x"d0",x"0f"),
   530 => (x"00",x"00",x"17",x"50"),
   531 => (x"20",x"27",x"1e",x"bf"),
   532 => (x"0f",x"00",x"00",x"0e"),
   533 => (x"c1",x"c1",x"86",x"c4"),
   534 => (x"17",x"61",x"27",x"4d"),
   535 => (x"bf",x"97",x"00",x"00"),
   536 => (x"c0",x"c0",x"c1",x"49"),
   537 => (x"c4",x"91",x"c0",x"c0"),
   538 => (x"49",x"91",x"b7",x"c0"),
   539 => (x"a9",x"b7",x"c1",x"c1"),
   540 => (x"87",x"ff",x"c1",x"04"),
   541 => (x"75",x"1e",x"c3",x"c1"),
   542 => (x"c0",x"c0",x"c1",x"49"),
   543 => (x"c4",x"91",x"c0",x"c0"),
   544 => (x"49",x"91",x"b7",x"c0"),
   545 => (x"e0",x"27",x"1e",x"71"),
   546 => (x"0f",x"00",x"00",x"04"),
   547 => (x"66",x"c8",x"86",x"c8"),
   548 => (x"f5",x"c0",x"05",x"a8"),
   549 => (x"1e",x"a6",x"c8",x"87"),
   550 => (x"d2",x"27",x"1e",x"c0"),
   551 => (x"0f",x"00",x"00",x"03"),
   552 => (x"d8",x"27",x"86",x"c8"),
   553 => (x"4a",x"00",x"00",x"3f"),
   554 => (x"00",x"0f",x"f8",x"27"),
   555 => (x"42",x"20",x"48",x"00"),
   556 => (x"42",x"20",x"42",x"20"),
   557 => (x"42",x"20",x"42",x"20"),
   558 => (x"42",x"20",x"42",x"20"),
   559 => (x"52",x"10",x"52",x"10"),
   560 => (x"4b",x"74",x"52",x"10"),
   561 => (x"00",x"17",x"5c",x"27"),
   562 => (x"85",x"c1",x"5c",x"00"),
   563 => (x"c0",x"c1",x"4a",x"75"),
   564 => (x"92",x"c0",x"c0",x"c0"),
   565 => (x"92",x"b7",x"c0",x"c4"),
   566 => (x"17",x"61",x"27",x"4a"),
   567 => (x"bf",x"97",x"00",x"00"),
   568 => (x"c0",x"c0",x"c1",x"49"),
   569 => (x"c4",x"91",x"c0",x"c0"),
   570 => (x"49",x"91",x"b7",x"c0"),
   571 => (x"06",x"aa",x"b7",x"71"),
   572 => (x"6e",x"87",x"c1",x"fe"),
   573 => (x"72",x"1e",x"71",x"93"),
   574 => (x"d4",x"49",x"73",x"1e"),
   575 => (x"26",x"27",x"4a",x"66"),
   576 => (x"0f",x"00",x"00",x"06"),
   577 => (x"49",x"26",x"4a",x"26"),
   578 => (x"73",x"58",x"a6",x"c4"),
   579 => (x"89",x"66",x"cc",x"49"),
   580 => (x"4b",x"71",x"91",x"c7"),
   581 => (x"1e",x"76",x"8b",x"6e"),
   582 => (x"00",x"0e",x"af",x"27"),
   583 => (x"86",x"c4",x"0f",x"00"),
   584 => (x"3c",x"27",x"84",x"c1"),
   585 => (x"bf",x"00",x"00",x"17"),
   586 => (x"f9",x"06",x"ac",x"b7"),
   587 => (x"68",x"27",x"87",x"f1"),
   588 => (x"0f",x"00",x"00",x"06"),
   589 => (x"00",x"3f",x"48",x"27"),
   590 => (x"b1",x"27",x"58",x"00"),
   591 => (x"1e",x"00",x"00",x"11"),
   592 => (x"00",x"03",x"13",x"27"),
   593 => (x"86",x"c4",x"0f",x"00"),
   594 => (x"00",x"11",x"c1",x"27"),
   595 => (x"13",x"27",x"1e",x"00"),
   596 => (x"0f",x"00",x"00",x"03"),
   597 => (x"c3",x"27",x"86",x"c4"),
   598 => (x"1e",x"00",x"00",x"11"),
   599 => (x"00",x"03",x"13",x"27"),
   600 => (x"86",x"c4",x"0f",x"00"),
   601 => (x"00",x"11",x"f9",x"27"),
   602 => (x"13",x"27",x"1e",x"00"),
   603 => (x"0f",x"00",x"00",x"03"),
   604 => (x"58",x"27",x"86",x"c4"),
   605 => (x"bf",x"00",x"00",x"17"),
   606 => (x"11",x"fb",x"27",x"1e"),
   607 => (x"27",x"1e",x"00",x"00"),
   608 => (x"00",x"00",x"03",x"13"),
   609 => (x"c5",x"86",x"c8",x"0f"),
   610 => (x"12",x"14",x"27",x"1e"),
   611 => (x"27",x"1e",x"00",x"00"),
   612 => (x"00",x"00",x"03",x"13"),
   613 => (x"27",x"86",x"c8",x"0f"),
   614 => (x"00",x"00",x"17",x"5c"),
   615 => (x"2d",x"27",x"1e",x"bf"),
   616 => (x"1e",x"00",x"00",x"12"),
   617 => (x"00",x"03",x"13",x"27"),
   618 => (x"86",x"c8",x"0f",x"00"),
   619 => (x"46",x"27",x"1e",x"c1"),
   620 => (x"1e",x"00",x"00",x"12"),
   621 => (x"00",x"03",x"13",x"27"),
   622 => (x"86",x"c8",x"0f",x"00"),
   623 => (x"00",x"17",x"60",x"27"),
   624 => (x"49",x"bf",x"97",x"00"),
   625 => (x"c0",x"c0",x"c0",x"c1"),
   626 => (x"c0",x"c4",x"91",x"c0"),
   627 => (x"71",x"49",x"91",x"b7"),
   628 => (x"12",x"5f",x"27",x"1e"),
   629 => (x"27",x"1e",x"00",x"00"),
   630 => (x"00",x"00",x"03",x"13"),
   631 => (x"c1",x"86",x"c8",x"0f"),
   632 => (x"78",x"27",x"1e",x"c1"),
   633 => (x"1e",x"00",x"00",x"12"),
   634 => (x"00",x"03",x"13",x"27"),
   635 => (x"86",x"c8",x"0f",x"00"),
   636 => (x"00",x"17",x"61",x"27"),
   637 => (x"49",x"bf",x"97",x"00"),
   638 => (x"c0",x"c0",x"c0",x"c1"),
   639 => (x"c0",x"c4",x"91",x"c0"),
   640 => (x"71",x"49",x"91",x"b7"),
   641 => (x"12",x"91",x"27",x"1e"),
   642 => (x"27",x"1e",x"00",x"00"),
   643 => (x"00",x"00",x"03",x"13"),
   644 => (x"c1",x"86",x"c8",x"0f"),
   645 => (x"aa",x"27",x"1e",x"c2"),
   646 => (x"1e",x"00",x"00",x"12"),
   647 => (x"00",x"03",x"13",x"27"),
   648 => (x"86",x"c8",x"0f",x"00"),
   649 => (x"00",x"17",x"88",x"27"),
   650 => (x"27",x"1e",x"bf",x"00"),
   651 => (x"00",x"00",x"12",x"c3"),
   652 => (x"03",x"13",x"27",x"1e"),
   653 => (x"c8",x"0f",x"00",x"00"),
   654 => (x"27",x"1e",x"c7",x"86"),
   655 => (x"00",x"00",x"12",x"dc"),
   656 => (x"03",x"13",x"27",x"1e"),
   657 => (x"c8",x"0f",x"00",x"00"),
   658 => (x"1e",x"8c",x"27",x"86"),
   659 => (x"1e",x"bf",x"00",x"00"),
   660 => (x"00",x"12",x"f5",x"27"),
   661 => (x"13",x"27",x"1e",x"00"),
   662 => (x"0f",x"00",x"00",x"03"),
   663 => (x"0e",x"27",x"86",x"c8"),
   664 => (x"1e",x"00",x"00",x"13"),
   665 => (x"00",x"03",x"13",x"27"),
   666 => (x"86",x"c4",x"0f",x"00"),
   667 => (x"00",x"13",x"38",x"27"),
   668 => (x"13",x"27",x"1e",x"00"),
   669 => (x"0f",x"00",x"00",x"03"),
   670 => (x"50",x"27",x"86",x"c4"),
   671 => (x"bf",x"00",x"00",x"17"),
   672 => (x"44",x"27",x"1e",x"bf"),
   673 => (x"1e",x"00",x"00",x"13"),
   674 => (x"00",x"03",x"13",x"27"),
   675 => (x"86",x"c8",x"0f",x"00"),
   676 => (x"00",x"13",x"5d",x"27"),
   677 => (x"13",x"27",x"1e",x"00"),
   678 => (x"0f",x"00",x"00",x"03"),
   679 => (x"50",x"27",x"86",x"c4"),
   680 => (x"bf",x"00",x"00",x"17"),
   681 => (x"69",x"81",x"c4",x"49"),
   682 => (x"13",x"8e",x"27",x"1e"),
   683 => (x"27",x"1e",x"00",x"00"),
   684 => (x"00",x"00",x"03",x"13"),
   685 => (x"c0",x"86",x"c8",x"0f"),
   686 => (x"13",x"a7",x"27",x"1e"),
   687 => (x"27",x"1e",x"00",x"00"),
   688 => (x"00",x"00",x"03",x"13"),
   689 => (x"27",x"86",x"c8",x"0f"),
   690 => (x"00",x"00",x"17",x"50"),
   691 => (x"81",x"c8",x"49",x"bf"),
   692 => (x"c0",x"27",x"1e",x"69"),
   693 => (x"1e",x"00",x"00",x"13"),
   694 => (x"00",x"03",x"13",x"27"),
   695 => (x"86",x"c8",x"0f",x"00"),
   696 => (x"d9",x"27",x"1e",x"c2"),
   697 => (x"1e",x"00",x"00",x"13"),
   698 => (x"00",x"03",x"13",x"27"),
   699 => (x"86",x"c8",x"0f",x"00"),
   700 => (x"00",x"17",x"50",x"27"),
   701 => (x"cc",x"49",x"bf",x"00"),
   702 => (x"27",x"1e",x"69",x"81"),
   703 => (x"00",x"00",x"13",x"f2"),
   704 => (x"03",x"13",x"27",x"1e"),
   705 => (x"c8",x"0f",x"00",x"00"),
   706 => (x"27",x"1e",x"d1",x"86"),
   707 => (x"00",x"00",x"14",x"0b"),
   708 => (x"03",x"13",x"27",x"1e"),
   709 => (x"c8",x"0f",x"00",x"00"),
   710 => (x"17",x"50",x"27",x"86"),
   711 => (x"49",x"bf",x"00",x"00"),
   712 => (x"1e",x"71",x"81",x"d0"),
   713 => (x"00",x"14",x"24",x"27"),
   714 => (x"13",x"27",x"1e",x"00"),
   715 => (x"0f",x"00",x"00",x"03"),
   716 => (x"3d",x"27",x"86",x"c8"),
   717 => (x"1e",x"00",x"00",x"14"),
   718 => (x"00",x"03",x"13",x"27"),
   719 => (x"86",x"c4",x"0f",x"00"),
   720 => (x"00",x"14",x"72",x"27"),
   721 => (x"13",x"27",x"1e",x"00"),
   722 => (x"0f",x"00",x"00",x"03"),
   723 => (x"54",x"27",x"86",x"c4"),
   724 => (x"bf",x"00",x"00",x"17"),
   725 => (x"83",x"27",x"1e",x"bf"),
   726 => (x"1e",x"00",x"00",x"14"),
   727 => (x"00",x"03",x"13",x"27"),
   728 => (x"86",x"c8",x"0f",x"00"),
   729 => (x"00",x"14",x"9c",x"27"),
   730 => (x"13",x"27",x"1e",x"00"),
   731 => (x"0f",x"00",x"00",x"03"),
   732 => (x"54",x"27",x"86",x"c4"),
   733 => (x"bf",x"00",x"00",x"17"),
   734 => (x"69",x"81",x"c4",x"49"),
   735 => (x"14",x"dc",x"27",x"1e"),
   736 => (x"27",x"1e",x"00",x"00"),
   737 => (x"00",x"00",x"03",x"13"),
   738 => (x"c0",x"86",x"c8",x"0f"),
   739 => (x"14",x"f5",x"27",x"1e"),
   740 => (x"27",x"1e",x"00",x"00"),
   741 => (x"00",x"00",x"03",x"13"),
   742 => (x"27",x"86",x"c8",x"0f"),
   743 => (x"00",x"00",x"17",x"54"),
   744 => (x"81",x"c8",x"49",x"bf"),
   745 => (x"0e",x"27",x"1e",x"69"),
   746 => (x"1e",x"00",x"00",x"15"),
   747 => (x"00",x"03",x"13",x"27"),
   748 => (x"86",x"c8",x"0f",x"00"),
   749 => (x"27",x"27",x"1e",x"c1"),
   750 => (x"1e",x"00",x"00",x"15"),
   751 => (x"00",x"03",x"13",x"27"),
   752 => (x"86",x"c8",x"0f",x"00"),
   753 => (x"00",x"17",x"54",x"27"),
   754 => (x"cc",x"49",x"bf",x"00"),
   755 => (x"27",x"1e",x"69",x"81"),
   756 => (x"00",x"00",x"15",x"40"),
   757 => (x"03",x"13",x"27",x"1e"),
   758 => (x"c8",x"0f",x"00",x"00"),
   759 => (x"27",x"1e",x"d2",x"86"),
   760 => (x"00",x"00",x"15",x"59"),
   761 => (x"03",x"13",x"27",x"1e"),
   762 => (x"c8",x"0f",x"00",x"00"),
   763 => (x"17",x"54",x"27",x"86"),
   764 => (x"49",x"bf",x"00",x"00"),
   765 => (x"1e",x"71",x"81",x"d0"),
   766 => (x"00",x"15",x"72",x"27"),
   767 => (x"13",x"27",x"1e",x"00"),
   768 => (x"0f",x"00",x"00",x"03"),
   769 => (x"8b",x"27",x"86",x"c8"),
   770 => (x"1e",x"00",x"00",x"15"),
   771 => (x"00",x"03",x"13",x"27"),
   772 => (x"86",x"c4",x"0f",x"00"),
   773 => (x"c0",x"27",x"1e",x"6e"),
   774 => (x"1e",x"00",x"00",x"15"),
   775 => (x"00",x"03",x"13",x"27"),
   776 => (x"86",x"c8",x"0f",x"00"),
   777 => (x"d9",x"27",x"1e",x"c5"),
   778 => (x"1e",x"00",x"00",x"15"),
   779 => (x"00",x"03",x"13",x"27"),
   780 => (x"86",x"c8",x"0f",x"00"),
   781 => (x"f2",x"27",x"1e",x"73"),
   782 => (x"1e",x"00",x"00",x"15"),
   783 => (x"00",x"03",x"13",x"27"),
   784 => (x"86",x"c8",x"0f",x"00"),
   785 => (x"0b",x"27",x"1e",x"cd"),
   786 => (x"1e",x"00",x"00",x"16"),
   787 => (x"00",x"03",x"13",x"27"),
   788 => (x"86",x"c8",x"0f",x"00"),
   789 => (x"27",x"1e",x"66",x"cc"),
   790 => (x"00",x"00",x"16",x"24"),
   791 => (x"03",x"13",x"27",x"1e"),
   792 => (x"c8",x"0f",x"00",x"00"),
   793 => (x"27",x"1e",x"c7",x"86"),
   794 => (x"00",x"00",x"16",x"3d"),
   795 => (x"03",x"13",x"27",x"1e"),
   796 => (x"c8",x"0f",x"00",x"00"),
   797 => (x"1e",x"66",x"c8",x"86"),
   798 => (x"00",x"16",x"56",x"27"),
   799 => (x"13",x"27",x"1e",x"00"),
   800 => (x"0f",x"00",x"00",x"03"),
   801 => (x"1e",x"c1",x"86",x"c8"),
   802 => (x"00",x"16",x"6f",x"27"),
   803 => (x"13",x"27",x"1e",x"00"),
   804 => (x"0f",x"00",x"00",x"03"),
   805 => (x"b8",x"27",x"86",x"c8"),
   806 => (x"1e",x"00",x"00",x"3f"),
   807 => (x"00",x"16",x"88",x"27"),
   808 => (x"13",x"27",x"1e",x"00"),
   809 => (x"0f",x"00",x"00",x"03"),
   810 => (x"a1",x"27",x"86",x"c8"),
   811 => (x"1e",x"00",x"00",x"16"),
   812 => (x"00",x"03",x"13",x"27"),
   813 => (x"86",x"c4",x"0f",x"00"),
   814 => (x"00",x"3f",x"d8",x"27"),
   815 => (x"d6",x"27",x"1e",x"00"),
   816 => (x"1e",x"00",x"00",x"16"),
   817 => (x"00",x"03",x"13",x"27"),
   818 => (x"86",x"c8",x"0f",x"00"),
   819 => (x"00",x"16",x"ef",x"27"),
   820 => (x"13",x"27",x"1e",x"00"),
   821 => (x"0f",x"00",x"00",x"03"),
   822 => (x"24",x"27",x"86",x"c4"),
   823 => (x"1e",x"00",x"00",x"17"),
   824 => (x"00",x"03",x"13",x"27"),
   825 => (x"86",x"c4",x"0f",x"00"),
   826 => (x"00",x"3f",x"44",x"27"),
   827 => (x"27",x"49",x"bf",x"00"),
   828 => (x"00",x"00",x"3f",x"40"),
   829 => (x"4c",x"27",x"89",x"bf"),
   830 => (x"59",x"00",x"00",x"3f"),
   831 => (x"26",x"27",x"1e",x"71"),
   832 => (x"1e",x"00",x"00",x"17"),
   833 => (x"00",x"03",x"13",x"27"),
   834 => (x"86",x"c8",x"0f",x"00"),
   835 => (x"00",x"3f",x"48",x"27"),
   836 => (x"c1",x"48",x"bf",x"00"),
   837 => (x"03",x"a8",x"b7",x"f8"),
   838 => (x"27",x"87",x"ea",x"c0"),
   839 => (x"00",x"00",x"10",x"36"),
   840 => (x"03",x"13",x"27",x"1e"),
   841 => (x"c4",x"0f",x"00",x"00"),
   842 => (x"10",x"6c",x"27",x"86"),
   843 => (x"27",x"1e",x"00",x"00"),
   844 => (x"00",x"00",x"03",x"13"),
   845 => (x"27",x"86",x"c4",x"0f"),
   846 => (x"00",x"00",x"10",x"8c"),
   847 => (x"03",x"13",x"27",x"1e"),
   848 => (x"c4",x"0f",x"00",x"00"),
   849 => (x"3f",x"48",x"27",x"86"),
   850 => (x"49",x"bf",x"00",x"00"),
   851 => (x"e8",x"cf",x"4a",x"71"),
   852 => (x"72",x"1e",x"71",x"92"),
   853 => (x"27",x"49",x"72",x"1e"),
   854 => (x"00",x"00",x"17",x"3c"),
   855 => (x"26",x"27",x"4a",x"bf"),
   856 => (x"0f",x"00",x"00",x"06"),
   857 => (x"49",x"26",x"4a",x"26"),
   858 => (x"00",x"3f",x"50",x"27"),
   859 => (x"3c",x"27",x"58",x"00"),
   860 => (x"bf",x"00",x"00",x"17"),
   861 => (x"cf",x"4b",x"72",x"4a"),
   862 => (x"1e",x"71",x"93",x"e8"),
   863 => (x"09",x"73",x"1e",x"72"),
   864 => (x"06",x"26",x"27",x"4a"),
   865 => (x"26",x"0f",x"00",x"00"),
   866 => (x"27",x"49",x"26",x"4a"),
   867 => (x"00",x"00",x"3f",x"54"),
   868 => (x"92",x"f9",x"c8",x"58"),
   869 => (x"1e",x"72",x"1e",x"71"),
   870 => (x"27",x"4a",x"09",x"72"),
   871 => (x"00",x"00",x"06",x"26"),
   872 => (x"26",x"4a",x"26",x"0f"),
   873 => (x"3f",x"58",x"27",x"49"),
   874 => (x"27",x"58",x"00",x"00"),
   875 => (x"00",x"00",x"10",x"8e"),
   876 => (x"03",x"13",x"27",x"1e"),
   877 => (x"c4",x"0f",x"00",x"00"),
   878 => (x"3f",x"4c",x"27",x"86"),
   879 => (x"1e",x"bf",x"00",x"00"),
   880 => (x"00",x"10",x"bb",x"27"),
   881 => (x"13",x"27",x"1e",x"00"),
   882 => (x"0f",x"00",x"00",x"03"),
   883 => (x"c0",x"27",x"86",x"c8"),
   884 => (x"1e",x"00",x"00",x"10"),
   885 => (x"00",x"03",x"13",x"27"),
   886 => (x"86",x"c4",x"0f",x"00"),
   887 => (x"00",x"3f",x"50",x"27"),
   888 => (x"27",x"1e",x"bf",x"00"),
   889 => (x"00",x"00",x"10",x"ed"),
   890 => (x"03",x"13",x"27",x"1e"),
   891 => (x"c8",x"0f",x"00",x"00"),
   892 => (x"3f",x"54",x"27",x"86"),
   893 => (x"1e",x"bf",x"00",x"00"),
   894 => (x"00",x"10",x"f2",x"27"),
   895 => (x"13",x"27",x"1e",x"00"),
   896 => (x"0f",x"00",x"00",x"03"),
   897 => (x"10",x"27",x"86",x"c8"),
   898 => (x"1e",x"00",x"00",x"11"),
   899 => (x"00",x"03",x"13",x"27"),
   900 => (x"86",x"c4",x"0f",x"00"),
   901 => (x"8e",x"f0",x"48",x"c0"),
   902 => (x"4c",x"26",x"4d",x"26"),
   903 => (x"4f",x"26",x"4b",x"26"),
   904 => (x"5c",x"5b",x"5e",x"0e"),
   905 => (x"66",x"d0",x"0e",x"5d"),
   906 => (x"73",x"4b",x"6d",x"4d"),
   907 => (x"27",x"1e",x"73",x"4c"),
   908 => (x"00",x"00",x"17",x"50"),
   909 => (x"f0",x"c0",x"48",x"bf"),
   910 => (x"43",x"20",x"4a",x"a3"),
   911 => (x"f9",x"05",x"aa",x"73"),
   912 => (x"75",x"4a",x"26",x"87"),
   913 => (x"c5",x"82",x"cc",x"4a"),
   914 => (x"cc",x"49",x"73",x"7a"),
   915 => (x"6d",x"79",x"6a",x"81"),
   916 => (x"27",x"1e",x"73",x"7b"),
   917 => (x"00",x"00",x"0f",x"02"),
   918 => (x"73",x"86",x"c4",x"0f"),
   919 => (x"69",x"81",x"c4",x"49"),
   920 => (x"87",x"f3",x"c0",x"05"),
   921 => (x"81",x"c8",x"49",x"74"),
   922 => (x"83",x"cc",x"4b",x"74"),
   923 => (x"1e",x"71",x"7b",x"c6"),
   924 => (x"81",x"c8",x"49",x"75"),
   925 => (x"d2",x"27",x"1e",x"69"),
   926 => (x"0f",x"00",x"00",x"03"),
   927 => (x"50",x"27",x"86",x"c8"),
   928 => (x"bf",x"00",x"00",x"17"),
   929 => (x"1e",x"73",x"7c",x"bf"),
   930 => (x"1e",x"6b",x"1e",x"ca"),
   931 => (x"00",x"04",x"3e",x"27"),
   932 => (x"86",x"cc",x"0f",x"00"),
   933 => (x"6d",x"87",x"d0",x"c0"),
   934 => (x"48",x"4a",x"75",x"49"),
   935 => (x"4b",x"a2",x"f0",x"c0"),
   936 => (x"ab",x"72",x"42",x"20"),
   937 => (x"26",x"87",x"f9",x"05"),
   938 => (x"26",x"4c",x"26",x"4d"),
   939 => (x"0e",x"4f",x"26",x"4b"),
   940 => (x"5d",x"5c",x"5b",x"5e"),
   941 => (x"27",x"86",x"fc",x"0e"),
   942 => (x"00",x"00",x"17",x"60"),
   943 => (x"6e",x"4d",x"bf",x"97"),
   944 => (x"4b",x"66",x"d4",x"4c"),
   945 => (x"82",x"ca",x"4a",x"6b"),
   946 => (x"c0",x"c1",x"49",x"75"),
   947 => (x"91",x"c0",x"c0",x"c0"),
   948 => (x"91",x"b7",x"c0",x"c4"),
   949 => (x"a9",x"c1",x"c1",x"49"),
   950 => (x"87",x"cf",x"c0",x"05"),
   951 => (x"48",x"72",x"8a",x"c1"),
   952 => (x"00",x"17",x"58",x"27"),
   953 => (x"70",x"88",x"bf",x"00"),
   954 => (x"74",x"4c",x"c0",x"7b"),
   955 => (x"d7",x"ff",x"05",x"9c"),
   956 => (x"17",x"64",x"27",x"87"),
   957 => (x"5d",x"97",x"00",x"00"),
   958 => (x"4d",x"26",x"8e",x"fc"),
   959 => (x"4b",x"26",x"4c",x"26"),
   960 => (x"27",x"1e",x"4f",x"26"),
   961 => (x"00",x"00",x"17",x"50"),
   962 => (x"cb",x"c0",x"02",x"bf"),
   963 => (x"48",x"66",x"c4",x"87"),
   964 => (x"00",x"17",x"50",x"27"),
   965 => (x"78",x"bf",x"bf",x"00"),
   966 => (x"00",x"17",x"50",x"27"),
   967 => (x"cc",x"49",x"bf",x"00"),
   968 => (x"27",x"1e",x"71",x"81"),
   969 => (x"00",x"00",x"17",x"58"),
   970 => (x"1e",x"ca",x"1e",x"bf"),
   971 => (x"00",x"04",x"3e",x"27"),
   972 => (x"86",x"cc",x"0f",x"00"),
   973 => (x"27",x"1e",x"4f",x"26"),
   974 => (x"00",x"00",x"17",x"60"),
   975 => (x"c1",x"49",x"bf",x"97"),
   976 => (x"c0",x"c0",x"c0",x"c0"),
   977 => (x"b7",x"c0",x"c4",x"91"),
   978 => (x"c1",x"c1",x"49",x"91"),
   979 => (x"c5",x"c0",x"02",x"a9"),
   980 => (x"c0",x"49",x"c0",x"87"),
   981 => (x"49",x"c1",x"87",x"c2"),
   982 => (x"00",x"17",x"5c",x"27"),
   983 => (x"71",x"48",x"bf",x"00"),
   984 => (x"17",x"60",x"27",x"b0"),
   985 => (x"27",x"58",x"00",x"00"),
   986 => (x"00",x"00",x"17",x"61"),
   987 => (x"50",x"c2",x"c1",x"48"),
   988 => (x"27",x"1e",x"4f",x"26"),
   989 => (x"00",x"00",x"17",x"60"),
   990 => (x"50",x"c1",x"c1",x"48"),
   991 => (x"00",x"17",x"5c",x"27"),
   992 => (x"78",x"c0",x"48",x"00"),
   993 => (x"00",x"00",x"4f",x"26"),
   994 => (x"33",x"32",x"31",x"30"),
   995 => (x"37",x"36",x"35",x"34"),
   996 => (x"42",x"41",x"39",x"38"),
   997 => (x"46",x"45",x"44",x"43"),
   998 => (x"6f",x"72",x"50",x"00"),
   999 => (x"6d",x"61",x"72",x"67"),
  1000 => (x"6d",x"6f",x"63",x"20"),
  1001 => (x"65",x"6c",x"69",x"70"),
  1002 => (x"69",x"77",x"20",x"64"),
  1003 => (x"27",x"20",x"68",x"74"),
  1004 => (x"69",x"67",x"65",x"72"),
  1005 => (x"72",x"65",x"74",x"73"),
  1006 => (x"74",x"61",x"20",x"27"),
  1007 => (x"62",x"69",x"72",x"74"),
  1008 => (x"0a",x"65",x"74",x"75"),
  1009 => (x"50",x"00",x"0a",x"00"),
  1010 => (x"72",x"67",x"6f",x"72"),
  1011 => (x"63",x"20",x"6d",x"61"),
  1012 => (x"69",x"70",x"6d",x"6f"),
  1013 => (x"20",x"64",x"65",x"6c"),
  1014 => (x"68",x"74",x"69",x"77"),
  1015 => (x"20",x"74",x"75",x"6f"),
  1016 => (x"67",x"65",x"72",x"27"),
  1017 => (x"65",x"74",x"73",x"69"),
  1018 => (x"61",x"20",x"27",x"72"),
  1019 => (x"69",x"72",x"74",x"74"),
  1020 => (x"65",x"74",x"75",x"62"),
  1021 => (x"00",x"0a",x"00",x"0a"),
  1022 => (x"59",x"52",x"48",x"44"),
  1023 => (x"4e",x"4f",x"54",x"53"),
  1024 => (x"52",x"50",x"20",x"45"),
  1025 => (x"41",x"52",x"47",x"4f"),
  1026 => (x"33",x"20",x"2c",x"4d"),
  1027 => (x"20",x"44",x"52",x"27"),
  1028 => (x"49",x"52",x"54",x"53"),
  1029 => (x"44",x"00",x"47",x"4e"),
  1030 => (x"53",x"59",x"52",x"48"),
  1031 => (x"45",x"4e",x"4f",x"54"),
  1032 => (x"4f",x"52",x"50",x"20"),
  1033 => (x"4d",x"41",x"52",x"47"),
  1034 => (x"27",x"32",x"20",x"2c"),
  1035 => (x"53",x"20",x"44",x"4e"),
  1036 => (x"4e",x"49",x"52",x"54"),
  1037 => (x"65",x"4d",x"00",x"47"),
  1038 => (x"72",x"75",x"73",x"61"),
  1039 => (x"74",x"20",x"64",x"65"),
  1040 => (x"20",x"65",x"6d",x"69"),
  1041 => (x"20",x"6f",x"6f",x"74"),
  1042 => (x"6c",x"61",x"6d",x"73"),
  1043 => (x"6f",x"74",x"20",x"6c"),
  1044 => (x"74",x"62",x"6f",x"20"),
  1045 => (x"20",x"6e",x"69",x"61"),
  1046 => (x"6e",x"61",x"65",x"6d"),
  1047 => (x"66",x"67",x"6e",x"69"),
  1048 => (x"72",x"20",x"6c",x"75"),
  1049 => (x"6c",x"75",x"73",x"65"),
  1050 => (x"00",x"0a",x"73",x"74"),
  1051 => (x"61",x"65",x"6c",x"50"),
  1052 => (x"69",x"20",x"65",x"73"),
  1053 => (x"65",x"72",x"63",x"6e"),
  1054 => (x"20",x"65",x"73",x"61"),
  1055 => (x"62",x"6d",x"75",x"6e"),
  1056 => (x"6f",x"20",x"72",x"65"),
  1057 => (x"75",x"72",x"20",x"66"),
  1058 => (x"00",x"0a",x"73",x"6e"),
  1059 => (x"69",x"4d",x"00",x"0a"),
  1060 => (x"73",x"6f",x"72",x"63"),
  1061 => (x"6e",x"6f",x"63",x"65"),
  1062 => (x"66",x"20",x"73",x"64"),
  1063 => (x"6f",x"20",x"72",x"6f"),
  1064 => (x"72",x"20",x"65",x"6e"),
  1065 => (x"74",x"20",x"6e",x"75"),
  1066 => (x"75",x"6f",x"72",x"68"),
  1067 => (x"44",x"20",x"68",x"67"),
  1068 => (x"73",x"79",x"72",x"68"),
  1069 => (x"65",x"6e",x"6f",x"74"),
  1070 => (x"25",x"00",x"20",x"3a"),
  1071 => (x"00",x"0a",x"20",x"64"),
  1072 => (x"79",x"72",x"68",x"44"),
  1073 => (x"6e",x"6f",x"74",x"73"),
  1074 => (x"70",x"20",x"73",x"65"),
  1075 => (x"53",x"20",x"72",x"65"),
  1076 => (x"6e",x"6f",x"63",x"65"),
  1077 => (x"20",x"20",x"3a",x"64"),
  1078 => (x"20",x"20",x"20",x"20"),
  1079 => (x"20",x"20",x"20",x"20"),
  1080 => (x"20",x"20",x"20",x"20"),
  1081 => (x"20",x"20",x"20",x"20"),
  1082 => (x"20",x"20",x"20",x"20"),
  1083 => (x"20",x"64",x"25",x"00"),
  1084 => (x"41",x"56",x"00",x"0a"),
  1085 => (x"49",x"4d",x"20",x"58"),
  1086 => (x"72",x"20",x"53",x"50"),
  1087 => (x"6e",x"69",x"74",x"61"),
  1088 => (x"20",x"2a",x"20",x"67"),
  1089 => (x"30",x"30",x"30",x"31"),
  1090 => (x"25",x"20",x"3d",x"20"),
  1091 => (x"00",x"0a",x"20",x"64"),
  1092 => (x"48",x"44",x"00",x"0a"),
  1093 => (x"54",x"53",x"59",x"52"),
  1094 => (x"20",x"45",x"4e",x"4f"),
  1095 => (x"47",x"4f",x"52",x"50"),
  1096 => (x"2c",x"4d",x"41",x"52"),
  1097 => (x"4d",x"4f",x"53",x"20"),
  1098 => (x"54",x"53",x"20",x"45"),
  1099 => (x"47",x"4e",x"49",x"52"),
  1100 => (x"52",x"48",x"44",x"00"),
  1101 => (x"4f",x"54",x"53",x"59"),
  1102 => (x"50",x"20",x"45",x"4e"),
  1103 => (x"52",x"47",x"4f",x"52"),
  1104 => (x"20",x"2c",x"4d",x"41"),
  1105 => (x"54",x"53",x"27",x"31"),
  1106 => (x"52",x"54",x"53",x"20"),
  1107 => (x"00",x"47",x"4e",x"49"),
  1108 => (x"68",x"44",x"00",x"0a"),
  1109 => (x"74",x"73",x"79",x"72"),
  1110 => (x"20",x"65",x"6e",x"6f"),
  1111 => (x"63",x"6e",x"65",x"42"),
  1112 => (x"72",x"61",x"6d",x"68"),
  1113 => (x"56",x"20",x"2c",x"6b"),
  1114 => (x"69",x"73",x"72",x"65"),
  1115 => (x"32",x"20",x"6e",x"6f"),
  1116 => (x"28",x"20",x"31",x"2e"),
  1117 => (x"67",x"6e",x"61",x"4c"),
  1118 => (x"65",x"67",x"61",x"75"),
  1119 => (x"29",x"43",x"20",x"3a"),
  1120 => (x"00",x"0a",x"00",x"0a"),
  1121 => (x"63",x"65",x"78",x"45"),
  1122 => (x"6f",x"69",x"74",x"75"),
  1123 => (x"74",x"73",x"20",x"6e"),
  1124 => (x"73",x"74",x"72",x"61"),
  1125 => (x"64",x"25",x"20",x"2c"),
  1126 => (x"6e",x"75",x"72",x"20"),
  1127 => (x"68",x"74",x"20",x"73"),
  1128 => (x"67",x"75",x"6f",x"72"),
  1129 => (x"68",x"44",x"20",x"68"),
  1130 => (x"74",x"73",x"79",x"72"),
  1131 => (x"0a",x"65",x"6e",x"6f"),
  1132 => (x"65",x"78",x"45",x"00"),
  1133 => (x"69",x"74",x"75",x"63"),
  1134 => (x"65",x"20",x"6e",x"6f"),
  1135 => (x"0a",x"73",x"64",x"6e"),
  1136 => (x"46",x"00",x"0a",x"00"),
  1137 => (x"6c",x"61",x"6e",x"69"),
  1138 => (x"6c",x"61",x"76",x"20"),
  1139 => (x"20",x"73",x"65",x"75"),
  1140 => (x"74",x"20",x"66",x"6f"),
  1141 => (x"76",x"20",x"65",x"68"),
  1142 => (x"61",x"69",x"72",x"61"),
  1143 => (x"73",x"65",x"6c",x"62"),
  1144 => (x"65",x"73",x"75",x"20"),
  1145 => (x"6e",x"69",x"20",x"64"),
  1146 => (x"65",x"68",x"74",x"20"),
  1147 => (x"6e",x"65",x"62",x"20"),
  1148 => (x"61",x"6d",x"68",x"63"),
  1149 => (x"0a",x"3a",x"6b",x"72"),
  1150 => (x"49",x"00",x"0a",x"00"),
  1151 => (x"47",x"5f",x"74",x"6e"),
  1152 => (x"3a",x"62",x"6f",x"6c"),
  1153 => (x"20",x"20",x"20",x"20"),
  1154 => (x"20",x"20",x"20",x"20"),
  1155 => (x"20",x"20",x"20",x"20"),
  1156 => (x"00",x"0a",x"64",x"25"),
  1157 => (x"20",x"20",x"20",x"20"),
  1158 => (x"20",x"20",x"20",x"20"),
  1159 => (x"75",x"6f",x"68",x"73"),
  1160 => (x"62",x"20",x"64",x"6c"),
  1161 => (x"20",x"20",x"3a",x"65"),
  1162 => (x"0a",x"64",x"25",x"20"),
  1163 => (x"6f",x"6f",x"42",x"00"),
  1164 => (x"6c",x"47",x"5f",x"6c"),
  1165 => (x"20",x"3a",x"62",x"6f"),
  1166 => (x"20",x"20",x"20",x"20"),
  1167 => (x"20",x"20",x"20",x"20"),
  1168 => (x"64",x"25",x"20",x"20"),
  1169 => (x"20",x"20",x"00",x"0a"),
  1170 => (x"20",x"20",x"20",x"20"),
  1171 => (x"68",x"73",x"20",x"20"),
  1172 => (x"64",x"6c",x"75",x"6f"),
  1173 => (x"3a",x"65",x"62",x"20"),
  1174 => (x"25",x"20",x"20",x"20"),
  1175 => (x"43",x"00",x"0a",x"64"),
  1176 => (x"5f",x"31",x"5f",x"68"),
  1177 => (x"62",x"6f",x"6c",x"47"),
  1178 => (x"20",x"20",x"20",x"3a"),
  1179 => (x"20",x"20",x"20",x"20"),
  1180 => (x"20",x"20",x"20",x"20"),
  1181 => (x"00",x"0a",x"63",x"25"),
  1182 => (x"20",x"20",x"20",x"20"),
  1183 => (x"20",x"20",x"20",x"20"),
  1184 => (x"75",x"6f",x"68",x"73"),
  1185 => (x"62",x"20",x"64",x"6c"),
  1186 => (x"20",x"20",x"3a",x"65"),
  1187 => (x"0a",x"63",x"25",x"20"),
  1188 => (x"5f",x"68",x"43",x"00"),
  1189 => (x"6c",x"47",x"5f",x"32"),
  1190 => (x"20",x"3a",x"62",x"6f"),
  1191 => (x"20",x"20",x"20",x"20"),
  1192 => (x"20",x"20",x"20",x"20"),
  1193 => (x"63",x"25",x"20",x"20"),
  1194 => (x"20",x"20",x"00",x"0a"),
  1195 => (x"20",x"20",x"20",x"20"),
  1196 => (x"68",x"73",x"20",x"20"),
  1197 => (x"64",x"6c",x"75",x"6f"),
  1198 => (x"3a",x"65",x"62",x"20"),
  1199 => (x"25",x"20",x"20",x"20"),
  1200 => (x"41",x"00",x"0a",x"63"),
  1201 => (x"31",x"5f",x"72",x"72"),
  1202 => (x"6f",x"6c",x"47",x"5f"),
  1203 => (x"5d",x"38",x"5b",x"62"),
  1204 => (x"20",x"20",x"20",x"3a"),
  1205 => (x"20",x"20",x"20",x"20"),
  1206 => (x"00",x"0a",x"64",x"25"),
  1207 => (x"20",x"20",x"20",x"20"),
  1208 => (x"20",x"20",x"20",x"20"),
  1209 => (x"75",x"6f",x"68",x"73"),
  1210 => (x"62",x"20",x"64",x"6c"),
  1211 => (x"20",x"20",x"3a",x"65"),
  1212 => (x"0a",x"64",x"25",x"20"),
  1213 => (x"72",x"72",x"41",x"00"),
  1214 => (x"47",x"5f",x"32",x"5f"),
  1215 => (x"5b",x"62",x"6f",x"6c"),
  1216 => (x"37",x"5b",x"5d",x"38"),
  1217 => (x"20",x"20",x"3a",x"5d"),
  1218 => (x"64",x"25",x"20",x"20"),
  1219 => (x"20",x"20",x"00",x"0a"),
  1220 => (x"20",x"20",x"20",x"20"),
  1221 => (x"68",x"73",x"20",x"20"),
  1222 => (x"64",x"6c",x"75",x"6f"),
  1223 => (x"3a",x"65",x"62",x"20"),
  1224 => (x"4e",x"20",x"20",x"20"),
  1225 => (x"65",x"62",x"6d",x"75"),
  1226 => (x"66",x"4f",x"5f",x"72"),
  1227 => (x"6e",x"75",x"52",x"5f"),
  1228 => (x"20",x"2b",x"20",x"73"),
  1229 => (x"00",x"0a",x"30",x"31"),
  1230 => (x"5f",x"72",x"74",x"50"),
  1231 => (x"62",x"6f",x"6c",x"47"),
  1232 => (x"00",x"0a",x"3e",x"2d"),
  1233 => (x"74",x"50",x"20",x"20"),
  1234 => (x"6f",x"43",x"5f",x"72"),
  1235 => (x"20",x"3a",x"70",x"6d"),
  1236 => (x"20",x"20",x"20",x"20"),
  1237 => (x"20",x"20",x"20",x"20"),
  1238 => (x"0a",x"64",x"25",x"20"),
  1239 => (x"20",x"20",x"20",x"00"),
  1240 => (x"20",x"20",x"20",x"20"),
  1241 => (x"6f",x"68",x"73",x"20"),
  1242 => (x"20",x"64",x"6c",x"75"),
  1243 => (x"20",x"3a",x"65",x"62"),
  1244 => (x"69",x"28",x"20",x"20"),
  1245 => (x"65",x"6c",x"70",x"6d"),
  1246 => (x"74",x"6e",x"65",x"6d"),
  1247 => (x"6f",x"69",x"74",x"61"),
  1248 => (x"65",x"64",x"2d",x"6e"),
  1249 => (x"64",x"6e",x"65",x"70"),
  1250 => (x"29",x"74",x"6e",x"65"),
  1251 => (x"20",x"20",x"00",x"0a"),
  1252 => (x"63",x"73",x"69",x"44"),
  1253 => (x"20",x"20",x"3a",x"72"),
  1254 => (x"20",x"20",x"20",x"20"),
  1255 => (x"20",x"20",x"20",x"20"),
  1256 => (x"25",x"20",x"20",x"20"),
  1257 => (x"20",x"00",x"0a",x"64"),
  1258 => (x"20",x"20",x"20",x"20"),
  1259 => (x"73",x"20",x"20",x"20"),
  1260 => (x"6c",x"75",x"6f",x"68"),
  1261 => (x"65",x"62",x"20",x"64"),
  1262 => (x"20",x"20",x"20",x"3a"),
  1263 => (x"00",x"0a",x"64",x"25"),
  1264 => (x"6e",x"45",x"20",x"20"),
  1265 => (x"43",x"5f",x"6d",x"75"),
  1266 => (x"3a",x"70",x"6d",x"6f"),
  1267 => (x"20",x"20",x"20",x"20"),
  1268 => (x"20",x"20",x"20",x"20"),
  1269 => (x"0a",x"64",x"25",x"20"),
  1270 => (x"20",x"20",x"20",x"00"),
  1271 => (x"20",x"20",x"20",x"20"),
  1272 => (x"6f",x"68",x"73",x"20"),
  1273 => (x"20",x"64",x"6c",x"75"),
  1274 => (x"20",x"3a",x"65",x"62"),
  1275 => (x"64",x"25",x"20",x"20"),
  1276 => (x"20",x"20",x"00",x"0a"),
  1277 => (x"5f",x"74",x"6e",x"49"),
  1278 => (x"70",x"6d",x"6f",x"43"),
  1279 => (x"20",x"20",x"20",x"3a"),
  1280 => (x"20",x"20",x"20",x"20"),
  1281 => (x"25",x"20",x"20",x"20"),
  1282 => (x"20",x"00",x"0a",x"64"),
  1283 => (x"20",x"20",x"20",x"20"),
  1284 => (x"73",x"20",x"20",x"20"),
  1285 => (x"6c",x"75",x"6f",x"68"),
  1286 => (x"65",x"62",x"20",x"64"),
  1287 => (x"20",x"20",x"20",x"3a"),
  1288 => (x"00",x"0a",x"64",x"25"),
  1289 => (x"74",x"53",x"20",x"20"),
  1290 => (x"6f",x"43",x"5f",x"72"),
  1291 => (x"20",x"3a",x"70",x"6d"),
  1292 => (x"20",x"20",x"20",x"20"),
  1293 => (x"20",x"20",x"20",x"20"),
  1294 => (x"0a",x"73",x"25",x"20"),
  1295 => (x"20",x"20",x"20",x"00"),
  1296 => (x"20",x"20",x"20",x"20"),
  1297 => (x"6f",x"68",x"73",x"20"),
  1298 => (x"20",x"64",x"6c",x"75"),
  1299 => (x"20",x"3a",x"65",x"62"),
  1300 => (x"48",x"44",x"20",x"20"),
  1301 => (x"54",x"53",x"59",x"52"),
  1302 => (x"20",x"45",x"4e",x"4f"),
  1303 => (x"47",x"4f",x"52",x"50"),
  1304 => (x"2c",x"4d",x"41",x"52"),
  1305 => (x"4d",x"4f",x"53",x"20"),
  1306 => (x"54",x"53",x"20",x"45"),
  1307 => (x"47",x"4e",x"49",x"52"),
  1308 => (x"65",x"4e",x"00",x"0a"),
  1309 => (x"50",x"5f",x"74",x"78"),
  1310 => (x"47",x"5f",x"72",x"74"),
  1311 => (x"2d",x"62",x"6f",x"6c"),
  1312 => (x"20",x"00",x"0a",x"3e"),
  1313 => (x"72",x"74",x"50",x"20"),
  1314 => (x"6d",x"6f",x"43",x"5f"),
  1315 => (x"20",x"20",x"3a",x"70"),
  1316 => (x"20",x"20",x"20",x"20"),
  1317 => (x"20",x"20",x"20",x"20"),
  1318 => (x"00",x"0a",x"64",x"25"),
  1319 => (x"20",x"20",x"20",x"20"),
  1320 => (x"20",x"20",x"20",x"20"),
  1321 => (x"75",x"6f",x"68",x"73"),
  1322 => (x"62",x"20",x"64",x"6c"),
  1323 => (x"20",x"20",x"3a",x"65"),
  1324 => (x"6d",x"69",x"28",x"20"),
  1325 => (x"6d",x"65",x"6c",x"70"),
  1326 => (x"61",x"74",x"6e",x"65"),
  1327 => (x"6e",x"6f",x"69",x"74"),
  1328 => (x"70",x"65",x"64",x"2d"),
  1329 => (x"65",x"64",x"6e",x"65"),
  1330 => (x"2c",x"29",x"74",x"6e"),
  1331 => (x"6d",x"61",x"73",x"20"),
  1332 => (x"73",x"61",x"20",x"65"),
  1333 => (x"6f",x"62",x"61",x"20"),
  1334 => (x"00",x"0a",x"65",x"76"),
  1335 => (x"69",x"44",x"20",x"20"),
  1336 => (x"3a",x"72",x"63",x"73"),
  1337 => (x"20",x"20",x"20",x"20"),
  1338 => (x"20",x"20",x"20",x"20"),
  1339 => (x"20",x"20",x"20",x"20"),
  1340 => (x"0a",x"64",x"25",x"20"),
  1341 => (x"20",x"20",x"20",x"00"),
  1342 => (x"20",x"20",x"20",x"20"),
  1343 => (x"6f",x"68",x"73",x"20"),
  1344 => (x"20",x"64",x"6c",x"75"),
  1345 => (x"20",x"3a",x"65",x"62"),
  1346 => (x"64",x"25",x"20",x"20"),
  1347 => (x"20",x"20",x"00",x"0a"),
  1348 => (x"6d",x"75",x"6e",x"45"),
  1349 => (x"6d",x"6f",x"43",x"5f"),
  1350 => (x"20",x"20",x"3a",x"70"),
  1351 => (x"20",x"20",x"20",x"20"),
  1352 => (x"25",x"20",x"20",x"20"),
  1353 => (x"20",x"00",x"0a",x"64"),
  1354 => (x"20",x"20",x"20",x"20"),
  1355 => (x"73",x"20",x"20",x"20"),
  1356 => (x"6c",x"75",x"6f",x"68"),
  1357 => (x"65",x"62",x"20",x"64"),
  1358 => (x"20",x"20",x"20",x"3a"),
  1359 => (x"00",x"0a",x"64",x"25"),
  1360 => (x"6e",x"49",x"20",x"20"),
  1361 => (x"6f",x"43",x"5f",x"74"),
  1362 => (x"20",x"3a",x"70",x"6d"),
  1363 => (x"20",x"20",x"20",x"20"),
  1364 => (x"20",x"20",x"20",x"20"),
  1365 => (x"0a",x"64",x"25",x"20"),
  1366 => (x"20",x"20",x"20",x"00"),
  1367 => (x"20",x"20",x"20",x"20"),
  1368 => (x"6f",x"68",x"73",x"20"),
  1369 => (x"20",x"64",x"6c",x"75"),
  1370 => (x"20",x"3a",x"65",x"62"),
  1371 => (x"64",x"25",x"20",x"20"),
  1372 => (x"20",x"20",x"00",x"0a"),
  1373 => (x"5f",x"72",x"74",x"53"),
  1374 => (x"70",x"6d",x"6f",x"43"),
  1375 => (x"20",x"20",x"20",x"3a"),
  1376 => (x"20",x"20",x"20",x"20"),
  1377 => (x"25",x"20",x"20",x"20"),
  1378 => (x"20",x"00",x"0a",x"73"),
  1379 => (x"20",x"20",x"20",x"20"),
  1380 => (x"73",x"20",x"20",x"20"),
  1381 => (x"6c",x"75",x"6f",x"68"),
  1382 => (x"65",x"62",x"20",x"64"),
  1383 => (x"20",x"20",x"20",x"3a"),
  1384 => (x"59",x"52",x"48",x"44"),
  1385 => (x"4e",x"4f",x"54",x"53"),
  1386 => (x"52",x"50",x"20",x"45"),
  1387 => (x"41",x"52",x"47",x"4f"),
  1388 => (x"53",x"20",x"2c",x"4d"),
  1389 => (x"20",x"45",x"4d",x"4f"),
  1390 => (x"49",x"52",x"54",x"53"),
  1391 => (x"00",x"0a",x"47",x"4e"),
  1392 => (x"5f",x"74",x"6e",x"49"),
  1393 => (x"6f",x"4c",x"5f",x"31"),
  1394 => (x"20",x"20",x"3a",x"63"),
  1395 => (x"20",x"20",x"20",x"20"),
  1396 => (x"20",x"20",x"20",x"20"),
  1397 => (x"0a",x"64",x"25",x"20"),
  1398 => (x"20",x"20",x"20",x"00"),
  1399 => (x"20",x"20",x"20",x"20"),
  1400 => (x"6f",x"68",x"73",x"20"),
  1401 => (x"20",x"64",x"6c",x"75"),
  1402 => (x"20",x"3a",x"65",x"62"),
  1403 => (x"64",x"25",x"20",x"20"),
  1404 => (x"6e",x"49",x"00",x"0a"),
  1405 => (x"5f",x"32",x"5f",x"74"),
  1406 => (x"3a",x"63",x"6f",x"4c"),
  1407 => (x"20",x"20",x"20",x"20"),
  1408 => (x"20",x"20",x"20",x"20"),
  1409 => (x"25",x"20",x"20",x"20"),
  1410 => (x"20",x"00",x"0a",x"64"),
  1411 => (x"20",x"20",x"20",x"20"),
  1412 => (x"73",x"20",x"20",x"20"),
  1413 => (x"6c",x"75",x"6f",x"68"),
  1414 => (x"65",x"62",x"20",x"64"),
  1415 => (x"20",x"20",x"20",x"3a"),
  1416 => (x"00",x"0a",x"64",x"25"),
  1417 => (x"5f",x"74",x"6e",x"49"),
  1418 => (x"6f",x"4c",x"5f",x"33"),
  1419 => (x"20",x"20",x"3a",x"63"),
  1420 => (x"20",x"20",x"20",x"20"),
  1421 => (x"20",x"20",x"20",x"20"),
  1422 => (x"0a",x"64",x"25",x"20"),
  1423 => (x"20",x"20",x"20",x"00"),
  1424 => (x"20",x"20",x"20",x"20"),
  1425 => (x"6f",x"68",x"73",x"20"),
  1426 => (x"20",x"64",x"6c",x"75"),
  1427 => (x"20",x"3a",x"65",x"62"),
  1428 => (x"64",x"25",x"20",x"20"),
  1429 => (x"6e",x"45",x"00",x"0a"),
  1430 => (x"4c",x"5f",x"6d",x"75"),
  1431 => (x"20",x"3a",x"63",x"6f"),
  1432 => (x"20",x"20",x"20",x"20"),
  1433 => (x"20",x"20",x"20",x"20"),
  1434 => (x"25",x"20",x"20",x"20"),
  1435 => (x"20",x"00",x"0a",x"64"),
  1436 => (x"20",x"20",x"20",x"20"),
  1437 => (x"73",x"20",x"20",x"20"),
  1438 => (x"6c",x"75",x"6f",x"68"),
  1439 => (x"65",x"62",x"20",x"64"),
  1440 => (x"20",x"20",x"20",x"3a"),
  1441 => (x"00",x"0a",x"64",x"25"),
  1442 => (x"5f",x"72",x"74",x"53"),
  1443 => (x"6f",x"4c",x"5f",x"31"),
  1444 => (x"20",x"20",x"3a",x"63"),
  1445 => (x"20",x"20",x"20",x"20"),
  1446 => (x"20",x"20",x"20",x"20"),
  1447 => (x"0a",x"73",x"25",x"20"),
  1448 => (x"20",x"20",x"20",x"00"),
  1449 => (x"20",x"20",x"20",x"20"),
  1450 => (x"6f",x"68",x"73",x"20"),
  1451 => (x"20",x"64",x"6c",x"75"),
  1452 => (x"20",x"3a",x"65",x"62"),
  1453 => (x"48",x"44",x"20",x"20"),
  1454 => (x"54",x"53",x"59",x"52"),
  1455 => (x"20",x"45",x"4e",x"4f"),
  1456 => (x"47",x"4f",x"52",x"50"),
  1457 => (x"2c",x"4d",x"41",x"52"),
  1458 => (x"53",x"27",x"31",x"20"),
  1459 => (x"54",x"53",x"20",x"54"),
  1460 => (x"47",x"4e",x"49",x"52"),
  1461 => (x"74",x"53",x"00",x"0a"),
  1462 => (x"5f",x"32",x"5f",x"72"),
  1463 => (x"3a",x"63",x"6f",x"4c"),
  1464 => (x"20",x"20",x"20",x"20"),
  1465 => (x"20",x"20",x"20",x"20"),
  1466 => (x"25",x"20",x"20",x"20"),
  1467 => (x"20",x"00",x"0a",x"73"),
  1468 => (x"20",x"20",x"20",x"20"),
  1469 => (x"73",x"20",x"20",x"20"),
  1470 => (x"6c",x"75",x"6f",x"68"),
  1471 => (x"65",x"62",x"20",x"64"),
  1472 => (x"20",x"20",x"20",x"3a"),
  1473 => (x"59",x"52",x"48",x"44"),
  1474 => (x"4e",x"4f",x"54",x"53"),
  1475 => (x"52",x"50",x"20",x"45"),
  1476 => (x"41",x"52",x"47",x"4f"),
  1477 => (x"32",x"20",x"2c",x"4d"),
  1478 => (x"20",x"44",x"4e",x"27"),
  1479 => (x"49",x"52",x"54",x"53"),
  1480 => (x"00",x"0a",x"47",x"4e"),
  1481 => (x"73",x"55",x"00",x"0a"),
  1482 => (x"74",x"20",x"72",x"65"),
  1483 => (x"3a",x"65",x"6d",x"69"),
  1484 => (x"0a",x"64",x"25",x"20"),
  1485 => (x"00",x"00",x"00",x"00"),
  1486 => (x"00",x"00",x"00",x"00"),
  1487 => (x"00",x"00",x"61",x"a8"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
