
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"3b",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"38"),
    10 => (x"20",x"00",x"27",x"4f"),
    11 => (x"27",x"4e",x"00",x"00"),
    12 => (x"00",x"00",x"03",x"0f"),
    13 => (x"87",x"fd",x"00",x"0f"),
    14 => (x"4f",x"87",x"fd",x"00"),
    15 => (x"ff",x"86",x"fc",x"1e"),
    16 => (x"48",x"69",x"49",x"c0"),
    17 => (x"c4",x"98",x"c0",x"c4"),
    18 => (x"02",x"6e",x"58",x"a6"),
    19 => (x"66",x"c8",x"87",x"f4"),
    20 => (x"8e",x"fc",x"48",x"79"),
    21 => (x"73",x"1e",x"4f",x"26"),
    22 => (x"75",x"1e",x"74",x"1e"),
    23 => (x"c0",x"86",x"e4",x"1e"),
    24 => (x"c4",x"4d",x"66",x"f4"),
    25 => (x"78",x"c0",x"48",x"a6"),
    26 => (x"78",x"c0",x"80",x"c4"),
    27 => (x"97",x"66",x"ec",x"c0"),
    28 => (x"ec",x"c0",x"4b",x"bf"),
    29 => (x"80",x"c1",x"48",x"66"),
    30 => (x"58",x"a6",x"f0",x"c0"),
    31 => (x"c7",x"02",x"9b",x"73"),
    32 => (x"66",x"c8",x"87",x"e3"),
    33 => (x"87",x"f0",x"c6",x"02"),
    34 => (x"c0",x"48",x"a6",x"d0"),
    35 => (x"c0",x"80",x"f8",x"78"),
    36 => (x"ab",x"f0",x"c0",x"78"),
    37 => (x"87",x"e1",x"c2",x"02"),
    38 => (x"02",x"ab",x"e3",x"c1"),
    39 => (x"c1",x"87",x"e2",x"c2"),
    40 => (x"c0",x"02",x"ab",x"e4"),
    41 => (x"ec",x"c1",x"87",x"e2"),
    42 => (x"cc",x"c2",x"02",x"ab"),
    43 => (x"ab",x"f0",x"c1",x"87"),
    44 => (x"c1",x"87",x"dd",x"02"),
    45 => (x"df",x"02",x"ab",x"f3"),
    46 => (x"ab",x"f5",x"c1",x"87"),
    47 => (x"c1",x"87",x"c9",x"02"),
    48 => (x"cb",x"02",x"ab",x"f8"),
    49 => (x"87",x"de",x"c2",x"87"),
    50 => (x"ca",x"48",x"a6",x"d0"),
    51 => (x"87",x"f9",x"c2",x"78"),
    52 => (x"d0",x"48",x"a6",x"d0"),
    53 => (x"87",x"f1",x"c2",x"78"),
    54 => (x"48",x"66",x"f0",x"c0"),
    55 => (x"f4",x"c0",x"80",x"c4"),
    56 => (x"f0",x"c0",x"58",x"a6"),
    57 => (x"89",x"c4",x"49",x"66"),
    58 => (x"a6",x"d4",x"7e",x"69"),
    59 => (x"6e",x"78",x"ff",x"48"),
    60 => (x"dc",x"48",x"bf",x"97"),
    61 => (x"48",x"6e",x"58",x"a6"),
    62 => (x"a6",x"c4",x"80",x"c1"),
    63 => (x"5b",x"a6",x"d0",x"58"),
    64 => (x"c0",x"02",x"66",x"d8"),
    65 => (x"66",x"d8",x"87",x"e4"),
    66 => (x"d4",x"4b",x"6e",x"4c"),
    67 => (x"80",x"c1",x"48",x"66"),
    68 => (x"c0",x"58",x"a6",x"d8"),
    69 => (x"74",x"1e",x"66",x"f8"),
    70 => (x"c8",x"0f",x"75",x"1e"),
    71 => (x"05",x"a8",x"74",x"86"),
    72 => (x"4c",x"13",x"87",x"c8"),
    73 => (x"ff",x"05",x"9c",x"74"),
    74 => (x"66",x"cc",x"87",x"e1"),
    75 => (x"48",x"66",x"d4",x"4b"),
    76 => (x"c8",x"80",x"66",x"c4"),
    77 => (x"d0",x"c1",x"58",x"a6"),
    78 => (x"48",x"a6",x"c8",x"87"),
    79 => (x"c8",x"c1",x"78",x"c1"),
    80 => (x"66",x"f8",x"c0",x"87"),
    81 => (x"66",x"f4",x"c0",x"1e"),
    82 => (x"c0",x"80",x"c4",x"48"),
    83 => (x"c0",x"58",x"a6",x"f8"),
    84 => (x"c4",x"49",x"66",x"f4"),
    85 => (x"75",x"1e",x"69",x"89"),
    86 => (x"c4",x"86",x"c8",x"0f"),
    87 => (x"80",x"c1",x"48",x"66"),
    88 => (x"c0",x"58",x"a6",x"c8"),
    89 => (x"e5",x"c0",x"87",x"e3"),
    90 => (x"87",x"cb",x"02",x"ab"),
    91 => (x"1e",x"66",x"f8",x"c0"),
    92 => (x"75",x"1e",x"e5",x"c0"),
    93 => (x"c0",x"86",x"c8",x"0f"),
    94 => (x"73",x"1e",x"66",x"f8"),
    95 => (x"c8",x"0f",x"75",x"1e"),
    96 => (x"48",x"66",x"c4",x"86"),
    97 => (x"a6",x"c8",x"80",x"c1"),
    98 => (x"02",x"66",x"d0",x"58"),
    99 => (x"c0",x"87",x"c0",x"c3"),
   100 => (x"c4",x"48",x"66",x"f0"),
   101 => (x"a6",x"f4",x"c0",x"80"),
   102 => (x"66",x"f0",x"c0",x"58"),
   103 => (x"69",x"89",x"c4",x"49"),
   104 => (x"ab",x"e4",x"c1",x"7e"),
   105 => (x"6e",x"87",x"d8",x"05"),
   106 => (x"a8",x"b7",x"c0",x"48"),
   107 => (x"c0",x"87",x"d0",x"03"),
   108 => (x"c7",x"fa",x"1e",x"ed"),
   109 => (x"6e",x"86",x"c4",x"87"),
   110 => (x"88",x"08",x"c0",x"48"),
   111 => (x"6e",x"58",x"a6",x"c4"),
   112 => (x"ec",x"ce",x"c1",x"4a"),
   113 => (x"48",x"a6",x"cc",x"4c"),
   114 => (x"05",x"6e",x"78",x"c0"),
   115 => (x"ce",x"c1",x"87",x"ce"),
   116 => (x"ce",x"c1",x"4c",x"ed"),
   117 => (x"f0",x"c0",x"48",x"ec"),
   118 => (x"87",x"eb",x"c0",x"50"),
   119 => (x"e6",x"c0",x"02",x"6e"),
   120 => (x"4b",x"66",x"d0",x"87"),
   121 => (x"49",x"72",x"1e",x"72"),
   122 => (x"ec",x"c2",x"4a",x"73"),
   123 => (x"ca",x"4a",x"26",x"87"),
   124 => (x"54",x"11",x"81",x"c8"),
   125 => (x"49",x"72",x"1e",x"71"),
   126 => (x"dc",x"c2",x"4a",x"73"),
   127 => (x"26",x"4a",x"70",x"87"),
   128 => (x"05",x"9a",x"72",x"49"),
   129 => (x"c1",x"87",x"dd",x"ff"),
   130 => (x"02",x"ac",x"ec",x"ce"),
   131 => (x"f8",x"c0",x"87",x"df"),
   132 => (x"8c",x"c1",x"1e",x"66"),
   133 => (x"71",x"49",x"6c",x"97"),
   134 => (x"c8",x"0f",x"75",x"1e"),
   135 => (x"48",x"66",x"cc",x"86"),
   136 => (x"a6",x"d0",x"80",x"c1"),
   137 => (x"ec",x"ce",x"c1",x"58"),
   138 => (x"e1",x"ff",x"05",x"ac"),
   139 => (x"48",x"66",x"cc",x"87"),
   140 => (x"c8",x"80",x"66",x"c4"),
   141 => (x"87",x"d7",x"58",x"a6"),
   142 => (x"05",x"ab",x"e5",x"c0"),
   143 => (x"a6",x"c8",x"87",x"c7"),
   144 => (x"ca",x"78",x"c1",x"48"),
   145 => (x"66",x"f8",x"c0",x"87"),
   146 => (x"75",x"1e",x"73",x"1e"),
   147 => (x"c0",x"86",x"c8",x"0f"),
   148 => (x"bf",x"97",x"66",x"ec"),
   149 => (x"66",x"ec",x"c0",x"4b"),
   150 => (x"c0",x"80",x"c1",x"48"),
   151 => (x"73",x"58",x"a6",x"f0"),
   152 => (x"dd",x"f8",x"05",x"9b"),
   153 => (x"48",x"66",x"c4",x"87"),
   154 => (x"4d",x"26",x"8e",x"e4"),
   155 => (x"4b",x"26",x"4c",x"26"),
   156 => (x"c0",x"1e",x"4f",x"26"),
   157 => (x"1e",x"fc",x"c0",x"1e"),
   158 => (x"d0",x"1e",x"a6",x"d0"),
   159 => (x"d5",x"f7",x"1e",x"66"),
   160 => (x"26",x"86",x"d0",x"87"),
   161 => (x"00",x"00",x"00",x"4f"),
   162 => (x"33",x"32",x"31",x"30"),
   163 => (x"37",x"36",x"35",x"34"),
   164 => (x"42",x"41",x"39",x"38"),
   165 => (x"46",x"45",x"44",x"43"),
   166 => (x"1e",x"73",x"1e",x"00"),
   167 => (x"c0",x"02",x"9a",x"72"),
   168 => (x"48",x"c0",x"87",x"e7"),
   169 => (x"a9",x"72",x"4b",x"c1"),
   170 => (x"72",x"87",x"d1",x"06"),
   171 => (x"87",x"c9",x"06",x"82"),
   172 => (x"a9",x"72",x"83",x"73"),
   173 => (x"c3",x"87",x"f4",x"01"),
   174 => (x"3a",x"b2",x"c1",x"87"),
   175 => (x"89",x"03",x"a9",x"72"),
   176 => (x"c1",x"07",x"80",x"73"),
   177 => (x"f3",x"05",x"2b",x"2a"),
   178 => (x"26",x"4b",x"26",x"87"),
   179 => (x"1e",x"75",x"1e",x"4f"),
   180 => (x"b7",x"71",x"4d",x"c4"),
   181 => (x"b9",x"ff",x"04",x"a1"),
   182 => (x"bd",x"c3",x"81",x"c1"),
   183 => (x"a2",x"b7",x"72",x"07"),
   184 => (x"c1",x"ba",x"ff",x"04"),
   185 => (x"07",x"bd",x"c1",x"82"),
   186 => (x"c1",x"87",x"ee",x"fe"),
   187 => (x"b8",x"ff",x"04",x"2d"),
   188 => (x"2d",x"07",x"80",x"c1"),
   189 => (x"c1",x"b9",x"ff",x"04"),
   190 => (x"4d",x"26",x"07",x"81"),
   191 => (x"72",x"1e",x"4f",x"26"),
   192 => (x"11",x"48",x"12",x"1e"),
   193 => (x"88",x"87",x"c4",x"02"),
   194 => (x"26",x"87",x"f6",x"02"),
   195 => (x"1e",x"4f",x"26",x"4a"),
   196 => (x"1e",x"74",x"1e",x"73"),
   197 => (x"dc",x"ff",x"1e",x"75"),
   198 => (x"c0",x"cf",x"c1",x"86"),
   199 => (x"c4",x"ef",x"c3",x"48"),
   200 => (x"fc",x"ce",x"c1",x"78"),
   201 => (x"f4",x"ef",x"c3",x"48"),
   202 => (x"ef",x"c3",x"48",x"78"),
   203 => (x"ef",x"c3",x"78",x"c4"),
   204 => (x"78",x"c0",x"48",x"f8"),
   205 => (x"78",x"c2",x"80",x"c4"),
   206 => (x"48",x"c0",x"f0",x"c3"),
   207 => (x"71",x"78",x"e8",x"c0"),
   208 => (x"c4",x"f0",x"c3",x"1e"),
   209 => (x"d4",x"ed",x"c0",x"49"),
   210 => (x"20",x"41",x"20",x"48"),
   211 => (x"20",x"41",x"20",x"41"),
   212 => (x"20",x"41",x"20",x"41"),
   213 => (x"10",x"41",x"20",x"41"),
   214 => (x"10",x"51",x"10",x"51"),
   215 => (x"71",x"49",x"26",x"51"),
   216 => (x"e4",x"f0",x"c3",x"1e"),
   217 => (x"f4",x"ed",x"c0",x"49"),
   218 => (x"20",x"41",x"20",x"48"),
   219 => (x"20",x"41",x"20",x"41"),
   220 => (x"20",x"41",x"20",x"41"),
   221 => (x"10",x"41",x"20",x"41"),
   222 => (x"10",x"51",x"10",x"51"),
   223 => (x"c1",x"49",x"26",x"51"),
   224 => (x"ca",x"48",x"f8",x"eb"),
   225 => (x"d4",x"ee",x"c0",x"78"),
   226 => (x"87",x"e6",x"fb",x"1e"),
   227 => (x"ee",x"c0",x"86",x"c4"),
   228 => (x"dd",x"fb",x"1e",x"d8"),
   229 => (x"c0",x"86",x"c4",x"87"),
   230 => (x"fb",x"1e",x"c8",x"ef"),
   231 => (x"86",x"c4",x"87",x"d4"),
   232 => (x"bf",x"f8",x"e6",x"c0"),
   233 => (x"c0",x"87",x"d4",x"02"),
   234 => (x"fb",x"1e",x"c0",x"e7"),
   235 => (x"86",x"c4",x"87",x"c4"),
   236 => (x"1e",x"ec",x"e7",x"c0"),
   237 => (x"c4",x"87",x"fb",x"fa"),
   238 => (x"c0",x"87",x"d2",x"86"),
   239 => (x"fa",x"1e",x"f0",x"e7"),
   240 => (x"86",x"c4",x"87",x"f0"),
   241 => (x"1e",x"e0",x"e8",x"c0"),
   242 => (x"c4",x"87",x"e7",x"fa"),
   243 => (x"fc",x"e6",x"c0",x"86"),
   244 => (x"ef",x"c0",x"1e",x"bf"),
   245 => (x"d9",x"fa",x"1e",x"cc"),
   246 => (x"c3",x"86",x"c8",x"87"),
   247 => (x"ff",x"48",x"ec",x"ee"),
   248 => (x"c8",x"78",x"bf",x"c8"),
   249 => (x"78",x"c1",x"48",x"a6"),
   250 => (x"bf",x"fc",x"e6",x"c0"),
   251 => (x"a8",x"b7",x"c0",x"48"),
   252 => (x"87",x"f5",x"c8",x"06"),
   253 => (x"d4",x"48",x"a6",x"cc"),
   254 => (x"80",x"c8",x"58",x"a6"),
   255 => (x"dc",x"58",x"a6",x"dc"),
   256 => (x"a6",x"c8",x"48",x"a6"),
   257 => (x"cc",x"cf",x"c1",x"58"),
   258 => (x"50",x"c1",x"c1",x"48"),
   259 => (x"48",x"c8",x"cf",x"c1"),
   260 => (x"cf",x"c1",x"78",x"c0"),
   261 => (x"49",x"bf",x"97",x"cc"),
   262 => (x"02",x"a9",x"c1",x"c1"),
   263 => (x"c0",x"87",x"c5",x"c0"),
   264 => (x"87",x"c2",x"c0",x"7e"),
   265 => (x"cf",x"c1",x"7e",x"c1"),
   266 => (x"6e",x"48",x"bf",x"c8"),
   267 => (x"cc",x"cf",x"c1",x"b0"),
   268 => (x"d0",x"cf",x"c1",x"58"),
   269 => (x"50",x"c2",x"c1",x"48"),
   270 => (x"c2",x"48",x"a6",x"dc"),
   271 => (x"c3",x"80",x"c4",x"78"),
   272 => (x"c4",x"f1",x"c3",x"78"),
   273 => (x"c4",x"e9",x"c0",x"49"),
   274 => (x"20",x"41",x"20",x"48"),
   275 => (x"20",x"41",x"20",x"41"),
   276 => (x"20",x"41",x"20",x"41"),
   277 => (x"10",x"41",x"20",x"41"),
   278 => (x"10",x"51",x"10",x"51"),
   279 => (x"48",x"a6",x"d4",x"51"),
   280 => (x"f1",x"c3",x"78",x"c1"),
   281 => (x"f0",x"c3",x"1e",x"c4"),
   282 => (x"fb",x"c0",x"1e",x"e4"),
   283 => (x"86",x"c8",x"87",x"cc"),
   284 => (x"c0",x"05",x"98",x"70"),
   285 => (x"49",x"c1",x"87",x"c5"),
   286 => (x"c0",x"87",x"c2",x"c0"),
   287 => (x"cc",x"cf",x"c1",x"49"),
   288 => (x"48",x"66",x"dc",x"59"),
   289 => (x"03",x"a8",x"b7",x"c3"),
   290 => (x"dc",x"87",x"ee",x"c0"),
   291 => (x"91",x"c5",x"49",x"66"),
   292 => (x"88",x"c3",x"48",x"71"),
   293 => (x"d0",x"58",x"a6",x"d0"),
   294 => (x"1e",x"c3",x"1e",x"66"),
   295 => (x"1e",x"66",x"e4",x"c0"),
   296 => (x"87",x"c3",x"f7",x"c0"),
   297 => (x"66",x"dc",x"86",x"cc"),
   298 => (x"c0",x"80",x"c1",x"48"),
   299 => (x"dc",x"58",x"a6",x"e0"),
   300 => (x"b7",x"c3",x"48",x"66"),
   301 => (x"d2",x"ff",x"04",x"a8"),
   302 => (x"1e",x"66",x"cc",x"87"),
   303 => (x"1e",x"66",x"e0",x"c0"),
   304 => (x"1e",x"dc",x"d2",x"c1"),
   305 => (x"1e",x"d4",x"cf",x"c1"),
   306 => (x"87",x"ed",x"f6",x"c0"),
   307 => (x"ce",x"c1",x"86",x"d0"),
   308 => (x"c1",x"4c",x"bf",x"fc"),
   309 => (x"bf",x"bf",x"fc",x"ce"),
   310 => (x"73",x"1e",x"72",x"4b"),
   311 => (x"fc",x"ce",x"c1",x"49"),
   312 => (x"f0",x"c0",x"48",x"bf"),
   313 => (x"41",x"20",x"4a",x"a1"),
   314 => (x"ff",x"05",x"aa",x"71"),
   315 => (x"4a",x"26",x"87",x"f8"),
   316 => (x"cc",x"7e",x"a4",x"c8"),
   317 => (x"79",x"c5",x"49",x"a4"),
   318 => (x"69",x"4d",x"a3",x"cc"),
   319 => (x"73",x"7b",x"6c",x"7d"),
   320 => (x"87",x"c9",x"d2",x"1e"),
   321 => (x"a3",x"c4",x"86",x"c4"),
   322 => (x"c0",x"05",x"69",x"49"),
   323 => (x"a3",x"c8",x"87",x"e6"),
   324 => (x"71",x"7d",x"c6",x"49"),
   325 => (x"bf",x"66",x"c4",x"1e"),
   326 => (x"ee",x"f3",x"c0",x"1e"),
   327 => (x"c1",x"86",x"c8",x"87"),
   328 => (x"bf",x"bf",x"fc",x"ce"),
   329 => (x"ca",x"1e",x"75",x"7b"),
   330 => (x"c0",x"1e",x"6d",x"1e"),
   331 => (x"cc",x"87",x"f8",x"f4"),
   332 => (x"87",x"d9",x"c0",x"86"),
   333 => (x"1e",x"71",x"49",x"6c"),
   334 => (x"49",x"74",x"1e",x"72"),
   335 => (x"a1",x"f0",x"c0",x"48"),
   336 => (x"71",x"41",x"20",x"4a"),
   337 => (x"f8",x"ff",x"05",x"aa"),
   338 => (x"26",x"4a",x"26",x"87"),
   339 => (x"97",x"c1",x"c1",x"49"),
   340 => (x"d0",x"cf",x"c1",x"7e"),
   341 => (x"c1",x"49",x"bf",x"97"),
   342 => (x"04",x"a9",x"b7",x"c1"),
   343 => (x"97",x"87",x"e1",x"c1"),
   344 => (x"c3",x"c1",x"4b",x"6e"),
   345 => (x"71",x"49",x"73",x"1e"),
   346 => (x"eb",x"f6",x"c0",x"1e"),
   347 => (x"d4",x"86",x"c8",x"87"),
   348 => (x"c0",x"05",x"a8",x"66"),
   349 => (x"66",x"d8",x"87",x"f9"),
   350 => (x"c0",x"1e",x"c0",x"1e"),
   351 => (x"c8",x"87",x"cc",x"f2"),
   352 => (x"c3",x"1e",x"71",x"86"),
   353 => (x"c0",x"49",x"c4",x"f1"),
   354 => (x"20",x"48",x"e4",x"e8"),
   355 => (x"20",x"41",x"20",x"41"),
   356 => (x"20",x"41",x"20",x"41"),
   357 => (x"20",x"41",x"20",x"41"),
   358 => (x"10",x"51",x"10",x"41"),
   359 => (x"26",x"51",x"10",x"51"),
   360 => (x"a6",x"e0",x"c0",x"49"),
   361 => (x"78",x"66",x"c8",x"48"),
   362 => (x"48",x"c4",x"cf",x"c1"),
   363 => (x"c1",x"78",x"66",x"c8"),
   364 => (x"c1",x"4a",x"73",x"83"),
   365 => (x"bf",x"97",x"d0",x"cf"),
   366 => (x"aa",x"b7",x"71",x"49"),
   367 => (x"87",x"e2",x"fe",x"06"),
   368 => (x"48",x"66",x"e0",x"c0"),
   369 => (x"c0",x"90",x"66",x"dc"),
   370 => (x"71",x"58",x"a6",x"e4"),
   371 => (x"c0",x"1e",x"72",x"1e"),
   372 => (x"d4",x"49",x"66",x"e8"),
   373 => (x"f4",x"f3",x"4a",x"66"),
   374 => (x"26",x"4a",x"26",x"87"),
   375 => (x"a6",x"e0",x"c0",x"49"),
   376 => (x"66",x"e0",x"c0",x"58"),
   377 => (x"89",x"66",x"cc",x"49"),
   378 => (x"48",x"71",x"91",x"c7"),
   379 => (x"c0",x"88",x"66",x"dc"),
   380 => (x"c4",x"58",x"a6",x"e4"),
   381 => (x"ca",x"4a",x"bf",x"66"),
   382 => (x"cc",x"cf",x"c1",x"82"),
   383 => (x"c1",x"49",x"bf",x"97"),
   384 => (x"c0",x"05",x"a9",x"c1"),
   385 => (x"8a",x"c1",x"87",x"ce"),
   386 => (x"cf",x"c1",x"48",x"72"),
   387 => (x"c4",x"88",x"bf",x"c4"),
   388 => (x"08",x"78",x"08",x"66"),
   389 => (x"c1",x"48",x"66",x"c8"),
   390 => (x"58",x"a6",x"cc",x"80"),
   391 => (x"c0",x"48",x"66",x"c8"),
   392 => (x"b7",x"bf",x"fc",x"e6"),
   393 => (x"dc",x"f7",x"06",x"a8"),
   394 => (x"f0",x"ee",x"c3",x"87"),
   395 => (x"bf",x"c8",x"ff",x"48"),
   396 => (x"fc",x"ef",x"c0",x"78"),
   397 => (x"87",x"fa",x"f0",x"1e"),
   398 => (x"f0",x"c0",x"86",x"c4"),
   399 => (x"f1",x"f0",x"1e",x"cc"),
   400 => (x"c0",x"86",x"c4",x"87"),
   401 => (x"f0",x"1e",x"d0",x"f0"),
   402 => (x"86",x"c4",x"87",x"e8"),
   403 => (x"1e",x"c8",x"f1",x"c0"),
   404 => (x"c4",x"87",x"df",x"f0"),
   405 => (x"c4",x"cf",x"c1",x"86"),
   406 => (x"f1",x"c0",x"1e",x"bf"),
   407 => (x"d1",x"f0",x"1e",x"cc"),
   408 => (x"c5",x"86",x"c8",x"87"),
   409 => (x"e8",x"f1",x"c0",x"1e"),
   410 => (x"87",x"c6",x"f0",x"1e"),
   411 => (x"cf",x"c1",x"86",x"c8"),
   412 => (x"c0",x"1e",x"bf",x"c8"),
   413 => (x"ef",x"1e",x"c4",x"f2"),
   414 => (x"86",x"c8",x"87",x"f8"),
   415 => (x"f2",x"c0",x"1e",x"c1"),
   416 => (x"ed",x"ef",x"1e",x"e0"),
   417 => (x"c1",x"86",x"c8",x"87"),
   418 => (x"bf",x"97",x"cc",x"cf"),
   419 => (x"c0",x"1e",x"71",x"49"),
   420 => (x"ef",x"1e",x"fc",x"f2"),
   421 => (x"86",x"c8",x"87",x"dc"),
   422 => (x"c0",x"1e",x"c1",x"c1"),
   423 => (x"ef",x"1e",x"d8",x"f3"),
   424 => (x"86",x"c8",x"87",x"d0"),
   425 => (x"97",x"d0",x"cf",x"c1"),
   426 => (x"1e",x"71",x"49",x"bf"),
   427 => (x"1e",x"f4",x"f3",x"c0"),
   428 => (x"c8",x"87",x"ff",x"ee"),
   429 => (x"1e",x"c2",x"c1",x"86"),
   430 => (x"1e",x"d0",x"f4",x"c0"),
   431 => (x"c8",x"87",x"f3",x"ee"),
   432 => (x"f4",x"cf",x"c1",x"86"),
   433 => (x"f4",x"c0",x"1e",x"bf"),
   434 => (x"e5",x"ee",x"1e",x"ec"),
   435 => (x"c7",x"86",x"c8",x"87"),
   436 => (x"c8",x"f5",x"c0",x"1e"),
   437 => (x"87",x"da",x"ee",x"1e"),
   438 => (x"eb",x"c1",x"86",x"c8"),
   439 => (x"c0",x"1e",x"bf",x"f8"),
   440 => (x"ee",x"1e",x"e4",x"f5"),
   441 => (x"86",x"c8",x"87",x"cc"),
   442 => (x"1e",x"c0",x"f6",x"c0"),
   443 => (x"c4",x"87",x"c3",x"ee"),
   444 => (x"ec",x"f6",x"c0",x"86"),
   445 => (x"87",x"fa",x"ed",x"1e"),
   446 => (x"ce",x"c1",x"86",x"c4"),
   447 => (x"1e",x"bf",x"bf",x"fc"),
   448 => (x"1e",x"f8",x"f6",x"c0"),
   449 => (x"c8",x"87",x"eb",x"ed"),
   450 => (x"d4",x"f7",x"c0",x"86"),
   451 => (x"87",x"e2",x"ed",x"1e"),
   452 => (x"ce",x"c1",x"86",x"c4"),
   453 => (x"c4",x"49",x"bf",x"fc"),
   454 => (x"c0",x"1e",x"69",x"81"),
   455 => (x"ed",x"1e",x"c8",x"f8"),
   456 => (x"86",x"c8",x"87",x"d0"),
   457 => (x"f8",x"c0",x"1e",x"c0"),
   458 => (x"c5",x"ed",x"1e",x"e4"),
   459 => (x"c1",x"86",x"c8",x"87"),
   460 => (x"49",x"bf",x"fc",x"ce"),
   461 => (x"1e",x"69",x"81",x"c8"),
   462 => (x"1e",x"c0",x"f9",x"c0"),
   463 => (x"c8",x"87",x"f3",x"ec"),
   464 => (x"c0",x"1e",x"c2",x"86"),
   465 => (x"ec",x"1e",x"dc",x"f9"),
   466 => (x"86",x"c8",x"87",x"e8"),
   467 => (x"bf",x"fc",x"ce",x"c1"),
   468 => (x"69",x"81",x"cc",x"49"),
   469 => (x"f8",x"f9",x"c0",x"1e"),
   470 => (x"87",x"d6",x"ec",x"1e"),
   471 => (x"1e",x"d1",x"86",x"c8"),
   472 => (x"1e",x"d4",x"fa",x"c0"),
   473 => (x"c8",x"87",x"cb",x"ec"),
   474 => (x"fc",x"ce",x"c1",x"86"),
   475 => (x"81",x"d0",x"49",x"bf"),
   476 => (x"fa",x"c0",x"1e",x"71"),
   477 => (x"f9",x"eb",x"1e",x"f0"),
   478 => (x"c0",x"86",x"c8",x"87"),
   479 => (x"eb",x"1e",x"cc",x"fb"),
   480 => (x"86",x"c4",x"87",x"f0"),
   481 => (x"1e",x"c4",x"fc",x"c0"),
   482 => (x"c4",x"87",x"e7",x"eb"),
   483 => (x"c0",x"cf",x"c1",x"86"),
   484 => (x"c0",x"1e",x"bf",x"bf"),
   485 => (x"eb",x"1e",x"d8",x"fc"),
   486 => (x"86",x"c8",x"87",x"d8"),
   487 => (x"1e",x"f4",x"fc",x"c0"),
   488 => (x"c4",x"87",x"cf",x"eb"),
   489 => (x"c0",x"cf",x"c1",x"86"),
   490 => (x"81",x"c4",x"49",x"bf"),
   491 => (x"fd",x"c0",x"1e",x"69"),
   492 => (x"fd",x"ea",x"1e",x"f4"),
   493 => (x"c0",x"86",x"c8",x"87"),
   494 => (x"d0",x"fe",x"c0",x"1e"),
   495 => (x"87",x"f2",x"ea",x"1e"),
   496 => (x"cf",x"c1",x"86",x"c8"),
   497 => (x"c8",x"49",x"bf",x"c0"),
   498 => (x"c0",x"1e",x"69",x"81"),
   499 => (x"ea",x"1e",x"ec",x"fe"),
   500 => (x"86",x"c8",x"87",x"e0"),
   501 => (x"ff",x"c0",x"1e",x"c1"),
   502 => (x"d5",x"ea",x"1e",x"c8"),
   503 => (x"c1",x"86",x"c8",x"87"),
   504 => (x"49",x"bf",x"c0",x"cf"),
   505 => (x"1e",x"69",x"81",x"cc"),
   506 => (x"1e",x"e4",x"ff",x"c0"),
   507 => (x"c8",x"87",x"c3",x"ea"),
   508 => (x"c1",x"1e",x"d2",x"86"),
   509 => (x"e9",x"1e",x"c0",x"c0"),
   510 => (x"86",x"c8",x"87",x"f8"),
   511 => (x"bf",x"c0",x"cf",x"c1"),
   512 => (x"71",x"81",x"d0",x"49"),
   513 => (x"dc",x"c0",x"c1",x"1e"),
   514 => (x"87",x"e6",x"e9",x"1e"),
   515 => (x"c0",x"c1",x"86",x"c8"),
   516 => (x"dd",x"e9",x"1e",x"f8"),
   517 => (x"dc",x"86",x"c4",x"87"),
   518 => (x"c1",x"c1",x"1e",x"66"),
   519 => (x"d1",x"e9",x"1e",x"f0"),
   520 => (x"c5",x"86",x"c8",x"87"),
   521 => (x"cc",x"c2",x"c1",x"1e"),
   522 => (x"87",x"c6",x"e9",x"1e"),
   523 => (x"e0",x"c0",x"86",x"c8"),
   524 => (x"c2",x"c1",x"1e",x"66"),
   525 => (x"f9",x"e8",x"1e",x"e8"),
   526 => (x"cd",x"86",x"c8",x"87"),
   527 => (x"c4",x"c3",x"c1",x"1e"),
   528 => (x"87",x"ee",x"e8",x"1e"),
   529 => (x"66",x"cc",x"86",x"c8"),
   530 => (x"e0",x"c3",x"c1",x"1e"),
   531 => (x"87",x"e2",x"e8",x"1e"),
   532 => (x"1e",x"c7",x"86",x"c8"),
   533 => (x"1e",x"fc",x"c3",x"c1"),
   534 => (x"c8",x"87",x"d7",x"e8"),
   535 => (x"1e",x"66",x"d4",x"86"),
   536 => (x"1e",x"d8",x"c4",x"c1"),
   537 => (x"c8",x"87",x"cb",x"e8"),
   538 => (x"c1",x"1e",x"c1",x"86"),
   539 => (x"e8",x"1e",x"f4",x"c4"),
   540 => (x"86",x"c8",x"87",x"c0"),
   541 => (x"1e",x"e4",x"f0",x"c3"),
   542 => (x"1e",x"d0",x"c5",x"c1"),
   543 => (x"c8",x"87",x"f3",x"e7"),
   544 => (x"ec",x"c5",x"c1",x"86"),
   545 => (x"87",x"ea",x"e7",x"1e"),
   546 => (x"f1",x"c3",x"86",x"c4"),
   547 => (x"c6",x"c1",x"1e",x"c4"),
   548 => (x"dd",x"e7",x"1e",x"e4"),
   549 => (x"c1",x"86",x"c8",x"87"),
   550 => (x"e7",x"1e",x"c0",x"c7"),
   551 => (x"86",x"c4",x"87",x"d4"),
   552 => (x"1e",x"f8",x"c7",x"c1"),
   553 => (x"c4",x"87",x"cb",x"e7"),
   554 => (x"f0",x"ee",x"c3",x"86"),
   555 => (x"ee",x"c3",x"49",x"bf"),
   556 => (x"c3",x"89",x"bf",x"ec"),
   557 => (x"71",x"59",x"f8",x"ee"),
   558 => (x"fc",x"c7",x"c1",x"1e"),
   559 => (x"87",x"f2",x"e6",x"1e"),
   560 => (x"ee",x"c3",x"86",x"c8"),
   561 => (x"c1",x"48",x"bf",x"f4"),
   562 => (x"03",x"a8",x"b7",x"f8"),
   563 => (x"c0",x"87",x"db",x"c0"),
   564 => (x"e6",x"1e",x"e4",x"e9"),
   565 => (x"86",x"c4",x"87",x"dc"),
   566 => (x"1e",x"dc",x"ea",x"c0"),
   567 => (x"c4",x"87",x"d3",x"e6"),
   568 => (x"fc",x"ea",x"c0",x"86"),
   569 => (x"87",x"ca",x"e6",x"1e"),
   570 => (x"ee",x"c3",x"86",x"c4"),
   571 => (x"71",x"49",x"bf",x"f4"),
   572 => (x"92",x"e8",x"cf",x"4a"),
   573 => (x"1e",x"72",x"1e",x"71"),
   574 => (x"e6",x"c0",x"49",x"72"),
   575 => (x"e7",x"4a",x"bf",x"fc"),
   576 => (x"4a",x"26",x"87",x"cb"),
   577 => (x"ee",x"c3",x"49",x"26"),
   578 => (x"e6",x"c0",x"58",x"fc"),
   579 => (x"72",x"4a",x"bf",x"fc"),
   580 => (x"93",x"e8",x"cf",x"4b"),
   581 => (x"1e",x"72",x"1e",x"71"),
   582 => (x"e6",x"4a",x"09",x"73"),
   583 => (x"4a",x"26",x"87",x"ef"),
   584 => (x"ef",x"c3",x"49",x"26"),
   585 => (x"f9",x"c8",x"58",x"c0"),
   586 => (x"72",x"1e",x"71",x"92"),
   587 => (x"4a",x"09",x"72",x"1e"),
   588 => (x"26",x"87",x"da",x"e6"),
   589 => (x"c3",x"49",x"26",x"4a"),
   590 => (x"c0",x"58",x"c4",x"ef"),
   591 => (x"e4",x"1e",x"c0",x"eb"),
   592 => (x"86",x"c4",x"87",x"f0"),
   593 => (x"bf",x"f8",x"ee",x"c3"),
   594 => (x"f0",x"eb",x"c0",x"1e"),
   595 => (x"87",x"e2",x"e4",x"1e"),
   596 => (x"eb",x"c0",x"86",x"c8"),
   597 => (x"d9",x"e4",x"1e",x"f8"),
   598 => (x"c3",x"86",x"c4",x"87"),
   599 => (x"1e",x"bf",x"fc",x"ee"),
   600 => (x"1e",x"e8",x"ec",x"c0"),
   601 => (x"c8",x"87",x"cb",x"e4"),
   602 => (x"c0",x"ef",x"c3",x"86"),
   603 => (x"ec",x"c0",x"1e",x"bf"),
   604 => (x"fd",x"e3",x"1e",x"f0"),
   605 => (x"c0",x"86",x"c8",x"87"),
   606 => (x"e3",x"1e",x"d0",x"ed"),
   607 => (x"86",x"c4",x"87",x"f4"),
   608 => (x"dc",x"ff",x"48",x"c0"),
   609 => (x"26",x"4d",x"26",x"8e"),
   610 => (x"26",x"4b",x"26",x"4c"),
   611 => (x"ce",x"c1",x"1e",x"4f"),
   612 => (x"c9",x"02",x"bf",x"fc"),
   613 => (x"48",x"66",x"c4",x"87"),
   614 => (x"bf",x"fc",x"ce",x"c1"),
   615 => (x"ce",x"c1",x"78",x"bf"),
   616 => (x"cc",x"49",x"bf",x"fc"),
   617 => (x"c1",x"1e",x"71",x"81"),
   618 => (x"1e",x"bf",x"c4",x"cf"),
   619 => (x"e2",x"c0",x"1e",x"ca"),
   620 => (x"86",x"cc",x"87",x"f5"),
   621 => (x"00",x"00",x"4f",x"26"),
   622 => (x"00",x"00",x"00",x"00"),
   623 => (x"00",x"00",x"61",x"a8"),
   624 => (x"67",x"6f",x"72",x"50"),
   625 => (x"20",x"6d",x"61",x"72"),
   626 => (x"70",x"6d",x"6f",x"63"),
   627 => (x"64",x"65",x"6c",x"69"),
   628 => (x"74",x"69",x"77",x"20"),
   629 => (x"72",x"27",x"20",x"68"),
   630 => (x"73",x"69",x"67",x"65"),
   631 => (x"27",x"72",x"65",x"74"),
   632 => (x"74",x"74",x"61",x"20"),
   633 => (x"75",x"62",x"69",x"72"),
   634 => (x"00",x"0a",x"65",x"74"),
   635 => (x"00",x"00",x"00",x"0a"),
   636 => (x"67",x"6f",x"72",x"50"),
   637 => (x"20",x"6d",x"61",x"72"),
   638 => (x"70",x"6d",x"6f",x"63"),
   639 => (x"64",x"65",x"6c",x"69"),
   640 => (x"74",x"69",x"77",x"20"),
   641 => (x"74",x"75",x"6f",x"68"),
   642 => (x"65",x"72",x"27",x"20"),
   643 => (x"74",x"73",x"69",x"67"),
   644 => (x"20",x"27",x"72",x"65"),
   645 => (x"72",x"74",x"74",x"61"),
   646 => (x"74",x"75",x"62",x"69"),
   647 => (x"00",x"00",x"0a",x"65"),
   648 => (x"00",x"00",x"00",x"0a"),
   649 => (x"59",x"52",x"48",x"44"),
   650 => (x"4e",x"4f",x"54",x"53"),
   651 => (x"52",x"50",x"20",x"45"),
   652 => (x"41",x"52",x"47",x"4f"),
   653 => (x"33",x"20",x"2c",x"4d"),
   654 => (x"20",x"44",x"52",x"27"),
   655 => (x"49",x"52",x"54",x"53"),
   656 => (x"00",x"00",x"47",x"4e"),
   657 => (x"59",x"52",x"48",x"44"),
   658 => (x"4e",x"4f",x"54",x"53"),
   659 => (x"52",x"50",x"20",x"45"),
   660 => (x"41",x"52",x"47",x"4f"),
   661 => (x"32",x"20",x"2c",x"4d"),
   662 => (x"20",x"44",x"4e",x"27"),
   663 => (x"49",x"52",x"54",x"53"),
   664 => (x"00",x"00",x"47",x"4e"),
   665 => (x"73",x"61",x"65",x"4d"),
   666 => (x"64",x"65",x"72",x"75"),
   667 => (x"6d",x"69",x"74",x"20"),
   668 => (x"6f",x"74",x"20",x"65"),
   669 => (x"6d",x"73",x"20",x"6f"),
   670 => (x"20",x"6c",x"6c",x"61"),
   671 => (x"6f",x"20",x"6f",x"74"),
   672 => (x"69",x"61",x"74",x"62"),
   673 => (x"65",x"6d",x"20",x"6e"),
   674 => (x"6e",x"69",x"6e",x"61"),
   675 => (x"6c",x"75",x"66",x"67"),
   676 => (x"73",x"65",x"72",x"20"),
   677 => (x"73",x"74",x"6c",x"75"),
   678 => (x"00",x"00",x"00",x"0a"),
   679 => (x"61",x"65",x"6c",x"50"),
   680 => (x"69",x"20",x"65",x"73"),
   681 => (x"65",x"72",x"63",x"6e"),
   682 => (x"20",x"65",x"73",x"61"),
   683 => (x"62",x"6d",x"75",x"6e"),
   684 => (x"6f",x"20",x"72",x"65"),
   685 => (x"75",x"72",x"20",x"66"),
   686 => (x"00",x"0a",x"73",x"6e"),
   687 => (x"00",x"00",x"00",x"0a"),
   688 => (x"72",x"63",x"69",x"4d"),
   689 => (x"63",x"65",x"73",x"6f"),
   690 => (x"73",x"64",x"6e",x"6f"),
   691 => (x"72",x"6f",x"66",x"20"),
   692 => (x"65",x"6e",x"6f",x"20"),
   693 => (x"6e",x"75",x"72",x"20"),
   694 => (x"72",x"68",x"74",x"20"),
   695 => (x"68",x"67",x"75",x"6f"),
   696 => (x"72",x"68",x"44",x"20"),
   697 => (x"6f",x"74",x"73",x"79"),
   698 => (x"20",x"3a",x"65",x"6e"),
   699 => (x"00",x"00",x"00",x"00"),
   700 => (x"0a",x"20",x"64",x"25"),
   701 => (x"00",x"00",x"00",x"00"),
   702 => (x"79",x"72",x"68",x"44"),
   703 => (x"6e",x"6f",x"74",x"73"),
   704 => (x"70",x"20",x"73",x"65"),
   705 => (x"53",x"20",x"72",x"65"),
   706 => (x"6e",x"6f",x"63",x"65"),
   707 => (x"20",x"20",x"3a",x"64"),
   708 => (x"20",x"20",x"20",x"20"),
   709 => (x"20",x"20",x"20",x"20"),
   710 => (x"20",x"20",x"20",x"20"),
   711 => (x"20",x"20",x"20",x"20"),
   712 => (x"20",x"20",x"20",x"20"),
   713 => (x"00",x"00",x"00",x"00"),
   714 => (x"0a",x"20",x"64",x"25"),
   715 => (x"00",x"00",x"00",x"00"),
   716 => (x"20",x"58",x"41",x"56"),
   717 => (x"53",x"50",x"49",x"4d"),
   718 => (x"74",x"61",x"72",x"20"),
   719 => (x"20",x"67",x"6e",x"69"),
   720 => (x"30",x"31",x"20",x"2a"),
   721 => (x"3d",x"20",x"30",x"30"),
   722 => (x"20",x"64",x"25",x"20"),
   723 => (x"00",x"00",x"00",x"0a"),
   724 => (x"00",x"00",x"00",x"0a"),
   725 => (x"59",x"52",x"48",x"44"),
   726 => (x"4e",x"4f",x"54",x"53"),
   727 => (x"52",x"50",x"20",x"45"),
   728 => (x"41",x"52",x"47",x"4f"),
   729 => (x"53",x"20",x"2c",x"4d"),
   730 => (x"20",x"45",x"4d",x"4f"),
   731 => (x"49",x"52",x"54",x"53"),
   732 => (x"00",x"00",x"47",x"4e"),
   733 => (x"59",x"52",x"48",x"44"),
   734 => (x"4e",x"4f",x"54",x"53"),
   735 => (x"52",x"50",x"20",x"45"),
   736 => (x"41",x"52",x"47",x"4f"),
   737 => (x"31",x"20",x"2c",x"4d"),
   738 => (x"20",x"54",x"53",x"27"),
   739 => (x"49",x"52",x"54",x"53"),
   740 => (x"00",x"00",x"47",x"4e"),
   741 => (x"00",x"00",x"00",x"0a"),
   742 => (x"79",x"72",x"68",x"44"),
   743 => (x"6e",x"6f",x"74",x"73"),
   744 => (x"65",x"42",x"20",x"65"),
   745 => (x"6d",x"68",x"63",x"6e"),
   746 => (x"2c",x"6b",x"72",x"61"),
   747 => (x"72",x"65",x"56",x"20"),
   748 => (x"6e",x"6f",x"69",x"73"),
   749 => (x"31",x"2e",x"32",x"20"),
   750 => (x"61",x"4c",x"28",x"20"),
   751 => (x"61",x"75",x"67",x"6e"),
   752 => (x"20",x"3a",x"65",x"67"),
   753 => (x"00",x"0a",x"29",x"43"),
   754 => (x"00",x"00",x"00",x"0a"),
   755 => (x"63",x"65",x"78",x"45"),
   756 => (x"6f",x"69",x"74",x"75"),
   757 => (x"74",x"73",x"20",x"6e"),
   758 => (x"73",x"74",x"72",x"61"),
   759 => (x"64",x"25",x"20",x"2c"),
   760 => (x"6e",x"75",x"72",x"20"),
   761 => (x"68",x"74",x"20",x"73"),
   762 => (x"67",x"75",x"6f",x"72"),
   763 => (x"68",x"44",x"20",x"68"),
   764 => (x"74",x"73",x"79",x"72"),
   765 => (x"0a",x"65",x"6e",x"6f"),
   766 => (x"00",x"00",x"00",x"00"),
   767 => (x"63",x"65",x"78",x"45"),
   768 => (x"6f",x"69",x"74",x"75"),
   769 => (x"6e",x"65",x"20",x"6e"),
   770 => (x"00",x"0a",x"73",x"64"),
   771 => (x"00",x"00",x"00",x"0a"),
   772 => (x"61",x"6e",x"69",x"46"),
   773 => (x"61",x"76",x"20",x"6c"),
   774 => (x"73",x"65",x"75",x"6c"),
   775 => (x"20",x"66",x"6f",x"20"),
   776 => (x"20",x"65",x"68",x"74"),
   777 => (x"69",x"72",x"61",x"76"),
   778 => (x"65",x"6c",x"62",x"61"),
   779 => (x"73",x"75",x"20",x"73"),
   780 => (x"69",x"20",x"64",x"65"),
   781 => (x"68",x"74",x"20",x"6e"),
   782 => (x"65",x"62",x"20",x"65"),
   783 => (x"6d",x"68",x"63",x"6e"),
   784 => (x"3a",x"6b",x"72",x"61"),
   785 => (x"00",x"00",x"00",x"0a"),
   786 => (x"00",x"00",x"00",x"0a"),
   787 => (x"5f",x"74",x"6e",x"49"),
   788 => (x"62",x"6f",x"6c",x"47"),
   789 => (x"20",x"20",x"20",x"3a"),
   790 => (x"20",x"20",x"20",x"20"),
   791 => (x"20",x"20",x"20",x"20"),
   792 => (x"0a",x"64",x"25",x"20"),
   793 => (x"00",x"00",x"00",x"00"),
   794 => (x"20",x"20",x"20",x"20"),
   795 => (x"20",x"20",x"20",x"20"),
   796 => (x"75",x"6f",x"68",x"73"),
   797 => (x"62",x"20",x"64",x"6c"),
   798 => (x"20",x"20",x"3a",x"65"),
   799 => (x"0a",x"64",x"25",x"20"),
   800 => (x"00",x"00",x"00",x"00"),
   801 => (x"6c",x"6f",x"6f",x"42"),
   802 => (x"6f",x"6c",x"47",x"5f"),
   803 => (x"20",x"20",x"3a",x"62"),
   804 => (x"20",x"20",x"20",x"20"),
   805 => (x"20",x"20",x"20",x"20"),
   806 => (x"0a",x"64",x"25",x"20"),
   807 => (x"00",x"00",x"00",x"00"),
   808 => (x"20",x"20",x"20",x"20"),
   809 => (x"20",x"20",x"20",x"20"),
   810 => (x"75",x"6f",x"68",x"73"),
   811 => (x"62",x"20",x"64",x"6c"),
   812 => (x"20",x"20",x"3a",x"65"),
   813 => (x"0a",x"64",x"25",x"20"),
   814 => (x"00",x"00",x"00",x"00"),
   815 => (x"31",x"5f",x"68",x"43"),
   816 => (x"6f",x"6c",x"47",x"5f"),
   817 => (x"20",x"20",x"3a",x"62"),
   818 => (x"20",x"20",x"20",x"20"),
   819 => (x"20",x"20",x"20",x"20"),
   820 => (x"0a",x"63",x"25",x"20"),
   821 => (x"00",x"00",x"00",x"00"),
   822 => (x"20",x"20",x"20",x"20"),
   823 => (x"20",x"20",x"20",x"20"),
   824 => (x"75",x"6f",x"68",x"73"),
   825 => (x"62",x"20",x"64",x"6c"),
   826 => (x"20",x"20",x"3a",x"65"),
   827 => (x"0a",x"63",x"25",x"20"),
   828 => (x"00",x"00",x"00",x"00"),
   829 => (x"32",x"5f",x"68",x"43"),
   830 => (x"6f",x"6c",x"47",x"5f"),
   831 => (x"20",x"20",x"3a",x"62"),
   832 => (x"20",x"20",x"20",x"20"),
   833 => (x"20",x"20",x"20",x"20"),
   834 => (x"0a",x"63",x"25",x"20"),
   835 => (x"00",x"00",x"00",x"00"),
   836 => (x"20",x"20",x"20",x"20"),
   837 => (x"20",x"20",x"20",x"20"),
   838 => (x"75",x"6f",x"68",x"73"),
   839 => (x"62",x"20",x"64",x"6c"),
   840 => (x"20",x"20",x"3a",x"65"),
   841 => (x"0a",x"63",x"25",x"20"),
   842 => (x"00",x"00",x"00",x"00"),
   843 => (x"5f",x"72",x"72",x"41"),
   844 => (x"6c",x"47",x"5f",x"31"),
   845 => (x"38",x"5b",x"62",x"6f"),
   846 => (x"20",x"20",x"3a",x"5d"),
   847 => (x"20",x"20",x"20",x"20"),
   848 => (x"0a",x"64",x"25",x"20"),
   849 => (x"00",x"00",x"00",x"00"),
   850 => (x"20",x"20",x"20",x"20"),
   851 => (x"20",x"20",x"20",x"20"),
   852 => (x"75",x"6f",x"68",x"73"),
   853 => (x"62",x"20",x"64",x"6c"),
   854 => (x"20",x"20",x"3a",x"65"),
   855 => (x"0a",x"64",x"25",x"20"),
   856 => (x"00",x"00",x"00",x"00"),
   857 => (x"5f",x"72",x"72",x"41"),
   858 => (x"6c",x"47",x"5f",x"32"),
   859 => (x"38",x"5b",x"62",x"6f"),
   860 => (x"5d",x"37",x"5b",x"5d"),
   861 => (x"20",x"20",x"20",x"3a"),
   862 => (x"0a",x"64",x"25",x"20"),
   863 => (x"00",x"00",x"00",x"00"),
   864 => (x"20",x"20",x"20",x"20"),
   865 => (x"20",x"20",x"20",x"20"),
   866 => (x"75",x"6f",x"68",x"73"),
   867 => (x"62",x"20",x"64",x"6c"),
   868 => (x"20",x"20",x"3a",x"65"),
   869 => (x"6d",x"75",x"4e",x"20"),
   870 => (x"5f",x"72",x"65",x"62"),
   871 => (x"52",x"5f",x"66",x"4f"),
   872 => (x"20",x"73",x"6e",x"75"),
   873 => (x"30",x"31",x"20",x"2b"),
   874 => (x"00",x"00",x"00",x"0a"),
   875 => (x"5f",x"72",x"74",x"50"),
   876 => (x"62",x"6f",x"6c",x"47"),
   877 => (x"00",x"0a",x"3e",x"2d"),
   878 => (x"74",x"50",x"20",x"20"),
   879 => (x"6f",x"43",x"5f",x"72"),
   880 => (x"20",x"3a",x"70",x"6d"),
   881 => (x"20",x"20",x"20",x"20"),
   882 => (x"20",x"20",x"20",x"20"),
   883 => (x"0a",x"64",x"25",x"20"),
   884 => (x"00",x"00",x"00",x"00"),
   885 => (x"20",x"20",x"20",x"20"),
   886 => (x"20",x"20",x"20",x"20"),
   887 => (x"75",x"6f",x"68",x"73"),
   888 => (x"62",x"20",x"64",x"6c"),
   889 => (x"20",x"20",x"3a",x"65"),
   890 => (x"6d",x"69",x"28",x"20"),
   891 => (x"6d",x"65",x"6c",x"70"),
   892 => (x"61",x"74",x"6e",x"65"),
   893 => (x"6e",x"6f",x"69",x"74"),
   894 => (x"70",x"65",x"64",x"2d"),
   895 => (x"65",x"64",x"6e",x"65"),
   896 => (x"0a",x"29",x"74",x"6e"),
   897 => (x"00",x"00",x"00",x"00"),
   898 => (x"69",x"44",x"20",x"20"),
   899 => (x"3a",x"72",x"63",x"73"),
   900 => (x"20",x"20",x"20",x"20"),
   901 => (x"20",x"20",x"20",x"20"),
   902 => (x"20",x"20",x"20",x"20"),
   903 => (x"0a",x"64",x"25",x"20"),
   904 => (x"00",x"00",x"00",x"00"),
   905 => (x"20",x"20",x"20",x"20"),
   906 => (x"20",x"20",x"20",x"20"),
   907 => (x"75",x"6f",x"68",x"73"),
   908 => (x"62",x"20",x"64",x"6c"),
   909 => (x"20",x"20",x"3a",x"65"),
   910 => (x"0a",x"64",x"25",x"20"),
   911 => (x"00",x"00",x"00",x"00"),
   912 => (x"6e",x"45",x"20",x"20"),
   913 => (x"43",x"5f",x"6d",x"75"),
   914 => (x"3a",x"70",x"6d",x"6f"),
   915 => (x"20",x"20",x"20",x"20"),
   916 => (x"20",x"20",x"20",x"20"),
   917 => (x"0a",x"64",x"25",x"20"),
   918 => (x"00",x"00",x"00",x"00"),
   919 => (x"20",x"20",x"20",x"20"),
   920 => (x"20",x"20",x"20",x"20"),
   921 => (x"75",x"6f",x"68",x"73"),
   922 => (x"62",x"20",x"64",x"6c"),
   923 => (x"20",x"20",x"3a",x"65"),
   924 => (x"0a",x"64",x"25",x"20"),
   925 => (x"00",x"00",x"00",x"00"),
   926 => (x"6e",x"49",x"20",x"20"),
   927 => (x"6f",x"43",x"5f",x"74"),
   928 => (x"20",x"3a",x"70",x"6d"),
   929 => (x"20",x"20",x"20",x"20"),
   930 => (x"20",x"20",x"20",x"20"),
   931 => (x"0a",x"64",x"25",x"20"),
   932 => (x"00",x"00",x"00",x"00"),
   933 => (x"20",x"20",x"20",x"20"),
   934 => (x"20",x"20",x"20",x"20"),
   935 => (x"75",x"6f",x"68",x"73"),
   936 => (x"62",x"20",x"64",x"6c"),
   937 => (x"20",x"20",x"3a",x"65"),
   938 => (x"0a",x"64",x"25",x"20"),
   939 => (x"00",x"00",x"00",x"00"),
   940 => (x"74",x"53",x"20",x"20"),
   941 => (x"6f",x"43",x"5f",x"72"),
   942 => (x"20",x"3a",x"70",x"6d"),
   943 => (x"20",x"20",x"20",x"20"),
   944 => (x"20",x"20",x"20",x"20"),
   945 => (x"0a",x"73",x"25",x"20"),
   946 => (x"00",x"00",x"00",x"00"),
   947 => (x"20",x"20",x"20",x"20"),
   948 => (x"20",x"20",x"20",x"20"),
   949 => (x"75",x"6f",x"68",x"73"),
   950 => (x"62",x"20",x"64",x"6c"),
   951 => (x"20",x"20",x"3a",x"65"),
   952 => (x"52",x"48",x"44",x"20"),
   953 => (x"4f",x"54",x"53",x"59"),
   954 => (x"50",x"20",x"45",x"4e"),
   955 => (x"52",x"47",x"4f",x"52"),
   956 => (x"20",x"2c",x"4d",x"41"),
   957 => (x"45",x"4d",x"4f",x"53"),
   958 => (x"52",x"54",x"53",x"20"),
   959 => (x"0a",x"47",x"4e",x"49"),
   960 => (x"00",x"00",x"00",x"00"),
   961 => (x"74",x"78",x"65",x"4e"),
   962 => (x"72",x"74",x"50",x"5f"),
   963 => (x"6f",x"6c",x"47",x"5f"),
   964 => (x"0a",x"3e",x"2d",x"62"),
   965 => (x"00",x"00",x"00",x"00"),
   966 => (x"74",x"50",x"20",x"20"),
   967 => (x"6f",x"43",x"5f",x"72"),
   968 => (x"20",x"3a",x"70",x"6d"),
   969 => (x"20",x"20",x"20",x"20"),
   970 => (x"20",x"20",x"20",x"20"),
   971 => (x"0a",x"64",x"25",x"20"),
   972 => (x"00",x"00",x"00",x"00"),
   973 => (x"20",x"20",x"20",x"20"),
   974 => (x"20",x"20",x"20",x"20"),
   975 => (x"75",x"6f",x"68",x"73"),
   976 => (x"62",x"20",x"64",x"6c"),
   977 => (x"20",x"20",x"3a",x"65"),
   978 => (x"6d",x"69",x"28",x"20"),
   979 => (x"6d",x"65",x"6c",x"70"),
   980 => (x"61",x"74",x"6e",x"65"),
   981 => (x"6e",x"6f",x"69",x"74"),
   982 => (x"70",x"65",x"64",x"2d"),
   983 => (x"65",x"64",x"6e",x"65"),
   984 => (x"2c",x"29",x"74",x"6e"),
   985 => (x"6d",x"61",x"73",x"20"),
   986 => (x"73",x"61",x"20",x"65"),
   987 => (x"6f",x"62",x"61",x"20"),
   988 => (x"00",x"0a",x"65",x"76"),
   989 => (x"69",x"44",x"20",x"20"),
   990 => (x"3a",x"72",x"63",x"73"),
   991 => (x"20",x"20",x"20",x"20"),
   992 => (x"20",x"20",x"20",x"20"),
   993 => (x"20",x"20",x"20",x"20"),
   994 => (x"0a",x"64",x"25",x"20"),
   995 => (x"00",x"00",x"00",x"00"),
   996 => (x"20",x"20",x"20",x"20"),
   997 => (x"20",x"20",x"20",x"20"),
   998 => (x"75",x"6f",x"68",x"73"),
   999 => (x"62",x"20",x"64",x"6c"),
  1000 => (x"20",x"20",x"3a",x"65"),
  1001 => (x"0a",x"64",x"25",x"20"),
  1002 => (x"00",x"00",x"00",x"00"),
  1003 => (x"6e",x"45",x"20",x"20"),
  1004 => (x"43",x"5f",x"6d",x"75"),
  1005 => (x"3a",x"70",x"6d",x"6f"),
  1006 => (x"20",x"20",x"20",x"20"),
  1007 => (x"20",x"20",x"20",x"20"),
  1008 => (x"0a",x"64",x"25",x"20"),
  1009 => (x"00",x"00",x"00",x"00"),
  1010 => (x"20",x"20",x"20",x"20"),
  1011 => (x"20",x"20",x"20",x"20"),
  1012 => (x"75",x"6f",x"68",x"73"),
  1013 => (x"62",x"20",x"64",x"6c"),
  1014 => (x"20",x"20",x"3a",x"65"),
  1015 => (x"0a",x"64",x"25",x"20"),
  1016 => (x"00",x"00",x"00",x"00"),
  1017 => (x"6e",x"49",x"20",x"20"),
  1018 => (x"6f",x"43",x"5f",x"74"),
  1019 => (x"20",x"3a",x"70",x"6d"),
  1020 => (x"20",x"20",x"20",x"20"),
  1021 => (x"20",x"20",x"20",x"20"),
  1022 => (x"0a",x"64",x"25",x"20"),
  1023 => (x"00",x"00",x"00",x"00"),
  1024 => (x"20",x"20",x"20",x"20"),
  1025 => (x"20",x"20",x"20",x"20"),
  1026 => (x"75",x"6f",x"68",x"73"),
  1027 => (x"62",x"20",x"64",x"6c"),
  1028 => (x"20",x"20",x"3a",x"65"),
  1029 => (x"0a",x"64",x"25",x"20"),
  1030 => (x"00",x"00",x"00",x"00"),
  1031 => (x"74",x"53",x"20",x"20"),
  1032 => (x"6f",x"43",x"5f",x"72"),
  1033 => (x"20",x"3a",x"70",x"6d"),
  1034 => (x"20",x"20",x"20",x"20"),
  1035 => (x"20",x"20",x"20",x"20"),
  1036 => (x"0a",x"73",x"25",x"20"),
  1037 => (x"00",x"00",x"00",x"00"),
  1038 => (x"20",x"20",x"20",x"20"),
  1039 => (x"20",x"20",x"20",x"20"),
  1040 => (x"75",x"6f",x"68",x"73"),
  1041 => (x"62",x"20",x"64",x"6c"),
  1042 => (x"20",x"20",x"3a",x"65"),
  1043 => (x"52",x"48",x"44",x"20"),
  1044 => (x"4f",x"54",x"53",x"59"),
  1045 => (x"50",x"20",x"45",x"4e"),
  1046 => (x"52",x"47",x"4f",x"52"),
  1047 => (x"20",x"2c",x"4d",x"41"),
  1048 => (x"45",x"4d",x"4f",x"53"),
  1049 => (x"52",x"54",x"53",x"20"),
  1050 => (x"0a",x"47",x"4e",x"49"),
  1051 => (x"00",x"00",x"00",x"00"),
  1052 => (x"5f",x"74",x"6e",x"49"),
  1053 => (x"6f",x"4c",x"5f",x"31"),
  1054 => (x"20",x"20",x"3a",x"63"),
  1055 => (x"20",x"20",x"20",x"20"),
  1056 => (x"20",x"20",x"20",x"20"),
  1057 => (x"0a",x"64",x"25",x"20"),
  1058 => (x"00",x"00",x"00",x"00"),
  1059 => (x"20",x"20",x"20",x"20"),
  1060 => (x"20",x"20",x"20",x"20"),
  1061 => (x"75",x"6f",x"68",x"73"),
  1062 => (x"62",x"20",x"64",x"6c"),
  1063 => (x"20",x"20",x"3a",x"65"),
  1064 => (x"0a",x"64",x"25",x"20"),
  1065 => (x"00",x"00",x"00",x"00"),
  1066 => (x"5f",x"74",x"6e",x"49"),
  1067 => (x"6f",x"4c",x"5f",x"32"),
  1068 => (x"20",x"20",x"3a",x"63"),
  1069 => (x"20",x"20",x"20",x"20"),
  1070 => (x"20",x"20",x"20",x"20"),
  1071 => (x"0a",x"64",x"25",x"20"),
  1072 => (x"00",x"00",x"00",x"00"),
  1073 => (x"20",x"20",x"20",x"20"),
  1074 => (x"20",x"20",x"20",x"20"),
  1075 => (x"75",x"6f",x"68",x"73"),
  1076 => (x"62",x"20",x"64",x"6c"),
  1077 => (x"20",x"20",x"3a",x"65"),
  1078 => (x"0a",x"64",x"25",x"20"),
  1079 => (x"00",x"00",x"00",x"00"),
  1080 => (x"5f",x"74",x"6e",x"49"),
  1081 => (x"6f",x"4c",x"5f",x"33"),
  1082 => (x"20",x"20",x"3a",x"63"),
  1083 => (x"20",x"20",x"20",x"20"),
  1084 => (x"20",x"20",x"20",x"20"),
  1085 => (x"0a",x"64",x"25",x"20"),
  1086 => (x"00",x"00",x"00",x"00"),
  1087 => (x"20",x"20",x"20",x"20"),
  1088 => (x"20",x"20",x"20",x"20"),
  1089 => (x"75",x"6f",x"68",x"73"),
  1090 => (x"62",x"20",x"64",x"6c"),
  1091 => (x"20",x"20",x"3a",x"65"),
  1092 => (x"0a",x"64",x"25",x"20"),
  1093 => (x"00",x"00",x"00",x"00"),
  1094 => (x"6d",x"75",x"6e",x"45"),
  1095 => (x"63",x"6f",x"4c",x"5f"),
  1096 => (x"20",x"20",x"20",x"3a"),
  1097 => (x"20",x"20",x"20",x"20"),
  1098 => (x"20",x"20",x"20",x"20"),
  1099 => (x"0a",x"64",x"25",x"20"),
  1100 => (x"00",x"00",x"00",x"00"),
  1101 => (x"20",x"20",x"20",x"20"),
  1102 => (x"20",x"20",x"20",x"20"),
  1103 => (x"75",x"6f",x"68",x"73"),
  1104 => (x"62",x"20",x"64",x"6c"),
  1105 => (x"20",x"20",x"3a",x"65"),
  1106 => (x"0a",x"64",x"25",x"20"),
  1107 => (x"00",x"00",x"00",x"00"),
  1108 => (x"5f",x"72",x"74",x"53"),
  1109 => (x"6f",x"4c",x"5f",x"31"),
  1110 => (x"20",x"20",x"3a",x"63"),
  1111 => (x"20",x"20",x"20",x"20"),
  1112 => (x"20",x"20",x"20",x"20"),
  1113 => (x"0a",x"73",x"25",x"20"),
  1114 => (x"00",x"00",x"00",x"00"),
  1115 => (x"20",x"20",x"20",x"20"),
  1116 => (x"20",x"20",x"20",x"20"),
  1117 => (x"75",x"6f",x"68",x"73"),
  1118 => (x"62",x"20",x"64",x"6c"),
  1119 => (x"20",x"20",x"3a",x"65"),
  1120 => (x"52",x"48",x"44",x"20"),
  1121 => (x"4f",x"54",x"53",x"59"),
  1122 => (x"50",x"20",x"45",x"4e"),
  1123 => (x"52",x"47",x"4f",x"52"),
  1124 => (x"20",x"2c",x"4d",x"41"),
  1125 => (x"54",x"53",x"27",x"31"),
  1126 => (x"52",x"54",x"53",x"20"),
  1127 => (x"0a",x"47",x"4e",x"49"),
  1128 => (x"00",x"00",x"00",x"00"),
  1129 => (x"5f",x"72",x"74",x"53"),
  1130 => (x"6f",x"4c",x"5f",x"32"),
  1131 => (x"20",x"20",x"3a",x"63"),
  1132 => (x"20",x"20",x"20",x"20"),
  1133 => (x"20",x"20",x"20",x"20"),
  1134 => (x"0a",x"73",x"25",x"20"),
  1135 => (x"00",x"00",x"00",x"00"),
  1136 => (x"20",x"20",x"20",x"20"),
  1137 => (x"20",x"20",x"20",x"20"),
  1138 => (x"75",x"6f",x"68",x"73"),
  1139 => (x"62",x"20",x"64",x"6c"),
  1140 => (x"20",x"20",x"3a",x"65"),
  1141 => (x"52",x"48",x"44",x"20"),
  1142 => (x"4f",x"54",x"53",x"59"),
  1143 => (x"50",x"20",x"45",x"4e"),
  1144 => (x"52",x"47",x"4f",x"52"),
  1145 => (x"20",x"2c",x"4d",x"41"),
  1146 => (x"44",x"4e",x"27",x"32"),
  1147 => (x"52",x"54",x"53",x"20"),
  1148 => (x"0a",x"47",x"4e",x"49"),
  1149 => (x"00",x"00",x"00",x"00"),
  1150 => (x"00",x"00",x"00",x"0a"),
  1151 => (x"72",x"65",x"73",x"55"),
  1152 => (x"6d",x"69",x"74",x"20"),
  1153 => (x"25",x"20",x"3a",x"65"),
  1154 => (x"1e",x"00",x"0a",x"64"),
  1155 => (x"66",x"c8",x"1e",x"73"),
  1156 => (x"49",x"66",x"cc",x"4b"),
  1157 => (x"ab",x"c2",x"79",x"73"),
  1158 => (x"c1",x"87",x"c4",x"05"),
  1159 => (x"c0",x"87",x"c2",x"4a"),
  1160 => (x"05",x"9a",x"72",x"4a"),
  1161 => (x"79",x"c3",x"87",x"c2"),
  1162 => (x"d8",x"02",x"ab",x"c0"),
  1163 => (x"02",x"ab",x"c1",x"87"),
  1164 => (x"ab",x"c2",x"87",x"d7"),
  1165 => (x"87",x"e5",x"c0",x"02"),
  1166 => (x"c0",x"02",x"ab",x"c3"),
  1167 => (x"ab",x"c4",x"87",x"e5"),
  1168 => (x"de",x"87",x"de",x"02"),
  1169 => (x"da",x"79",x"c0",x"87"),
  1170 => (x"c4",x"cf",x"c1",x"87"),
  1171 => (x"e4",x"c1",x"48",x"bf"),
  1172 => (x"c4",x"06",x"a8",x"b7"),
  1173 => (x"ca",x"79",x"c0",x"87"),
  1174 => (x"c6",x"79",x"c3",x"87"),
  1175 => (x"c2",x"79",x"c1",x"87"),
  1176 => (x"26",x"79",x"c2",x"87"),
  1177 => (x"1e",x"4f",x"26",x"4b"),
  1178 => (x"c2",x"49",x"66",x"c4"),
  1179 => (x"48",x"66",x"c8",x"81"),
  1180 => (x"66",x"cc",x"80",x"71"),
  1181 => (x"26",x"08",x"78",x"08"),
  1182 => (x"1e",x"73",x"1e",x"4f"),
  1183 => (x"1e",x"75",x"1e",x"74"),
  1184 => (x"e4",x"c0",x"86",x"f4"),
  1185 => (x"84",x"c5",x"4c",x"66"),
  1186 => (x"90",x"c4",x"48",x"74"),
  1187 => (x"dc",x"58",x"a6",x"c8"),
  1188 => (x"66",x"c4",x"48",x"66"),
  1189 => (x"58",x"a6",x"c4",x"80"),
  1190 => (x"e8",x"c0",x"48",x"6e"),
  1191 => (x"a6",x"c8",x"78",x"66"),
  1192 => (x"78",x"a4",x"c1",x"48"),
  1193 => (x"dc",x"91",x"c4",x"49"),
  1194 => (x"e8",x"c0",x"81",x"66"),
  1195 => (x"a4",x"de",x"79",x"66"),
  1196 => (x"dc",x"91",x"c4",x"49"),
  1197 => (x"79",x"74",x"81",x"66"),
  1198 => (x"ac",x"b7",x"66",x"c8"),
  1199 => (x"87",x"e0",x"c0",x"01"),
  1200 => (x"c8",x"c3",x"49",x"74"),
  1201 => (x"66",x"e0",x"c0",x"91"),
  1202 => (x"71",x"4d",x"c4",x"81"),
  1203 => (x"82",x"66",x"c4",x"4a"),
  1204 => (x"74",x"4b",x"66",x"c8"),
  1205 => (x"74",x"83",x"c1",x"8b"),
  1206 => (x"c1",x"82",x"75",x"7a"),
  1207 => (x"87",x"f7",x"01",x"8b"),
  1208 => (x"c8",x"c3",x"4a",x"74"),
  1209 => (x"66",x"e0",x"c0",x"92"),
  1210 => (x"c1",x"49",x"74",x"82"),
  1211 => (x"72",x"91",x"c4",x"89"),
  1212 => (x"48",x"69",x"49",x"a1"),
  1213 => (x"79",x"70",x"80",x"c1"),
  1214 => (x"c3",x"49",x"a4",x"d4"),
  1215 => (x"e0",x"c0",x"91",x"c8"),
  1216 => (x"66",x"c4",x"81",x"66"),
  1217 => (x"79",x"bf",x"6e",x"81"),
  1218 => (x"48",x"c4",x"cf",x"c1"),
  1219 => (x"8e",x"f4",x"78",x"c5"),
  1220 => (x"4c",x"26",x"4d",x"26"),
  1221 => (x"4f",x"26",x"4b",x"26"),
  1222 => (x"97",x"1e",x"73",x"1e"),
  1223 => (x"73",x"4b",x"66",x"c8"),
  1224 => (x"66",x"cc",x"97",x"4a"),
  1225 => (x"aa",x"b7",x"71",x"49"),
  1226 => (x"c0",x"87",x"c4",x"02"),
  1227 => (x"c1",x"87",x"c7",x"48"),
  1228 => (x"5b",x"97",x"d0",x"cf"),
  1229 => (x"4b",x"26",x"48",x"c1"),
  1230 => (x"73",x"1e",x"4f",x"26"),
  1231 => (x"75",x"1e",x"74",x"1e"),
  1232 => (x"c2",x"86",x"f8",x"1e"),
  1233 => (x"49",x"66",x"dc",x"4d"),
  1234 => (x"66",x"d8",x"81",x"c1"),
  1235 => (x"a1",x"84",x"c2",x"4c"),
  1236 => (x"49",x"6b",x"97",x"4b"),
  1237 => (x"7e",x"97",x"6c",x"97"),
  1238 => (x"71",x"4a",x"6e",x"97"),
  1239 => (x"c7",x"02",x"aa",x"b7"),
  1240 => (x"48",x"a6",x"c4",x"87"),
  1241 => (x"87",x"cc",x"78",x"c0"),
  1242 => (x"48",x"cc",x"cf",x"c1"),
  1243 => (x"c4",x"50",x"6e",x"97"),
  1244 => (x"78",x"c1",x"48",x"a6"),
  1245 => (x"c4",x"05",x"66",x"c4"),
  1246 => (x"83",x"85",x"c1",x"87"),
  1247 => (x"ad",x"b7",x"c2",x"84"),
  1248 => (x"87",x"cd",x"ff",x"06"),
  1249 => (x"dc",x"4a",x"66",x"d8"),
  1250 => (x"fd",x"fe",x"49",x"66"),
  1251 => (x"b7",x"c0",x"87",x"f0"),
  1252 => (x"87",x"cb",x"06",x"a8"),
  1253 => (x"48",x"c4",x"cf",x"c1"),
  1254 => (x"c1",x"78",x"a5",x"c7"),
  1255 => (x"c0",x"87",x"c2",x"48"),
  1256 => (x"26",x"8e",x"f8",x"48"),
  1257 => (x"26",x"4c",x"26",x"4d"),
  1258 => (x"26",x"4f",x"26",x"4b"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
