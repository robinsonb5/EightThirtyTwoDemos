
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of OSDBoot_832_ROM is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"d4",x"01"),
     1 => (x"18",x"0e",x"87",x"d7"),
     2 => (x"3e",x"27",x"0e",x"1e"),
     3 => (x"0f",x"00",x"00",x"00"),
     4 => (x"80",x"ff",x"48",x"26"),
     5 => (x"27",x"4f",x"08",x"26"),
     6 => (x"00",x"00",x"00",x"23"),
     7 => (x"00",x"30",x"27",x"4f"),
     8 => (x"c2",x"4f",x"00",x"00"),
     9 => (x"27",x"4e",x"c0",x"c0"),
    10 => (x"00",x"00",x"05",x"96"),
    11 => (x"87",x"fd",x"00",x"0f"),
    12 => (x"4e",x"c0",x"f0",x"c1"),
    13 => (x"00",x"00",x"3d",x"27"),
    14 => (x"fd",x"00",x"0f",x"00"),
    15 => (x"0e",x"4f",x"4f",x"87"),
    16 => (x"5c",x"5b",x"5a",x"5e"),
    17 => (x"8e",x"d0",x"0e",x"5d"),
    18 => (x"a6",x"c4",x"4c",x"c0"),
    19 => (x"c0",x"79",x"c0",x"49"),
    20 => (x"c0",x"4b",x"a6",x"e8"),
    21 => (x"c0",x"4a",x"66",x"e4"),
    22 => (x"c1",x"48",x"66",x"e4"),
    23 => (x"a6",x"e8",x"c0",x"80"),
    24 => (x"c1",x"48",x"12",x"58"),
    25 => (x"c0",x"c0",x"c0",x"c0"),
    26 => (x"b7",x"c0",x"c4",x"90"),
    27 => (x"a6",x"c4",x"48",x"90"),
    28 => (x"c5",x"02",x"6e",x"58"),
    29 => (x"66",x"c4",x"87",x"c2"),
    30 => (x"87",x"fe",x"c3",x"02"),
    31 => (x"c0",x"49",x"a6",x"c4"),
    32 => (x"6e",x"4a",x"6e",x"79"),
    33 => (x"a9",x"f0",x"c0",x"49"),
    34 => (x"87",x"c4",x"c3",x"02"),
    35 => (x"02",x"aa",x"e3",x"c1"),
    36 => (x"c1",x"87",x"c5",x"c3"),
    37 => (x"c0",x"02",x"aa",x"e4"),
    38 => (x"ec",x"c1",x"87",x"e3"),
    39 => (x"ef",x"c2",x"02",x"aa"),
    40 => (x"aa",x"f0",x"c1",x"87"),
    41 => (x"87",x"d5",x"c0",x"02"),
    42 => (x"02",x"aa",x"f3",x"c1"),
    43 => (x"c1",x"87",x"c8",x"c2"),
    44 => (x"c0",x"02",x"aa",x"f5"),
    45 => (x"f8",x"c1",x"87",x"c7"),
    46 => (x"f0",x"c2",x"05",x"aa"),
    47 => (x"73",x"83",x"c4",x"87"),
    48 => (x"76",x"8a",x"c4",x"4a"),
    49 => (x"6e",x"79",x"6a",x"49"),
    50 => (x"87",x"db",x"c1",x"02"),
    51 => (x"c0",x"49",x"a6",x"c8"),
    52 => (x"49",x"a6",x"cc",x"79"),
    53 => (x"4a",x"6e",x"79",x"c0"),
    54 => (x"72",x"2a",x"b7",x"dc"),
    55 => (x"6e",x"9d",x"cf",x"4d"),
    56 => (x"c4",x"30",x"c4",x"48"),
    57 => (x"9d",x"75",x"58",x"a6"),
    58 => (x"87",x"c5",x"c0",x"02"),
    59 => (x"c1",x"49",x"a6",x"c8"),
    60 => (x"06",x"ad",x"c9",x"79"),
    61 => (x"c0",x"87",x"c6",x"c0"),
    62 => (x"c3",x"c0",x"85",x"f7"),
    63 => (x"85",x"f0",x"c0",x"87"),
    64 => (x"c0",x"02",x"66",x"c8"),
    65 => (x"1e",x"75",x"87",x"cc"),
    66 => (x"00",x"17",x"74",x"27"),
    67 => (x"86",x"c4",x"0f",x"00"),
    68 => (x"66",x"cc",x"84",x"c1"),
    69 => (x"d0",x"80",x"c1",x"48"),
    70 => (x"66",x"cc",x"58",x"a6"),
    71 => (x"a9",x"b7",x"c8",x"49"),
    72 => (x"87",x"f2",x"fe",x"04"),
    73 => (x"c0",x"87",x"ee",x"c1"),
    74 => (x"74",x"27",x"1e",x"f0"),
    75 => (x"0f",x"00",x"00",x"17"),
    76 => (x"84",x"c1",x"86",x"c4"),
    77 => (x"c4",x"87",x"de",x"c1"),
    78 => (x"c4",x"4a",x"73",x"83"),
    79 => (x"27",x"1e",x"6a",x"8a"),
    80 => (x"00",x"00",x"17",x"a3"),
    81 => (x"70",x"86",x"c4",x"0f"),
    82 => (x"72",x"4c",x"74",x"4a"),
    83 => (x"87",x"c5",x"c1",x"84"),
    84 => (x"c1",x"49",x"a6",x"c4"),
    85 => (x"87",x"fd",x"c0",x"79"),
    86 => (x"4a",x"73",x"83",x"c4"),
    87 => (x"1e",x"6a",x"8a",x"c4"),
    88 => (x"00",x"17",x"74",x"27"),
    89 => (x"86",x"c4",x"0f",x"00"),
    90 => (x"e8",x"c0",x"84",x"c1"),
    91 => (x"27",x"1e",x"6e",x"87"),
    92 => (x"00",x"00",x"17",x"74"),
    93 => (x"c0",x"86",x"c4",x"0f"),
    94 => (x"49",x"6e",x"87",x"db"),
    95 => (x"05",x"a9",x"e5",x"c0"),
    96 => (x"c4",x"87",x"c8",x"c0"),
    97 => (x"79",x"c1",x"49",x"a6"),
    98 => (x"6e",x"87",x"ca",x"c0"),
    99 => (x"17",x"74",x"27",x"1e"),
   100 => (x"c4",x"0f",x"00",x"00"),
   101 => (x"66",x"e4",x"c0",x"86"),
   102 => (x"66",x"e4",x"c0",x"4a"),
   103 => (x"c0",x"80",x"c1",x"48"),
   104 => (x"12",x"58",x"a6",x"e8"),
   105 => (x"c0",x"c0",x"c1",x"48"),
   106 => (x"c4",x"90",x"c0",x"c0"),
   107 => (x"48",x"90",x"b7",x"c0"),
   108 => (x"6e",x"58",x"a6",x"c4"),
   109 => (x"87",x"fe",x"fa",x"05"),
   110 => (x"86",x"d0",x"48",x"74"),
   111 => (x"4c",x"26",x"4d",x"26"),
   112 => (x"4a",x"26",x"4b",x"26"),
   113 => (x"5e",x"0e",x"4f",x"26"),
   114 => (x"cc",x"0e",x"5b",x"5a"),
   115 => (x"2a",x"d8",x"4a",x"66"),
   116 => (x"cc",x"9a",x"ff",x"c3"),
   117 => (x"2b",x"c8",x"4b",x"66"),
   118 => (x"9b",x"c0",x"fc",x"cf"),
   119 => (x"b2",x"73",x"4a",x"72"),
   120 => (x"c8",x"4b",x"66",x"cc"),
   121 => (x"f0",x"ff",x"c0",x"33"),
   122 => (x"72",x"9b",x"c0",x"c0"),
   123 => (x"cc",x"b2",x"73",x"4a"),
   124 => (x"33",x"d8",x"4b",x"66"),
   125 => (x"c0",x"c0",x"fc",x"cf"),
   126 => (x"4a",x"72",x"9b",x"c0"),
   127 => (x"48",x"72",x"b2",x"73"),
   128 => (x"4a",x"26",x"4b",x"26"),
   129 => (x"5e",x"0e",x"4f",x"26"),
   130 => (x"cc",x"0e",x"5b",x"5a"),
   131 => (x"2a",x"c8",x"4a",x"66"),
   132 => (x"cc",x"9a",x"ff",x"c3"),
   133 => (x"33",x"c8",x"4b",x"66"),
   134 => (x"9b",x"c0",x"fc",x"cf"),
   135 => (x"b2",x"73",x"4a",x"72"),
   136 => (x"4b",x"26",x"48",x"72"),
   137 => (x"4f",x"26",x"4a",x"26"),
   138 => (x"5b",x"5a",x"5e",x"0e"),
   139 => (x"4a",x"66",x"cc",x"0e"),
   140 => (x"ff",x"cf",x"2a",x"d0"),
   141 => (x"cc",x"4a",x"9a",x"ff"),
   142 => (x"33",x"d0",x"4b",x"66"),
   143 => (x"9b",x"c0",x"c0",x"f0"),
   144 => (x"b2",x"73",x"4a",x"72"),
   145 => (x"4b",x"26",x"48",x"72"),
   146 => (x"4f",x"26",x"4a",x"26"),
   147 => (x"00",x"00",x"27",x"1e"),
   148 => (x"ff",x"0f",x"10",x"00"),
   149 => (x"4f",x"26",x"87",x"fd"),
   150 => (x"cc",x"1e",x"72",x"1e"),
   151 => (x"df",x"c3",x"4a",x"66"),
   152 => (x"8a",x"f7",x"c0",x"9a"),
   153 => (x"03",x"aa",x"b7",x"c0"),
   154 => (x"c0",x"87",x"c3",x"c0"),
   155 => (x"66",x"c8",x"82",x"e7"),
   156 => (x"cc",x"30",x"c4",x"48"),
   157 => (x"66",x"c8",x"58",x"a6"),
   158 => (x"cc",x"b0",x"72",x"48"),
   159 => (x"66",x"c8",x"58",x"a6"),
   160 => (x"26",x"4a",x"26",x"48"),
   161 => (x"5a",x"5e",x"0e",x"4f"),
   162 => (x"0e",x"5d",x"5c",x"5b"),
   163 => (x"c0",x"e8",x"f6",x"c0"),
   164 => (x"18",x"27",x"4c",x"c0"),
   165 => (x"bf",x"00",x"00",x"1a"),
   166 => (x"27",x"80",x"c1",x"48"),
   167 => (x"00",x"00",x"1a",x"1c"),
   168 => (x"66",x"d4",x"97",x"58"),
   169 => (x"c0",x"c0",x"c1",x"4a"),
   170 => (x"c4",x"92",x"c0",x"c0"),
   171 => (x"4a",x"92",x"b7",x"c0"),
   172 => (x"aa",x"b7",x"d3",x"c1"),
   173 => (x"87",x"e6",x"c0",x"05"),
   174 => (x"00",x"1a",x"18",x"27"),
   175 => (x"79",x"c0",x"49",x"00"),
   176 => (x"00",x"1a",x"1c",x"27"),
   177 => (x"79",x"c0",x"49",x"00"),
   178 => (x"00",x"1a",x"24",x"27"),
   179 => (x"79",x"c0",x"49",x"00"),
   180 => (x"00",x"1a",x"28",x"27"),
   181 => (x"79",x"c0",x"49",x"00"),
   182 => (x"c9",x"7c",x"d3",x"c1"),
   183 => (x"18",x"27",x"87",x"e8"),
   184 => (x"bf",x"00",x"00",x"1a"),
   185 => (x"a9",x"b7",x"c1",x"49"),
   186 => (x"87",x"d5",x"c1",x"05"),
   187 => (x"97",x"7c",x"f4",x"c1"),
   188 => (x"c1",x"4a",x"66",x"d4"),
   189 => (x"c0",x"c0",x"c0",x"c0"),
   190 => (x"b7",x"c0",x"c4",x"92"),
   191 => (x"1e",x"72",x"4a",x"92"),
   192 => (x"00",x"1a",x"28",x"27"),
   193 => (x"27",x"1e",x"bf",x"00"),
   194 => (x"00",x"00",x"02",x"58"),
   195 => (x"27",x"86",x"c8",x"0f"),
   196 => (x"00",x"00",x"1a",x"2c"),
   197 => (x"1a",x"28",x"27",x"58"),
   198 => (x"4d",x"bf",x"00",x"00"),
   199 => (x"06",x"ad",x"b7",x"c3"),
   200 => (x"ca",x"87",x"c6",x"c0"),
   201 => (x"70",x"88",x"75",x"48"),
   202 => (x"c1",x"4a",x"75",x"4d"),
   203 => (x"c1",x"48",x"72",x"82"),
   204 => (x"1a",x"24",x"27",x"30"),
   205 => (x"75",x"58",x"00",x"00"),
   206 => (x"80",x"f0",x"c0",x"48"),
   207 => (x"c5",x"c8",x"7c",x"70"),
   208 => (x"1a",x"28",x"27",x"87"),
   209 => (x"49",x"bf",x"00",x"00"),
   210 => (x"01",x"a9",x"b7",x"c9"),
   211 => (x"27",x"87",x"f7",x"c7"),
   212 => (x"00",x"00",x"1a",x"28"),
   213 => (x"b7",x"c0",x"49",x"bf"),
   214 => (x"e9",x"c7",x"06",x"a9"),
   215 => (x"1a",x"28",x"27",x"87"),
   216 => (x"48",x"bf",x"00",x"00"),
   217 => (x"70",x"80",x"f0",x"c0"),
   218 => (x"1a",x"18",x"27",x"7c"),
   219 => (x"49",x"bf",x"00",x"00"),
   220 => (x"01",x"a9",x"b7",x"c3"),
   221 => (x"97",x"87",x"e9",x"c0"),
   222 => (x"c1",x"4a",x"66",x"d4"),
   223 => (x"c0",x"c0",x"c0",x"c0"),
   224 => (x"b7",x"c0",x"c4",x"92"),
   225 => (x"1e",x"72",x"4a",x"92"),
   226 => (x"00",x"1a",x"24",x"27"),
   227 => (x"27",x"1e",x"bf",x"00"),
   228 => (x"00",x"00",x"02",x"58"),
   229 => (x"27",x"86",x"c8",x"0f"),
   230 => (x"00",x"00",x"1a",x"28"),
   231 => (x"87",x"e6",x"c6",x"58"),
   232 => (x"00",x"1a",x"20",x"27"),
   233 => (x"c3",x"4a",x"bf",x"00"),
   234 => (x"1a",x"18",x"27",x"82"),
   235 => (x"49",x"bf",x"00",x"00"),
   236 => (x"01",x"a9",x"b7",x"72"),
   237 => (x"97",x"87",x"f1",x"c0"),
   238 => (x"c1",x"4a",x"66",x"d4"),
   239 => (x"c0",x"c0",x"c0",x"c0"),
   240 => (x"b7",x"c0",x"c4",x"92"),
   241 => (x"1e",x"72",x"4a",x"92"),
   242 => (x"00",x"1a",x"1c",x"27"),
   243 => (x"27",x"1e",x"bf",x"00"),
   244 => (x"00",x"00",x"02",x"58"),
   245 => (x"27",x"86",x"c8",x"0f"),
   246 => (x"00",x"00",x"1a",x"20"),
   247 => (x"1a",x"2c",x"27",x"58"),
   248 => (x"c1",x"49",x"00",x"00"),
   249 => (x"87",x"de",x"c5",x"79"),
   250 => (x"00",x"1a",x"28",x"27"),
   251 => (x"c0",x"49",x"bf",x"00"),
   252 => (x"c3",x"06",x"a9",x"b7"),
   253 => (x"28",x"27",x"87",x"d0"),
   254 => (x"bf",x"00",x"00",x"1a"),
   255 => (x"a9",x"b7",x"c3",x"49"),
   256 => (x"87",x"c2",x"c3",x"01"),
   257 => (x"00",x"1a",x"24",x"27"),
   258 => (x"c1",x"4a",x"bf",x"00"),
   259 => (x"27",x"82",x"c1",x"32"),
   260 => (x"00",x"00",x"1a",x"18"),
   261 => (x"b7",x"72",x"49",x"bf"),
   262 => (x"c2",x"c2",x"01",x"a9"),
   263 => (x"66",x"d4",x"97",x"87"),
   264 => (x"c0",x"c0",x"c1",x"4a"),
   265 => (x"c4",x"92",x"c0",x"c0"),
   266 => (x"4a",x"92",x"b7",x"c0"),
   267 => (x"30",x"27",x"1e",x"72"),
   268 => (x"bf",x"00",x"00",x"1a"),
   269 => (x"02",x"58",x"27",x"1e"),
   270 => (x"c8",x"0f",x"00",x"00"),
   271 => (x"1a",x"34",x"27",x"86"),
   272 => (x"27",x"58",x"00",x"00"),
   273 => (x"00",x"00",x"1a",x"2c"),
   274 => (x"8a",x"c1",x"4a",x"bf"),
   275 => (x"00",x"1a",x"2c",x"27"),
   276 => (x"79",x"72",x"49",x"00"),
   277 => (x"03",x"aa",x"b7",x"c0"),
   278 => (x"27",x"87",x"eb",x"c3"),
   279 => (x"00",x"00",x"1a",x"1c"),
   280 => (x"30",x"27",x"4a",x"bf"),
   281 => (x"97",x"00",x"00",x"1a"),
   282 => (x"1c",x"27",x"52",x"bf"),
   283 => (x"bf",x"00",x"00",x"1a"),
   284 => (x"27",x"82",x"c1",x"4a"),
   285 => (x"00",x"00",x"1a",x"1c"),
   286 => (x"27",x"79",x"72",x"49"),
   287 => (x"00",x"00",x"1a",x"34"),
   288 => (x"06",x"aa",x"b7",x"bf"),
   289 => (x"27",x"87",x"cd",x"c0"),
   290 => (x"00",x"00",x"1a",x"34"),
   291 => (x"1a",x"1c",x"27",x"49"),
   292 => (x"79",x"bf",x"00",x"00"),
   293 => (x"00",x"1a",x"2c",x"27"),
   294 => (x"79",x"c1",x"49",x"00"),
   295 => (x"27",x"87",x"e7",x"c2"),
   296 => (x"00",x"00",x"1a",x"2c"),
   297 => (x"dd",x"c2",x"05",x"bf"),
   298 => (x"1a",x"30",x"27",x"87"),
   299 => (x"4b",x"bf",x"00",x"00"),
   300 => (x"30",x"27",x"33",x"c4"),
   301 => (x"49",x"00",x"00",x"1a"),
   302 => (x"1c",x"27",x"79",x"73"),
   303 => (x"bf",x"00",x"00",x"1a"),
   304 => (x"c2",x"52",x"73",x"4a"),
   305 => (x"28",x"27",x"87",x"c0"),
   306 => (x"bf",x"00",x"00",x"1a"),
   307 => (x"a9",x"b7",x"c7",x"49"),
   308 => (x"87",x"e6",x"c1",x"04"),
   309 => (x"f4",x"fe",x"4b",x"c0"),
   310 => (x"27",x"79",x"c1",x"49"),
   311 => (x"00",x"00",x"1a",x"1c"),
   312 => (x"27",x"79",x"c0",x"49"),
   313 => (x"00",x"00",x"1a",x"34"),
   314 => (x"b7",x"c0",x"49",x"bf"),
   315 => (x"e5",x"c0",x"06",x"a9"),
   316 => (x"1a",x"1c",x"27",x"87"),
   317 => (x"bf",x"bf",x"00",x"00"),
   318 => (x"1a",x"1c",x"27",x"83"),
   319 => (x"4a",x"bf",x"00",x"00"),
   320 => (x"1c",x"27",x"82",x"c4"),
   321 => (x"49",x"00",x"00",x"1a"),
   322 => (x"34",x"27",x"79",x"72"),
   323 => (x"bf",x"00",x"00",x"1a"),
   324 => (x"ff",x"04",x"aa",x"b7"),
   325 => (x"1e",x"73",x"87",x"db"),
   326 => (x"00",x"1a",x"34",x"27"),
   327 => (x"27",x"1e",x"bf",x"00"),
   328 => (x"00",x"00",x"18",x"62"),
   329 => (x"00",x"3f",x"27",x"1e"),
   330 => (x"cc",x"0f",x"00",x"00"),
   331 => (x"7c",x"c2",x"c1",x"86"),
   332 => (x"00",x"00",x"00",x"27"),
   333 => (x"c0",x"0f",x"bf",x"10"),
   334 => (x"28",x"27",x"87",x"cc"),
   335 => (x"bf",x"00",x"00",x"1a"),
   336 => (x"80",x"f0",x"c0",x"48"),
   337 => (x"4d",x"26",x"7c",x"70"),
   338 => (x"4b",x"26",x"4c",x"26"),
   339 => (x"4f",x"26",x"4a",x"26"),
   340 => (x"5b",x"5a",x"5e",x"0e"),
   341 => (x"d8",x"0e",x"5d",x"5c"),
   342 => (x"4c",x"c0",x"4d",x"66"),
   343 => (x"dc",x"4a",x"66",x"d4"),
   344 => (x"4b",x"72",x"2a",x"b7"),
   345 => (x"66",x"d4",x"9b",x"cf"),
   346 => (x"d8",x"30",x"c4",x"48"),
   347 => (x"b7",x"c9",x"58",x"a6"),
   348 => (x"c6",x"c0",x"06",x"ab"),
   349 => (x"83",x"f7",x"c0",x"87"),
   350 => (x"c0",x"87",x"c3",x"c0"),
   351 => (x"97",x"73",x"83",x"f0"),
   352 => (x"c1",x"85",x"c1",x"7d"),
   353 => (x"ac",x"b7",x"c8",x"84"),
   354 => (x"87",x"d0",x"ff",x"04"),
   355 => (x"4c",x"26",x"4d",x"26"),
   356 => (x"4a",x"26",x"4b",x"26"),
   357 => (x"5e",x"0e",x"4f",x"26"),
   358 => (x"5d",x"5c",x"5b",x"5a"),
   359 => (x"27",x"8e",x"d0",x"0e"),
   360 => (x"00",x"00",x"07",x"99"),
   361 => (x"17",x"a3",x"27",x"1e"),
   362 => (x"c4",x"0f",x"00",x"00"),
   363 => (x"15",x"d7",x"27",x"86"),
   364 => (x"70",x"0f",x"00",x"00"),
   365 => (x"02",x"9a",x"72",x"4a"),
   366 => (x"27",x"87",x"ed",x"c4"),
   367 => (x"00",x"00",x"07",x"82"),
   368 => (x"17",x"a3",x"27",x"1e"),
   369 => (x"c4",x"0f",x"00",x"00"),
   370 => (x"08",x"20",x"27",x"86"),
   371 => (x"70",x"0f",x"00",x"00"),
   372 => (x"02",x"9a",x"72",x"4a"),
   373 => (x"27",x"87",x"c3",x"c4"),
   374 => (x"10",x"00",x"00",x"00"),
   375 => (x"07",x"5a",x"27",x"1e"),
   376 => (x"27",x"1e",x"00",x"00"),
   377 => (x"00",x"00",x"0e",x"df"),
   378 => (x"70",x"86",x"c8",x"0f"),
   379 => (x"02",x"9b",x"73",x"4b"),
   380 => (x"c8",x"87",x"f5",x"c3"),
   381 => (x"79",x"c0",x"49",x"a6"),
   382 => (x"27",x"49",x"a6",x"c4"),
   383 => (x"10",x"00",x"00",x"00"),
   384 => (x"49",x"a6",x"cc",x"79"),
   385 => (x"83",x"c3",x"79",x"c0"),
   386 => (x"00",x"27",x"9b",x"fc"),
   387 => (x"4d",x"10",x"00",x"00"),
   388 => (x"1e",x"75",x"85",x"73"),
   389 => (x"00",x"07",x"4e",x"27"),
   390 => (x"df",x"27",x"1e",x"00"),
   391 => (x"0f",x"00",x"00",x"0e"),
   392 => (x"4a",x"70",x"86",x"c8"),
   393 => (x"c2",x"02",x"9a",x"72"),
   394 => (x"ff",x"c7",x"87",x"e0"),
   395 => (x"c2",x"06",x"ab",x"b7"),
   396 => (x"c0",x"c8",x"87",x"d8"),
   397 => (x"4a",x"66",x"c8",x"1e"),
   398 => (x"72",x"82",x"66",x"d0"),
   399 => (x"17",x"d7",x"27",x"1e"),
   400 => (x"c8",x"0f",x"00",x"00"),
   401 => (x"72",x"4a",x"70",x"86"),
   402 => (x"25",x"49",x"76",x"4c"),
   403 => (x"48",x"66",x"cc",x"79"),
   404 => (x"d0",x"80",x"c0",x"c8"),
   405 => (x"c0",x"c8",x"58",x"a6"),
   406 => (x"ac",x"b7",x"6e",x"8b"),
   407 => (x"87",x"e2",x"c1",x"02"),
   408 => (x"c1",x"48",x"66",x"c8"),
   409 => (x"58",x"a6",x"cc",x"80"),
   410 => (x"00",x"19",x"f8",x"27"),
   411 => (x"66",x"d0",x"1e",x"00"),
   412 => (x"05",x"50",x"27",x"1e"),
   413 => (x"c8",x"0f",x"00",x"00"),
   414 => (x"1a",x"00",x"27",x"86"),
   415 => (x"c0",x"49",x"00",x"00"),
   416 => (x"01",x"27",x"51",x"e0"),
   417 => (x"1e",x"00",x"00",x"1a"),
   418 => (x"50",x"27",x"1e",x"74"),
   419 => (x"0f",x"00",x"00",x"05"),
   420 => (x"09",x"27",x"86",x"c8"),
   421 => (x"49",x"00",x"00",x"1a"),
   422 => (x"27",x"51",x"e0",x"c0"),
   423 => (x"00",x"00",x"1a",x"0a"),
   424 => (x"1e",x"66",x"c4",x"1e"),
   425 => (x"00",x"05",x"50",x"27"),
   426 => (x"86",x"c8",x"0f",x"00"),
   427 => (x"00",x"1a",x"12",x"27"),
   428 => (x"51",x"c0",x"49",x"00"),
   429 => (x"00",x"19",x"f8",x"27"),
   430 => (x"4a",x"27",x"1e",x"00"),
   431 => (x"0f",x"00",x"00",x"10"),
   432 => (x"ff",x"c7",x"86",x"c4"),
   433 => (x"fd",x"01",x"ab",x"b7"),
   434 => (x"66",x"c8",x"87",x"e8"),
   435 => (x"87",x"d8",x"c0",x"05"),
   436 => (x"00",x"00",x"00",x"27"),
   437 => (x"c0",x"0f",x"bf",x"10"),
   438 => (x"66",x"27",x"87",x"ce"),
   439 => (x"1e",x"00",x"00",x"07"),
   440 => (x"00",x"17",x"a3",x"27"),
   441 => (x"86",x"c4",x"0f",x"00"),
   442 => (x"00",x"07",x"af",x"27"),
   443 => (x"a3",x"27",x"1e",x"00"),
   444 => (x"0f",x"00",x"00",x"17"),
   445 => (x"34",x"27",x"86",x"c4"),
   446 => (x"49",x"00",x"00",x"1a"),
   447 => (x"f6",x"c0",x"79",x"c0"),
   448 => (x"4d",x"c0",x"c0",x"e8"),
   449 => (x"27",x"1e",x"ee",x"c0"),
   450 => (x"00",x"00",x"17",x"74"),
   451 => (x"c3",x"86",x"c4",x"0f"),
   452 => (x"4b",x"ff",x"c8",x"f4"),
   453 => (x"4a",x"74",x"4c",x"6d"),
   454 => (x"72",x"9a",x"c0",x"c8"),
   455 => (x"d4",x"c0",x"02",x"9a"),
   456 => (x"c3",x"4a",x"74",x"87"),
   457 => (x"1e",x"72",x"9a",x"ff"),
   458 => (x"00",x"02",x"85",x"27"),
   459 => (x"86",x"c4",x"0f",x"00"),
   460 => (x"c0",x"c9",x"f4",x"c3"),
   461 => (x"c1",x"4a",x"73",x"4b"),
   462 => (x"05",x"9a",x"72",x"8b"),
   463 => (x"ff",x"87",x"d5",x"ff"),
   464 => (x"86",x"d0",x"87",x"c2"),
   465 => (x"4c",x"26",x"4d",x"26"),
   466 => (x"4a",x"26",x"4b",x"26"),
   467 => (x"48",x"43",x"4f",x"26"),
   468 => (x"53",x"4b",x"43",x"45"),
   469 => (x"49",x"42",x"4d",x"55"),
   470 => (x"53",x"4f",x"00",x"4e"),
   471 => (x"32",x"33",x"38",x"44"),
   472 => (x"59",x"53",x"31",x"30"),
   473 => (x"6e",x"55",x"00",x"53"),
   474 => (x"65",x"6c",x"62",x"61"),
   475 => (x"20",x"6f",x"74",x"20"),
   476 => (x"61",x"63",x"6f",x"6c"),
   477 => (x"70",x"20",x"65",x"74"),
   478 => (x"69",x"74",x"72",x"61"),
   479 => (x"6e",x"6f",x"69",x"74"),
   480 => (x"75",x"48",x"00",x"0a"),
   481 => (x"6e",x"69",x"74",x"6e"),
   482 => (x"6f",x"66",x"20",x"67"),
   483 => (x"61",x"70",x"20",x"72"),
   484 => (x"74",x"69",x"74",x"72"),
   485 => (x"0a",x"6e",x"6f",x"69"),
   486 => (x"69",x"6e",x"49",x"00"),
   487 => (x"6c",x"61",x"69",x"74"),
   488 => (x"6e",x"69",x"7a",x"69"),
   489 => (x"44",x"53",x"20",x"67"),
   490 => (x"72",x"61",x"63",x"20"),
   491 => (x"42",x"00",x"0a",x"64"),
   492 => (x"69",x"74",x"6f",x"6f"),
   493 => (x"66",x"20",x"67",x"6e"),
   494 => (x"20",x"6d",x"6f",x"72"),
   495 => (x"33",x"32",x"53",x"52"),
   496 => (x"0e",x"00",x"2e",x"32"),
   497 => (x"5c",x"5b",x"5a",x"5e"),
   498 => (x"66",x"d4",x"0e",x"5d"),
   499 => (x"dc",x"4c",x"c0",x"4d"),
   500 => (x"b7",x"c0",x"49",x"66"),
   501 => (x"fb",x"c0",x"06",x"a9"),
   502 => (x"c1",x"4b",x"15",x"87"),
   503 => (x"c0",x"c0",x"c0",x"c0"),
   504 => (x"b7",x"c0",x"c4",x"93"),
   505 => (x"66",x"d8",x"4b",x"93"),
   506 => (x"c1",x"4a",x"bf",x"97"),
   507 => (x"c0",x"c0",x"c0",x"c0"),
   508 => (x"b7",x"c0",x"c4",x"92"),
   509 => (x"66",x"d8",x"4a",x"92"),
   510 => (x"dc",x"80",x"c1",x"48"),
   511 => (x"b7",x"72",x"58",x"a6"),
   512 => (x"c5",x"c0",x"02",x"ab"),
   513 => (x"c0",x"48",x"c1",x"87"),
   514 => (x"84",x"c1",x"87",x"cc"),
   515 => (x"ac",x"b7",x"66",x"dc"),
   516 => (x"87",x"c5",x"ff",x"04"),
   517 => (x"4d",x"26",x"48",x"c0"),
   518 => (x"4b",x"26",x"4c",x"26"),
   519 => (x"4f",x"26",x"4a",x"26"),
   520 => (x"5b",x"5a",x"5e",x"0e"),
   521 => (x"27",x"0e",x"5d",x"5c"),
   522 => (x"00",x"00",x"1c",x"40"),
   523 => (x"27",x"79",x"c0",x"49"),
   524 => (x"00",x"00",x"19",x"4a"),
   525 => (x"17",x"a3",x"27",x"1e"),
   526 => (x"c4",x"0f",x"00",x"00"),
   527 => (x"1a",x"38",x"27",x"86"),
   528 => (x"c0",x"1e",x"00",x"00"),
   529 => (x"16",x"78",x"27",x"1e"),
   530 => (x"c8",x"0f",x"00",x"00"),
   531 => (x"72",x"4a",x"70",x"86"),
   532 => (x"d3",x"c0",x"05",x"9a"),
   533 => (x"18",x"76",x"27",x"87"),
   534 => (x"27",x"1e",x"00",x"00"),
   535 => (x"00",x"00",x"17",x"a3"),
   536 => (x"c0",x"86",x"c4",x"0f"),
   537 => (x"87",x"d8",x"cf",x"48"),
   538 => (x"00",x"19",x"57",x"27"),
   539 => (x"a3",x"27",x"1e",x"00"),
   540 => (x"0f",x"00",x"00",x"17"),
   541 => (x"4c",x"c0",x"86",x"c4"),
   542 => (x"00",x"1c",x"6c",x"27"),
   543 => (x"79",x"c1",x"49",x"00"),
   544 => (x"6e",x"27",x"1e",x"c8"),
   545 => (x"1e",x"00",x"00",x"19"),
   546 => (x"00",x"1a",x"6e",x"27"),
   547 => (x"c3",x"27",x"1e",x"00"),
   548 => (x"0f",x"00",x"00",x"07"),
   549 => (x"4a",x"70",x"86",x"cc"),
   550 => (x"c0",x"05",x"9a",x"72"),
   551 => (x"6c",x"27",x"87",x"c8"),
   552 => (x"49",x"00",x"00",x"1c"),
   553 => (x"1e",x"c8",x"79",x"c0"),
   554 => (x"00",x"19",x"77",x"27"),
   555 => (x"8a",x"27",x"1e",x"00"),
   556 => (x"1e",x"00",x"00",x"1a"),
   557 => (x"00",x"07",x"c3",x"27"),
   558 => (x"86",x"cc",x"0f",x"00"),
   559 => (x"9a",x"72",x"4a",x"70"),
   560 => (x"87",x"c8",x"c0",x"05"),
   561 => (x"00",x"1c",x"6c",x"27"),
   562 => (x"79",x"c0",x"49",x"00"),
   563 => (x"00",x"1c",x"6c",x"27"),
   564 => (x"27",x"1e",x"bf",x"00"),
   565 => (x"00",x"00",x"19",x"80"),
   566 => (x"00",x"3f",x"27",x"1e"),
   567 => (x"c8",x"0f",x"00",x"00"),
   568 => (x"1c",x"6c",x"27",x"86"),
   569 => (x"02",x"bf",x"00",x"00"),
   570 => (x"27",x"87",x"c0",x"c3"),
   571 => (x"00",x"00",x"1a",x"38"),
   572 => (x"1b",x"f6",x"27",x"4d"),
   573 => (x"27",x"4b",x"00",x"00"),
   574 => (x"00",x"00",x"1c",x"36"),
   575 => (x"72",x"4a",x"bf",x"9f"),
   576 => (x"1c",x"36",x"27",x"1e"),
   577 => (x"27",x"4a",x"00",x"00"),
   578 => (x"00",x"00",x"1a",x"38"),
   579 => (x"d0",x"1e",x"72",x"8a"),
   580 => (x"1e",x"c0",x"c8",x"1e"),
   581 => (x"00",x"18",x"a8",x"27"),
   582 => (x"3f",x"27",x"1e",x"00"),
   583 => (x"0f",x"00",x"00",x"00"),
   584 => (x"4a",x"73",x"86",x"d4"),
   585 => (x"4c",x"6a",x"82",x"c8"),
   586 => (x"00",x"1c",x"36",x"27"),
   587 => (x"4a",x"bf",x"9f",x"00"),
   588 => (x"b7",x"ea",x"d6",x"c5"),
   589 => (x"d3",x"c0",x"05",x"aa"),
   590 => (x"c8",x"4a",x"73",x"87"),
   591 => (x"27",x"1e",x"6a",x"82"),
   592 => (x"00",x"00",x"01",x"c6"),
   593 => (x"70",x"86",x"c4",x"0f"),
   594 => (x"87",x"e4",x"c0",x"4c"),
   595 => (x"fe",x"c7",x"4a",x"75"),
   596 => (x"4a",x"6a",x"9f",x"82"),
   597 => (x"b7",x"d5",x"e9",x"ca"),
   598 => (x"d3",x"c0",x"02",x"aa"),
   599 => (x"18",x"8a",x"27",x"87"),
   600 => (x"27",x"1e",x"00",x"00"),
   601 => (x"00",x"00",x"17",x"a3"),
   602 => (x"c0",x"86",x"c4",x"0f"),
   603 => (x"87",x"d0",x"cb",x"48"),
   604 => (x"e5",x"27",x"1e",x"74"),
   605 => (x"1e",x"00",x"00",x"18"),
   606 => (x"00",x"00",x"3f",x"27"),
   607 => (x"86",x"c8",x"0f",x"00"),
   608 => (x"00",x"1a",x"38",x"27"),
   609 => (x"1e",x"74",x"1e",x"00"),
   610 => (x"00",x"16",x"78",x"27"),
   611 => (x"86",x"c8",x"0f",x"00"),
   612 => (x"9a",x"72",x"4a",x"70"),
   613 => (x"87",x"c5",x"c0",x"05"),
   614 => (x"e3",x"ca",x"48",x"c0"),
   615 => (x"18",x"fd",x"27",x"87"),
   616 => (x"27",x"1e",x"00",x"00"),
   617 => (x"00",x"00",x"17",x"a3"),
   618 => (x"27",x"86",x"c4",x"0f"),
   619 => (x"00",x"00",x"19",x"93"),
   620 => (x"00",x"3f",x"27",x"1e"),
   621 => (x"c4",x"0f",x"00",x"00"),
   622 => (x"27",x"1e",x"c8",x"86"),
   623 => (x"00",x"00",x"19",x"ab"),
   624 => (x"1a",x"8a",x"27",x"1e"),
   625 => (x"27",x"1e",x"00",x"00"),
   626 => (x"00",x"00",x"07",x"c3"),
   627 => (x"70",x"86",x"cc",x"0f"),
   628 => (x"05",x"9a",x"72",x"4a"),
   629 => (x"27",x"87",x"cb",x"c0"),
   630 => (x"00",x"00",x"1c",x"40"),
   631 => (x"c0",x"79",x"c1",x"49"),
   632 => (x"1e",x"c8",x"87",x"f1"),
   633 => (x"00",x"19",x"b4",x"27"),
   634 => (x"6e",x"27",x"1e",x"00"),
   635 => (x"1e",x"00",x"00",x"1a"),
   636 => (x"00",x"07",x"c3",x"27"),
   637 => (x"86",x"cc",x"0f",x"00"),
   638 => (x"9a",x"72",x"4a",x"70"),
   639 => (x"87",x"d3",x"c0",x"02"),
   640 => (x"00",x"19",x"24",x"27"),
   641 => (x"3f",x"27",x"1e",x"00"),
   642 => (x"0f",x"00",x"00",x"00"),
   643 => (x"48",x"c0",x"86",x"c4"),
   644 => (x"27",x"87",x"ed",x"c8"),
   645 => (x"00",x"00",x"1c",x"36"),
   646 => (x"c1",x"4a",x"bf",x"97"),
   647 => (x"05",x"aa",x"b7",x"d5"),
   648 => (x"27",x"87",x"d0",x"c0"),
   649 => (x"00",x"00",x"1c",x"37"),
   650 => (x"c2",x"4a",x"bf",x"97"),
   651 => (x"02",x"aa",x"b7",x"ea"),
   652 => (x"c0",x"87",x"c5",x"c0"),
   653 => (x"87",x"c8",x"c8",x"48"),
   654 => (x"00",x"1a",x"38",x"27"),
   655 => (x"4a",x"bf",x"97",x"00"),
   656 => (x"aa",x"b7",x"e9",x"c3"),
   657 => (x"87",x"d5",x"c0",x"02"),
   658 => (x"00",x"1a",x"38",x"27"),
   659 => (x"4a",x"bf",x"97",x"00"),
   660 => (x"aa",x"b7",x"eb",x"c3"),
   661 => (x"87",x"c5",x"c0",x"02"),
   662 => (x"e3",x"c7",x"48",x"c0"),
   663 => (x"1a",x"43",x"27",x"87"),
   664 => (x"bf",x"97",x"00",x"00"),
   665 => (x"05",x"9a",x"72",x"4a"),
   666 => (x"27",x"87",x"cf",x"c0"),
   667 => (x"00",x"00",x"1a",x"44"),
   668 => (x"c2",x"4a",x"bf",x"97"),
   669 => (x"c0",x"02",x"aa",x"b7"),
   670 => (x"48",x"c0",x"87",x"c5"),
   671 => (x"27",x"87",x"c1",x"c7"),
   672 => (x"00",x"00",x"1a",x"45"),
   673 => (x"27",x"48",x"bf",x"97"),
   674 => (x"00",x"00",x"1c",x"3c"),
   675 => (x"1c",x"38",x"27",x"58"),
   676 => (x"4a",x"bf",x"00",x"00"),
   677 => (x"8b",x"c1",x"4b",x"72"),
   678 => (x"00",x"1c",x"3c",x"27"),
   679 => (x"79",x"73",x"49",x"00"),
   680 => (x"1e",x"72",x"1e",x"73"),
   681 => (x"00",x"19",x"bd",x"27"),
   682 => (x"3f",x"27",x"1e",x"00"),
   683 => (x"0f",x"00",x"00",x"00"),
   684 => (x"46",x"27",x"86",x"cc"),
   685 => (x"97",x"00",x"00",x"1a"),
   686 => (x"82",x"74",x"4a",x"bf"),
   687 => (x"00",x"1a",x"47",x"27"),
   688 => (x"4b",x"bf",x"97",x"00"),
   689 => (x"48",x"73",x"33",x"c8"),
   690 => (x"50",x"27",x"80",x"72"),
   691 => (x"58",x"00",x"00",x"1c"),
   692 => (x"00",x"1a",x"48",x"27"),
   693 => (x"48",x"bf",x"97",x"00"),
   694 => (x"00",x"1c",x"64",x"27"),
   695 => (x"40",x"27",x"58",x"00"),
   696 => (x"bf",x"00",x"00",x"1c"),
   697 => (x"87",x"df",x"c3",x"02"),
   698 => (x"41",x"27",x"1e",x"c8"),
   699 => (x"1e",x"00",x"00",x"19"),
   700 => (x"00",x"1a",x"8a",x"27"),
   701 => (x"c3",x"27",x"1e",x"00"),
   702 => (x"0f",x"00",x"00",x"07"),
   703 => (x"4a",x"70",x"86",x"cc"),
   704 => (x"c0",x"02",x"9a",x"72"),
   705 => (x"48",x"c0",x"87",x"c5"),
   706 => (x"27",x"87",x"f5",x"c4"),
   707 => (x"00",x"00",x"1c",x"38"),
   708 => (x"48",x"73",x"4b",x"bf"),
   709 => (x"68",x"27",x"30",x"c4"),
   710 => (x"58",x"00",x"00",x"1c"),
   711 => (x"00",x"1c",x"5c",x"27"),
   712 => (x"79",x"73",x"49",x"00"),
   713 => (x"00",x"1a",x"5d",x"27"),
   714 => (x"4a",x"bf",x"97",x"00"),
   715 => (x"5c",x"27",x"32",x"c8"),
   716 => (x"97",x"00",x"00",x"1a"),
   717 => (x"4a",x"72",x"4c",x"bf"),
   718 => (x"5e",x"27",x"82",x"74"),
   719 => (x"97",x"00",x"00",x"1a"),
   720 => (x"34",x"d0",x"4c",x"bf"),
   721 => (x"82",x"74",x"4a",x"72"),
   722 => (x"00",x"1a",x"5f",x"27"),
   723 => (x"4c",x"bf",x"97",x"00"),
   724 => (x"4a",x"72",x"34",x"d8"),
   725 => (x"68",x"27",x"82",x"74"),
   726 => (x"49",x"00",x"00",x"1c"),
   727 => (x"4a",x"72",x"79",x"72"),
   728 => (x"00",x"1c",x"60",x"27"),
   729 => (x"72",x"92",x"bf",x"00"),
   730 => (x"1c",x"4c",x"27",x"4a"),
   731 => (x"82",x"bf",x"00",x"00"),
   732 => (x"00",x"1c",x"50",x"27"),
   733 => (x"79",x"72",x"49",x"00"),
   734 => (x"00",x"1a",x"65",x"27"),
   735 => (x"4c",x"bf",x"97",x"00"),
   736 => (x"64",x"27",x"34",x"c8"),
   737 => (x"97",x"00",x"00",x"1a"),
   738 => (x"4c",x"74",x"4d",x"bf"),
   739 => (x"66",x"27",x"84",x"75"),
   740 => (x"97",x"00",x"00",x"1a"),
   741 => (x"35",x"d0",x"4d",x"bf"),
   742 => (x"84",x"75",x"4c",x"74"),
   743 => (x"00",x"1a",x"67",x"27"),
   744 => (x"4d",x"bf",x"97",x"00"),
   745 => (x"35",x"d8",x"9d",x"cf"),
   746 => (x"84",x"75",x"4c",x"74"),
   747 => (x"00",x"1c",x"54",x"27"),
   748 => (x"79",x"74",x"49",x"00"),
   749 => (x"4b",x"73",x"8c",x"c2"),
   750 => (x"48",x"73",x"93",x"74"),
   751 => (x"5c",x"27",x"80",x"72"),
   752 => (x"58",x"00",x"00",x"1c"),
   753 => (x"27",x"87",x"f7",x"c1"),
   754 => (x"00",x"00",x"1a",x"4a"),
   755 => (x"c8",x"4a",x"bf",x"97"),
   756 => (x"1a",x"49",x"27",x"32"),
   757 => (x"bf",x"97",x"00",x"00"),
   758 => (x"73",x"4a",x"72",x"4b"),
   759 => (x"1c",x"64",x"27",x"82"),
   760 => (x"72",x"49",x"00",x"00"),
   761 => (x"c7",x"32",x"c5",x"79"),
   762 => (x"2a",x"c9",x"82",x"ff"),
   763 => (x"00",x"1c",x"5c",x"27"),
   764 => (x"79",x"72",x"49",x"00"),
   765 => (x"00",x"1a",x"4f",x"27"),
   766 => (x"4b",x"bf",x"97",x"00"),
   767 => (x"4e",x"27",x"33",x"c8"),
   768 => (x"97",x"00",x"00",x"1a"),
   769 => (x"4b",x"73",x"4c",x"bf"),
   770 => (x"68",x"27",x"83",x"74"),
   771 => (x"49",x"00",x"00",x"1c"),
   772 => (x"4b",x"73",x"79",x"73"),
   773 => (x"00",x"1c",x"60",x"27"),
   774 => (x"73",x"93",x"bf",x"00"),
   775 => (x"1c",x"4c",x"27",x"4b"),
   776 => (x"83",x"bf",x"00",x"00"),
   777 => (x"00",x"1c",x"58",x"27"),
   778 => (x"79",x"73",x"49",x"00"),
   779 => (x"00",x"1c",x"54",x"27"),
   780 => (x"79",x"c0",x"49",x"00"),
   781 => (x"80",x"72",x"48",x"73"),
   782 => (x"00",x"1c",x"54",x"27"),
   783 => (x"48",x"c1",x"58",x"00"),
   784 => (x"4c",x"26",x"4d",x"26"),
   785 => (x"4a",x"26",x"4b",x"26"),
   786 => (x"5e",x"0e",x"4f",x"26"),
   787 => (x"5d",x"5c",x"5b",x"5a"),
   788 => (x"1c",x"40",x"27",x"0e"),
   789 => (x"02",x"bf",x"00",x"00"),
   790 => (x"d4",x"87",x"cf",x"c0"),
   791 => (x"b7",x"c7",x"4c",x"66"),
   792 => (x"4b",x"66",x"d4",x"2c"),
   793 => (x"c0",x"9b",x"ff",x"c1"),
   794 => (x"66",x"d4",x"87",x"cc"),
   795 => (x"2c",x"b7",x"c8",x"4c"),
   796 => (x"c3",x"4b",x"66",x"d4"),
   797 => (x"38",x"27",x"9b",x"ff"),
   798 => (x"1e",x"00",x"00",x"1a"),
   799 => (x"00",x"1c",x"4c",x"27"),
   800 => (x"74",x"4a",x"bf",x"00"),
   801 => (x"27",x"1e",x"72",x"82"),
   802 => (x"00",x"00",x"16",x"78"),
   803 => (x"70",x"86",x"c8",x"0f"),
   804 => (x"05",x"9a",x"72",x"4a"),
   805 => (x"c0",x"87",x"c5",x"c0"),
   806 => (x"87",x"f2",x"c0",x"48"),
   807 => (x"00",x"1c",x"40",x"27"),
   808 => (x"c0",x"02",x"bf",x"00"),
   809 => (x"4a",x"73",x"87",x"d7"),
   810 => (x"4a",x"72",x"92",x"c4"),
   811 => (x"00",x"1a",x"38",x"27"),
   812 => (x"4d",x"6a",x"82",x"00"),
   813 => (x"ff",x"ff",x"ff",x"cf"),
   814 => (x"cf",x"c0",x"9d",x"ff"),
   815 => (x"c2",x"4a",x"73",x"87"),
   816 => (x"27",x"4a",x"72",x"92"),
   817 => (x"00",x"00",x"1a",x"38"),
   818 => (x"4d",x"6a",x"9f",x"82"),
   819 => (x"4d",x"26",x"48",x"75"),
   820 => (x"4b",x"26",x"4c",x"26"),
   821 => (x"4f",x"26",x"4a",x"26"),
   822 => (x"5b",x"5a",x"5e",x"0e"),
   823 => (x"cc",x"0e",x"5d",x"5c"),
   824 => (x"ff",x"ff",x"cf",x"8e"),
   825 => (x"c0",x"4d",x"f8",x"ff"),
   826 => (x"27",x"49",x"76",x"4c"),
   827 => (x"00",x"00",x"1c",x"54"),
   828 => (x"a6",x"c4",x"79",x"bf"),
   829 => (x"1c",x"58",x"27",x"49"),
   830 => (x"79",x"bf",x"00",x"00"),
   831 => (x"00",x"1c",x"40",x"27"),
   832 => (x"c0",x"02",x"bf",x"00"),
   833 => (x"38",x"27",x"87",x"cc"),
   834 => (x"bf",x"00",x"00",x"1c"),
   835 => (x"c0",x"32",x"c4",x"4a"),
   836 => (x"5c",x"27",x"87",x"c9"),
   837 => (x"bf",x"00",x"00",x"1c"),
   838 => (x"c8",x"32",x"c4",x"4a"),
   839 => (x"79",x"72",x"49",x"a6"),
   840 => (x"66",x"c8",x"4b",x"c0"),
   841 => (x"06",x"a9",x"c0",x"49"),
   842 => (x"73",x"87",x"d0",x"c3"),
   843 => (x"72",x"9a",x"cf",x"4a"),
   844 => (x"e4",x"c0",x"05",x"9a"),
   845 => (x"1a",x"38",x"27",x"87"),
   846 => (x"c8",x"1e",x"00",x"00"),
   847 => (x"66",x"c8",x"4a",x"66"),
   848 => (x"cc",x"80",x"c1",x"48"),
   849 => (x"1e",x"72",x"58",x"a6"),
   850 => (x"00",x"16",x"78",x"27"),
   851 => (x"86",x"c8",x"0f",x"00"),
   852 => (x"00",x"1a",x"38",x"27"),
   853 => (x"c3",x"c0",x"4c",x"00"),
   854 => (x"84",x"e0",x"c0",x"87"),
   855 => (x"72",x"4a",x"6c",x"97"),
   856 => (x"cd",x"c2",x"02",x"9a"),
   857 => (x"4a",x"6c",x"97",x"87"),
   858 => (x"aa",x"b7",x"e5",x"c3"),
   859 => (x"87",x"c2",x"c2",x"02"),
   860 => (x"82",x"cb",x"4a",x"74"),
   861 => (x"d8",x"4a",x"6a",x"97"),
   862 => (x"05",x"9a",x"72",x"9a"),
   863 => (x"74",x"87",x"f3",x"c1"),
   864 => (x"17",x"a3",x"27",x"1e"),
   865 => (x"c4",x"0f",x"00",x"00"),
   866 => (x"c0",x"1e",x"cb",x"86"),
   867 => (x"74",x"1e",x"66",x"e8"),
   868 => (x"07",x"c3",x"27",x"1e"),
   869 => (x"cc",x"0f",x"00",x"00"),
   870 => (x"72",x"4a",x"70",x"86"),
   871 => (x"d1",x"c1",x"05",x"9a"),
   872 => (x"dc",x"4b",x"74",x"87"),
   873 => (x"66",x"e0",x"c0",x"83"),
   874 => (x"6b",x"82",x"c4",x"4a"),
   875 => (x"da",x"4b",x"74",x"7a"),
   876 => (x"66",x"e0",x"c0",x"83"),
   877 => (x"9f",x"82",x"c8",x"4a"),
   878 => (x"7a",x"70",x"48",x"6b"),
   879 => (x"40",x"27",x"4d",x"72"),
   880 => (x"bf",x"00",x"00",x"1c"),
   881 => (x"87",x"d5",x"c0",x"02"),
   882 => (x"82",x"d4",x"4a",x"74"),
   883 => (x"c0",x"4a",x"6a",x"9f"),
   884 => (x"72",x"9a",x"ff",x"ff"),
   885 => (x"c4",x"30",x"d0",x"48"),
   886 => (x"c4",x"c0",x"58",x"a6"),
   887 => (x"c0",x"49",x"76",x"87"),
   888 => (x"6d",x"48",x"6e",x"79"),
   889 => (x"c0",x"7d",x"70",x"80"),
   890 => (x"c0",x"49",x"66",x"e0"),
   891 => (x"c1",x"48",x"c1",x"79"),
   892 => (x"83",x"c1",x"87",x"ce"),
   893 => (x"04",x"ab",x"66",x"c8"),
   894 => (x"cf",x"87",x"f0",x"fc"),
   895 => (x"f8",x"ff",x"ff",x"ff"),
   896 => (x"1c",x"40",x"27",x"4d"),
   897 => (x"02",x"bf",x"00",x"00"),
   898 => (x"6e",x"87",x"f3",x"c0"),
   899 => (x"0c",x"4a",x"27",x"1e"),
   900 => (x"c4",x"0f",x"00",x"00"),
   901 => (x"58",x"a6",x"c4",x"86"),
   902 => (x"9a",x"75",x"4a",x"6e"),
   903 => (x"c0",x"02",x"aa",x"75"),
   904 => (x"4a",x"6e",x"87",x"dc"),
   905 => (x"4a",x"72",x"8a",x"c2"),
   906 => (x"00",x"1c",x"38",x"27"),
   907 => (x"27",x"92",x"bf",x"00"),
   908 => (x"00",x"00",x"1c",x"50"),
   909 => (x"80",x"72",x"48",x"bf"),
   910 => (x"fb",x"58",x"a6",x"c8"),
   911 => (x"48",x"c0",x"87",x"e2"),
   912 => (x"ff",x"ff",x"ff",x"cf"),
   913 => (x"86",x"cc",x"4d",x"f8"),
   914 => (x"4c",x"26",x"4d",x"26"),
   915 => (x"4a",x"26",x"4b",x"26"),
   916 => (x"5e",x"0e",x"4f",x"26"),
   917 => (x"cc",x"0e",x"5b",x"5a"),
   918 => (x"c1",x"4a",x"bf",x"66"),
   919 => (x"49",x"66",x"cc",x"82"),
   920 => (x"4a",x"72",x"79",x"72"),
   921 => (x"00",x"1c",x"3c",x"27"),
   922 => (x"72",x"9a",x"bf",x"00"),
   923 => (x"d3",x"c0",x"05",x"9a"),
   924 => (x"4a",x"66",x"cc",x"87"),
   925 => (x"1e",x"6a",x"82",x"c8"),
   926 => (x"00",x"0c",x"4a",x"27"),
   927 => (x"86",x"c4",x"0f",x"00"),
   928 => (x"7a",x"73",x"4b",x"70"),
   929 => (x"4b",x"26",x"48",x"c1"),
   930 => (x"4f",x"26",x"4a",x"26"),
   931 => (x"5b",x"5a",x"5e",x"0e"),
   932 => (x"1c",x"50",x"27",x"0e"),
   933 => (x"4a",x"bf",x"00",x"00"),
   934 => (x"c8",x"4b",x"66",x"cc"),
   935 => (x"c2",x"4b",x"6b",x"83"),
   936 => (x"27",x"4b",x"73",x"8b"),
   937 => (x"00",x"00",x"1c",x"38"),
   938 => (x"4a",x"72",x"93",x"bf"),
   939 => (x"3c",x"27",x"82",x"73"),
   940 => (x"bf",x"00",x"00",x"1c"),
   941 => (x"bf",x"66",x"cc",x"4b"),
   942 => (x"73",x"4a",x"72",x"9b"),
   943 => (x"1e",x"66",x"d0",x"82"),
   944 => (x"78",x"27",x"1e",x"72"),
   945 => (x"0f",x"00",x"00",x"16"),
   946 => (x"4a",x"70",x"86",x"c8"),
   947 => (x"c0",x"05",x"9a",x"72"),
   948 => (x"48",x"c0",x"87",x"c5"),
   949 => (x"c1",x"87",x"c2",x"c0"),
   950 => (x"26",x"4b",x"26",x"48"),
   951 => (x"0e",x"4f",x"26",x"4a"),
   952 => (x"5c",x"5b",x"5a",x"5e"),
   953 => (x"66",x"d8",x"0e",x"5d"),
   954 => (x"1e",x"66",x"d4",x"4c"),
   955 => (x"00",x"1c",x"70",x"27"),
   956 => (x"d8",x"27",x"1e",x"00"),
   957 => (x"0f",x"00",x"00",x"0c"),
   958 => (x"4a",x"70",x"86",x"c8"),
   959 => (x"c1",x"02",x"9a",x"72"),
   960 => (x"74",x"27",x"87",x"df"),
   961 => (x"bf",x"00",x"00",x"1c"),
   962 => (x"82",x"ff",x"c7",x"4a"),
   963 => (x"4d",x"72",x"2a",x"c9"),
   964 => (x"83",x"27",x"4b",x"c0"),
   965 => (x"1e",x"00",x"00",x"0f"),
   966 => (x"00",x"17",x"a3",x"27"),
   967 => (x"86",x"c4",x"0f",x"00"),
   968 => (x"06",x"ad",x"b7",x"c0"),
   969 => (x"74",x"87",x"d0",x"c1"),
   970 => (x"1c",x"70",x"27",x"1e"),
   971 => (x"27",x"1e",x"00",x"00"),
   972 => (x"00",x"00",x"0e",x"8c"),
   973 => (x"70",x"86",x"c8",x"0f"),
   974 => (x"05",x"9a",x"72",x"4a"),
   975 => (x"c0",x"87",x"c5",x"c0"),
   976 => (x"87",x"f5",x"c0",x"48"),
   977 => (x"00",x"1c",x"70",x"27"),
   978 => (x"52",x"27",x"1e",x"00"),
   979 => (x"0f",x"00",x"00",x"0e"),
   980 => (x"c0",x"c8",x"86",x"c4"),
   981 => (x"75",x"83",x"c1",x"84"),
   982 => (x"ff",x"04",x"ab",x"b7"),
   983 => (x"d6",x"c0",x"87",x"c9"),
   984 => (x"1e",x"66",x"d4",x"87"),
   985 => (x"00",x"0f",x"9c",x"27"),
   986 => (x"3f",x"27",x"1e",x"00"),
   987 => (x"0f",x"00",x"00",x"00"),
   988 => (x"48",x"c0",x"86",x"c8"),
   989 => (x"c1",x"87",x"c2",x"c0"),
   990 => (x"26",x"4d",x"26",x"48"),
   991 => (x"26",x"4b",x"26",x"4c"),
   992 => (x"4f",x"4f",x"26",x"4a"),
   993 => (x"65",x"6e",x"65",x"70"),
   994 => (x"69",x"66",x"20",x"64"),
   995 => (x"20",x"2c",x"65",x"6c"),
   996 => (x"64",x"61",x"6f",x"6c"),
   997 => (x"2e",x"67",x"6e",x"69"),
   998 => (x"00",x"0a",x"2e",x"2e"),
   999 => (x"27",x"6e",x"61",x"43"),
  1000 => (x"70",x"6f",x"20",x"74"),
  1001 => (x"25",x"20",x"6e",x"65"),
  1002 => (x"1e",x"00",x"0a",x"73"),
  1003 => (x"66",x"c8",x"1e",x"72"),
  1004 => (x"87",x"d1",x"c0",x"02"),
  1005 => (x"00",x"1c",x"7c",x"27"),
  1006 => (x"66",x"c8",x"49",x"00"),
  1007 => (x"1c",x"84",x"27",x"79"),
  1008 => (x"c0",x"49",x"00",x"00"),
  1009 => (x"1c",x"84",x"27",x"79"),
  1010 => (x"05",x"bf",x"00",x"00"),
  1011 => (x"27",x"87",x"dc",x"c0"),
  1012 => (x"00",x"00",x"1c",x"7c"),
  1013 => (x"48",x"72",x"4a",x"bf"),
  1014 => (x"80",x"27",x"80",x"c4"),
  1015 => (x"58",x"00",x"00",x"1c"),
  1016 => (x"00",x"1c",x"80",x"27"),
  1017 => (x"79",x"6a",x"49",x"00"),
  1018 => (x"27",x"87",x"cf",x"c0"),
  1019 => (x"00",x"00",x"1c",x"80"),
  1020 => (x"30",x"c8",x"48",x"bf"),
  1021 => (x"00",x"1c",x"84",x"27"),
  1022 => (x"84",x"27",x"58",x"00"),
  1023 => (x"bf",x"00",x"00",x"1c"),
  1024 => (x"72",x"82",x"c1",x"4a"),
  1025 => (x"27",x"98",x"c3",x"48"),
  1026 => (x"00",x"00",x"1c",x"88"),
  1027 => (x"1c",x"80",x"27",x"58"),
  1028 => (x"4a",x"bf",x"00",x"00"),
  1029 => (x"72",x"2a",x"b7",x"d8"),
  1030 => (x"26",x"4a",x"26",x"48"),
  1031 => (x"5a",x"5e",x"0e",x"4f"),
  1032 => (x"66",x"cc",x"0e",x"5b"),
  1033 => (x"87",x"c3",x"fe",x"1e"),
  1034 => (x"4b",x"70",x"86",x"c4"),
  1035 => (x"9b",x"73",x"4a",x"c0"),
  1036 => (x"87",x"ce",x"c0",x"02"),
  1037 => (x"1e",x"c0",x"82",x"c1"),
  1038 => (x"c4",x"87",x"f0",x"fd"),
  1039 => (x"ff",x"4b",x"70",x"86"),
  1040 => (x"48",x"72",x"87",x"ec"),
  1041 => (x"4a",x"26",x"4b",x"26"),
  1042 => (x"5e",x"0e",x"4f",x"26"),
  1043 => (x"5d",x"5c",x"5b",x"5a"),
  1044 => (x"c0",x"8e",x"c8",x"0e"),
  1045 => (x"c4",x"c0",x"e4",x"f6"),
  1046 => (x"e4",x"f6",x"c0",x"4c"),
  1047 => (x"dc",x"4b",x"c0",x"c0"),
  1048 => (x"f8",x"fe",x"1e",x"66"),
  1049 => (x"70",x"86",x"c4",x"87"),
  1050 => (x"c2",x"4d",x"72",x"4a"),
  1051 => (x"c1",x"49",x"76",x"85"),
  1052 => (x"7c",x"9f",x"d0",x"79"),
  1053 => (x"9f",x"c1",x"c0",x"c1"),
  1054 => (x"4a",x"6b",x"9f",x"7b"),
  1055 => (x"c0",x"7b",x"9f",x"c0"),
  1056 => (x"6b",x"9f",x"7b",x"9f"),
  1057 => (x"58",x"a6",x"c8",x"48"),
  1058 => (x"72",x"9a",x"c0",x"c4"),
  1059 => (x"fd",x"c1",x"02",x"9a"),
  1060 => (x"c0",x"02",x"6e",x"87"),
  1061 => (x"66",x"c4",x"87",x"e6"),
  1062 => (x"c6",x"c0",x"c8",x"49"),
  1063 => (x"ed",x"c1",x"05",x"a9"),
  1064 => (x"c0",x"49",x"76",x"87"),
  1065 => (x"ca",x"eb",x"fa",x"79"),
  1066 => (x"9f",x"c1",x"7b",x"9f"),
  1067 => (x"7b",x"9f",x"c0",x"7b"),
  1068 => (x"c0",x"7b",x"9f",x"75"),
  1069 => (x"9f",x"c0",x"7b",x"9f"),
  1070 => (x"87",x"d2",x"c1",x"7b"),
  1071 => (x"2a",x"c1",x"4a",x"75"),
  1072 => (x"b2",x"c0",x"c0",x"c8"),
  1073 => (x"72",x"49",x"66",x"c4"),
  1074 => (x"c1",x"c1",x"05",x"a9"),
  1075 => (x"1e",x"66",x"dc",x"87"),
  1076 => (x"c4",x"87",x"d8",x"fb"),
  1077 => (x"58",x"a6",x"c4",x"86"),
  1078 => (x"8d",x"c1",x"4a",x"75"),
  1079 => (x"c0",x"02",x"9a",x"72"),
  1080 => (x"4c",x"6e",x"87",x"de"),
  1081 => (x"74",x"7b",x"97",x"74"),
  1082 => (x"c9",x"c0",x"02",x"9c"),
  1083 => (x"fa",x"1e",x"c0",x"87"),
  1084 => (x"86",x"c4",x"87",x"f9"),
  1085 => (x"4a",x"75",x"4c",x"70"),
  1086 => (x"9a",x"72",x"8d",x"c1"),
  1087 => (x"87",x"e4",x"ff",x"05"),
  1088 => (x"c0",x"e4",x"f6",x"c0"),
  1089 => (x"9f",x"d1",x"4c",x"c4"),
  1090 => (x"c0",x"48",x"c1",x"7c"),
  1091 => (x"9f",x"d1",x"87",x"c6"),
  1092 => (x"87",x"dd",x"fd",x"7c"),
  1093 => (x"4d",x"26",x"86",x"c8"),
  1094 => (x"4b",x"26",x"4c",x"26"),
  1095 => (x"4f",x"26",x"4a",x"26"),
  1096 => (x"5b",x"5a",x"5e",x"0e"),
  1097 => (x"e4",x"c0",x"0e",x"5c"),
  1098 => (x"4c",x"ff",x"c3",x"8e"),
  1099 => (x"c0",x"e4",x"f6",x"c0"),
  1100 => (x"7b",x"74",x"4b",x"c0"),
  1101 => (x"9a",x"74",x"4a",x"6b"),
  1102 => (x"48",x"6b",x"7b",x"74"),
  1103 => (x"a6",x"c4",x"98",x"74"),
  1104 => (x"c8",x"48",x"6e",x"58"),
  1105 => (x"58",x"a6",x"c8",x"30"),
  1106 => (x"72",x"49",x"a6",x"c8"),
  1107 => (x"c4",x"4a",x"72",x"79"),
  1108 => (x"7b",x"74",x"b2",x"66"),
  1109 => (x"98",x"74",x"48",x"6b"),
  1110 => (x"cc",x"58",x"a6",x"d0"),
  1111 => (x"30",x"d0",x"48",x"66"),
  1112 => (x"d4",x"58",x"a6",x"d4"),
  1113 => (x"79",x"72",x"49",x"a6"),
  1114 => (x"66",x"d0",x"4a",x"72"),
  1115 => (x"6b",x"7b",x"74",x"b2"),
  1116 => (x"dc",x"98",x"74",x"48"),
  1117 => (x"66",x"d8",x"58",x"a6"),
  1118 => (x"c0",x"30",x"d8",x"48"),
  1119 => (x"c0",x"58",x"a6",x"e0"),
  1120 => (x"72",x"49",x"a6",x"e0"),
  1121 => (x"dc",x"4a",x"72",x"79"),
  1122 => (x"48",x"72",x"b2",x"66"),
  1123 => (x"26",x"86",x"e4",x"c0"),
  1124 => (x"26",x"4b",x"26",x"4c"),
  1125 => (x"0e",x"4f",x"26",x"4a"),
  1126 => (x"5c",x"5b",x"5a",x"5e"),
  1127 => (x"c3",x"8e",x"d8",x"0e"),
  1128 => (x"f6",x"c0",x"4c",x"ff"),
  1129 => (x"4b",x"c0",x"c0",x"e4"),
  1130 => (x"4a",x"6b",x"7b",x"74"),
  1131 => (x"7b",x"74",x"9a",x"74"),
  1132 => (x"48",x"6b",x"32",x"c8"),
  1133 => (x"a6",x"c4",x"98",x"74"),
  1134 => (x"49",x"a6",x"c4",x"58"),
  1135 => (x"4a",x"72",x"79",x"72"),
  1136 => (x"7b",x"74",x"b2",x"6e"),
  1137 => (x"48",x"6b",x"32",x"c8"),
  1138 => (x"a6",x"cc",x"98",x"74"),
  1139 => (x"49",x"a6",x"cc",x"58"),
  1140 => (x"4a",x"72",x"79",x"72"),
  1141 => (x"74",x"b2",x"66",x"c8"),
  1142 => (x"6b",x"32",x"c8",x"7b"),
  1143 => (x"d4",x"98",x"74",x"48"),
  1144 => (x"a6",x"d4",x"58",x"a6"),
  1145 => (x"72",x"79",x"72",x"49"),
  1146 => (x"b2",x"66",x"d0",x"4a"),
  1147 => (x"86",x"d8",x"48",x"72"),
  1148 => (x"4b",x"26",x"4c",x"26"),
  1149 => (x"4f",x"26",x"4a",x"26"),
  1150 => (x"5b",x"5a",x"5e",x"0e"),
  1151 => (x"c0",x"0e",x"5d",x"5c"),
  1152 => (x"c0",x"c0",x"e4",x"f6"),
  1153 => (x"48",x"66",x"d4",x"4b"),
  1154 => (x"70",x"98",x"ff",x"c3"),
  1155 => (x"1c",x"88",x"27",x"7b"),
  1156 => (x"05",x"bf",x"00",x"00"),
  1157 => (x"d8",x"87",x"c8",x"c0"),
  1158 => (x"30",x"c9",x"48",x"66"),
  1159 => (x"d8",x"58",x"a6",x"dc"),
  1160 => (x"2a",x"d8",x"4a",x"66"),
  1161 => (x"ff",x"c3",x"48",x"72"),
  1162 => (x"d8",x"7b",x"70",x"98"),
  1163 => (x"2a",x"d0",x"4a",x"66"),
  1164 => (x"ff",x"c3",x"48",x"72"),
  1165 => (x"d8",x"7b",x"70",x"98"),
  1166 => (x"2a",x"c8",x"4a",x"66"),
  1167 => (x"ff",x"c3",x"48",x"72"),
  1168 => (x"d8",x"7b",x"70",x"98"),
  1169 => (x"ff",x"c3",x"48",x"66"),
  1170 => (x"d4",x"7b",x"70",x"98"),
  1171 => (x"2a",x"d0",x"4a",x"66"),
  1172 => (x"ff",x"c3",x"48",x"72"),
  1173 => (x"6b",x"7b",x"70",x"98"),
  1174 => (x"9d",x"ff",x"c3",x"4d"),
  1175 => (x"4c",x"ff",x"f0",x"c9"),
  1176 => (x"ad",x"b7",x"ff",x"c3"),
  1177 => (x"87",x"d8",x"c0",x"05"),
  1178 => (x"72",x"4a",x"ff",x"c3"),
  1179 => (x"72",x"4d",x"6b",x"7b"),
  1180 => (x"74",x"8c",x"c1",x"9d"),
  1181 => (x"c7",x"c0",x"02",x"9c"),
  1182 => (x"ad",x"b7",x"72",x"87"),
  1183 => (x"87",x"eb",x"ff",x"02"),
  1184 => (x"e1",x"27",x"1e",x"75"),
  1185 => (x"1e",x"00",x"00",x"19"),
  1186 => (x"00",x"00",x"3f",x"27"),
  1187 => (x"86",x"c8",x"0f",x"00"),
  1188 => (x"4d",x"26",x"48",x"75"),
  1189 => (x"4b",x"26",x"4c",x"26"),
  1190 => (x"4f",x"26",x"4a",x"26"),
  1191 => (x"5b",x"5a",x"5e",x"0e"),
  1192 => (x"e4",x"f6",x"c0",x"0e"),
  1193 => (x"c0",x"4b",x"c0",x"c0"),
  1194 => (x"7b",x"ff",x"c3",x"4a"),
  1195 => (x"c8",x"c3",x"82",x"c1"),
  1196 => (x"ff",x"04",x"aa",x"b7"),
  1197 => (x"4b",x"26",x"87",x"f3"),
  1198 => (x"4f",x"26",x"4a",x"26"),
  1199 => (x"5b",x"5a",x"5e",x"0e"),
  1200 => (x"c1",x"0e",x"5d",x"5c"),
  1201 => (x"c0",x"c0",x"c0",x"c0"),
  1202 => (x"f6",x"c0",x"4c",x"c0"),
  1203 => (x"4b",x"c0",x"c0",x"e4"),
  1204 => (x"00",x"12",x"9c",x"27"),
  1205 => (x"f8",x"c4",x"0f",x"00"),
  1206 => (x"1e",x"c0",x"4d",x"df"),
  1207 => (x"c1",x"f0",x"ff",x"c0"),
  1208 => (x"f8",x"27",x"1e",x"f7"),
  1209 => (x"0f",x"00",x"00",x"11"),
  1210 => (x"4a",x"70",x"86",x"c8"),
  1211 => (x"05",x"aa",x"b7",x"c1"),
  1212 => (x"72",x"87",x"dc",x"c1"),
  1213 => (x"13",x"7d",x"27",x"1e"),
  1214 => (x"27",x"1e",x"00",x"00"),
  1215 => (x"00",x"00",x"00",x"3f"),
  1216 => (x"c3",x"86",x"c8",x"0f"),
  1217 => (x"1e",x"74",x"7b",x"ff"),
  1218 => (x"c1",x"f0",x"e1",x"c0"),
  1219 => (x"f8",x"27",x"1e",x"e9"),
  1220 => (x"0f",x"00",x"00",x"11"),
  1221 => (x"4a",x"70",x"86",x"c8"),
  1222 => (x"c0",x"05",x"9a",x"72"),
  1223 => (x"1e",x"72",x"87",x"d8"),
  1224 => (x"00",x"13",x"73",x"27"),
  1225 => (x"3f",x"27",x"1e",x"00"),
  1226 => (x"0f",x"00",x"00",x"00"),
  1227 => (x"ff",x"c3",x"86",x"c8"),
  1228 => (x"c0",x"48",x"c1",x"7b"),
  1229 => (x"1e",x"72",x"87",x"f3"),
  1230 => (x"00",x"13",x"87",x"27"),
  1231 => (x"3f",x"27",x"1e",x"00"),
  1232 => (x"0f",x"00",x"00",x"00"),
  1233 => (x"9c",x"27",x"86",x"c8"),
  1234 => (x"0f",x"00",x"00",x"12"),
  1235 => (x"72",x"87",x"d0",x"c0"),
  1236 => (x"13",x"91",x"27",x"1e"),
  1237 => (x"27",x"1e",x"00",x"00"),
  1238 => (x"00",x"00",x"00",x"3f"),
  1239 => (x"c1",x"86",x"c8",x"0f"),
  1240 => (x"05",x"9d",x"75",x"8d"),
  1241 => (x"c0",x"87",x"f3",x"fd"),
  1242 => (x"26",x"4d",x"26",x"48"),
  1243 => (x"26",x"4b",x"26",x"4c"),
  1244 => (x"43",x"4f",x"26",x"4a"),
  1245 => (x"31",x"34",x"44",x"4d"),
  1246 => (x"0a",x"64",x"25",x"20"),
  1247 => (x"44",x"4d",x"43",x"00"),
  1248 => (x"25",x"20",x"35",x"35"),
  1249 => (x"43",x"00",x"0a",x"64"),
  1250 => (x"31",x"34",x"44",x"4d"),
  1251 => (x"0a",x"64",x"25",x"20"),
  1252 => (x"44",x"4d",x"43",x"00"),
  1253 => (x"25",x"20",x"35",x"35"),
  1254 => (x"0e",x"00",x"0a",x"64"),
  1255 => (x"5c",x"5b",x"5a",x"5e"),
  1256 => (x"ff",x"c0",x"0e",x"5d"),
  1257 => (x"4d",x"c1",x"c1",x"f0"),
  1258 => (x"c0",x"e4",x"f6",x"c0"),
  1259 => (x"ff",x"c3",x"4b",x"c0"),
  1260 => (x"14",x"2d",x"27",x"7b"),
  1261 => (x"27",x"1e",x"00",x"00"),
  1262 => (x"00",x"00",x"17",x"a3"),
  1263 => (x"d3",x"86",x"c4",x"0f"),
  1264 => (x"75",x"1e",x"c0",x"4c"),
  1265 => (x"11",x"f8",x"27",x"1e"),
  1266 => (x"c8",x"0f",x"00",x"00"),
  1267 => (x"72",x"4a",x"70",x"86"),
  1268 => (x"d8",x"c0",x"05",x"9a"),
  1269 => (x"27",x"1e",x"72",x"87"),
  1270 => (x"00",x"00",x"14",x"17"),
  1271 => (x"00",x"3f",x"27",x"1e"),
  1272 => (x"c8",x"0f",x"00",x"00"),
  1273 => (x"7b",x"ff",x"c3",x"86"),
  1274 => (x"e0",x"c0",x"48",x"c1"),
  1275 => (x"27",x"1e",x"72",x"87"),
  1276 => (x"00",x"00",x"14",x"22"),
  1277 => (x"00",x"3f",x"27",x"1e"),
  1278 => (x"c8",x"0f",x"00",x"00"),
  1279 => (x"12",x"9c",x"27",x"86"),
  1280 => (x"c1",x"0f",x"00",x"00"),
  1281 => (x"05",x"9c",x"74",x"8c"),
  1282 => (x"c0",x"87",x"f6",x"fe"),
  1283 => (x"26",x"4d",x"26",x"48"),
  1284 => (x"26",x"4b",x"26",x"4c"),
  1285 => (x"69",x"4f",x"26",x"4a"),
  1286 => (x"20",x"74",x"69",x"6e"),
  1287 => (x"20",x"0a",x"64",x"25"),
  1288 => (x"6e",x"69",x"00",x"20"),
  1289 => (x"25",x"20",x"74",x"69"),
  1290 => (x"20",x"20",x"0a",x"64"),
  1291 => (x"64",x"6d",x"43",x"00"),
  1292 => (x"69",x"6e",x"69",x"5f"),
  1293 => (x"0e",x"00",x"0a",x"74"),
  1294 => (x"5c",x"5b",x"5a",x"5e"),
  1295 => (x"c3",x"1e",x"0e",x"5d"),
  1296 => (x"f6",x"c0",x"4d",x"ff"),
  1297 => (x"4b",x"c0",x"c0",x"e4"),
  1298 => (x"00",x"12",x"9c",x"27"),
  1299 => (x"ea",x"c6",x"0f",x"00"),
  1300 => (x"f0",x"e1",x"c0",x"1e"),
  1301 => (x"27",x"1e",x"c8",x"c1"),
  1302 => (x"00",x"00",x"11",x"f8"),
  1303 => (x"70",x"86",x"c8",x"0f"),
  1304 => (x"27",x"1e",x"72",x"4a"),
  1305 => (x"00",x"00",x"15",x"c0"),
  1306 => (x"00",x"3f",x"27",x"1e"),
  1307 => (x"c8",x"0f",x"00",x"00"),
  1308 => (x"aa",x"b7",x"c1",x"86"),
  1309 => (x"87",x"cb",x"c0",x"02"),
  1310 => (x"00",x"13",x"9b",x"27"),
  1311 => (x"48",x"c0",x"0f",x"00"),
  1312 => (x"27",x"87",x"db",x"c3"),
  1313 => (x"00",x"00",x"11",x"97"),
  1314 => (x"74",x"4c",x"70",x"0f"),
  1315 => (x"ff",x"ff",x"cf",x"4a"),
  1316 => (x"b7",x"ea",x"c6",x"9a"),
  1317 => (x"db",x"c0",x"02",x"aa"),
  1318 => (x"27",x"1e",x"74",x"87"),
  1319 => (x"00",x"00",x"15",x"69"),
  1320 => (x"00",x"3f",x"27",x"1e"),
  1321 => (x"c8",x"0f",x"00",x"00"),
  1322 => (x"13",x"9b",x"27",x"86"),
  1323 => (x"c0",x"0f",x"00",x"00"),
  1324 => (x"87",x"ea",x"c2",x"48"),
  1325 => (x"49",x"76",x"7b",x"75"),
  1326 => (x"27",x"79",x"f1",x"c0"),
  1327 => (x"00",x"00",x"12",x"bc"),
  1328 => (x"72",x"4a",x"70",x"0f"),
  1329 => (x"eb",x"c1",x"02",x"9a"),
  1330 => (x"c0",x"1e",x"c0",x"87"),
  1331 => (x"fa",x"c1",x"f0",x"ff"),
  1332 => (x"11",x"f8",x"27",x"1e"),
  1333 => (x"c8",x"0f",x"00",x"00"),
  1334 => (x"74",x"4c",x"70",x"86"),
  1335 => (x"c3",x"c1",x"05",x"9c"),
  1336 => (x"27",x"1e",x"74",x"87"),
  1337 => (x"00",x"00",x"15",x"7e"),
  1338 => (x"00",x"3f",x"27",x"1e"),
  1339 => (x"c8",x"0f",x"00",x"00"),
  1340 => (x"6b",x"7b",x"75",x"86"),
  1341 => (x"74",x"9c",x"75",x"4c"),
  1342 => (x"15",x"8a",x"27",x"1e"),
  1343 => (x"27",x"1e",x"00",x"00"),
  1344 => (x"00",x"00",x"00",x"3f"),
  1345 => (x"75",x"86",x"c8",x"0f"),
  1346 => (x"75",x"7b",x"75",x"7b"),
  1347 => (x"74",x"7b",x"75",x"7b"),
  1348 => (x"9a",x"c0",x"c1",x"4a"),
  1349 => (x"c0",x"02",x"9a",x"72"),
  1350 => (x"48",x"c1",x"87",x"c5"),
  1351 => (x"c0",x"87",x"ff",x"c0"),
  1352 => (x"87",x"fa",x"c0",x"48"),
  1353 => (x"98",x"27",x"1e",x"74"),
  1354 => (x"1e",x"00",x"00",x"15"),
  1355 => (x"00",x"00",x"3f",x"27"),
  1356 => (x"86",x"c8",x"0f",x"00"),
  1357 => (x"b7",x"c2",x"49",x"6e"),
  1358 => (x"d3",x"c0",x"05",x"a9"),
  1359 => (x"15",x"a4",x"27",x"87"),
  1360 => (x"27",x"1e",x"00",x"00"),
  1361 => (x"00",x"00",x"00",x"3f"),
  1362 => (x"c0",x"86",x"c4",x"0f"),
  1363 => (x"87",x"ce",x"c0",x"48"),
  1364 => (x"88",x"c1",x"48",x"6e"),
  1365 => (x"6e",x"58",x"a6",x"c4"),
  1366 => (x"87",x"df",x"fd",x"05"),
  1367 => (x"26",x"26",x"48",x"c0"),
  1368 => (x"26",x"4c",x"26",x"4d"),
  1369 => (x"26",x"4a",x"26",x"4b"),
  1370 => (x"44",x"4d",x"43",x"4f"),
  1371 => (x"20",x"34",x"5f",x"38"),
  1372 => (x"70",x"73",x"65",x"72"),
  1373 => (x"65",x"73",x"6e",x"6f"),
  1374 => (x"64",x"25",x"20",x"3a"),
  1375 => (x"4d",x"43",x"00",x"0a"),
  1376 => (x"20",x"38",x"35",x"44"),
  1377 => (x"20",x"0a",x"64",x"25"),
  1378 => (x"4d",x"43",x"00",x"20"),
  1379 => (x"5f",x"38",x"35",x"44"),
  1380 => (x"64",x"25",x"20",x"32"),
  1381 => (x"00",x"20",x"20",x"0a"),
  1382 => (x"35",x"44",x"4d",x"43"),
  1383 => (x"64",x"25",x"20",x"38"),
  1384 => (x"00",x"20",x"20",x"0a"),
  1385 => (x"43",x"48",x"44",x"53"),
  1386 => (x"69",x"6e",x"49",x"20"),
  1387 => (x"6c",x"61",x"69",x"74"),
  1388 => (x"74",x"61",x"7a",x"69"),
  1389 => (x"20",x"6e",x"6f",x"69"),
  1390 => (x"6f",x"72",x"72",x"65"),
  1391 => (x"00",x"0a",x"21",x"72"),
  1392 => (x"5f",x"64",x"6d",x"63"),
  1393 => (x"38",x"44",x"4d",x"43"),
  1394 => (x"73",x"65",x"72",x"20"),
  1395 => (x"73",x"6e",x"6f",x"70"),
  1396 => (x"25",x"20",x"3a",x"65"),
  1397 => (x"0e",x"00",x"0a",x"64"),
  1398 => (x"5c",x"5b",x"5a",x"5e"),
  1399 => (x"f6",x"c0",x"0e",x"5d"),
  1400 => (x"4d",x"c0",x"c0",x"e4"),
  1401 => (x"c0",x"e4",x"f6",x"c0"),
  1402 => (x"88",x"27",x"4b",x"c4"),
  1403 => (x"49",x"00",x"00",x"1c"),
  1404 => (x"f6",x"c0",x"79",x"c1"),
  1405 => (x"49",x"c8",x"c0",x"e4"),
  1406 => (x"c7",x"79",x"e0",x"c0"),
  1407 => (x"27",x"7b",x"c3",x"4c"),
  1408 => (x"00",x"00",x"12",x"9c"),
  1409 => (x"c3",x"7b",x"c2",x"0f"),
  1410 => (x"1e",x"c0",x"7d",x"ff"),
  1411 => (x"c1",x"d0",x"e5",x"c0"),
  1412 => (x"f8",x"27",x"1e",x"c0"),
  1413 => (x"0f",x"00",x"00",x"11"),
  1414 => (x"4a",x"70",x"86",x"c8"),
  1415 => (x"05",x"aa",x"b7",x"c1"),
  1416 => (x"c1",x"87",x"c2",x"c0"),
  1417 => (x"ac",x"b7",x"c2",x"4c"),
  1418 => (x"87",x"c5",x"c0",x"05"),
  1419 => (x"f8",x"c0",x"48",x"c0"),
  1420 => (x"74",x"8c",x"c1",x"87"),
  1421 => (x"c4",x"ff",x"05",x"9c"),
  1422 => (x"14",x"37",x"27",x"87"),
  1423 => (x"27",x"0f",x"00",x"00"),
  1424 => (x"00",x"00",x"1c",x"8c"),
  1425 => (x"1c",x"88",x"27",x"58"),
  1426 => (x"05",x"bf",x"00",x"00"),
  1427 => (x"c1",x"87",x"d0",x"c0"),
  1428 => (x"f0",x"ff",x"c0",x"1e"),
  1429 => (x"27",x"1e",x"d0",x"c1"),
  1430 => (x"00",x"00",x"11",x"f8"),
  1431 => (x"c3",x"86",x"c8",x"0f"),
  1432 => (x"7b",x"c3",x"7d",x"ff"),
  1433 => (x"c1",x"7d",x"ff",x"c3"),
  1434 => (x"26",x"4d",x"26",x"48"),
  1435 => (x"26",x"4b",x"26",x"4c"),
  1436 => (x"1e",x"4f",x"26",x"4a"),
  1437 => (x"4f",x"26",x"48",x"c0"),
  1438 => (x"5b",x"5a",x"5e",x"0e"),
  1439 => (x"c8",x"0e",x"5d",x"5c"),
  1440 => (x"66",x"e0",x"c0",x"8e"),
  1441 => (x"e4",x"f6",x"c0",x"4d"),
  1442 => (x"76",x"4b",x"c0",x"c0"),
  1443 => (x"75",x"79",x"c0",x"49"),
  1444 => (x"66",x"e0",x"c0",x"1e"),
  1445 => (x"17",x"5d",x"27",x"1e"),
  1446 => (x"27",x"1e",x"00",x"00"),
  1447 => (x"00",x"00",x"00",x"3f"),
  1448 => (x"c3",x"86",x"cc",x"0f"),
  1449 => (x"f6",x"c0",x"7b",x"ff"),
  1450 => (x"49",x"c4",x"c0",x"e4"),
  1451 => (x"f6",x"c0",x"79",x"c2"),
  1452 => (x"49",x"c8",x"c0",x"e4"),
  1453 => (x"ff",x"c3",x"79",x"c1"),
  1454 => (x"1e",x"66",x"dc",x"7b"),
  1455 => (x"c1",x"f0",x"ff",x"c0"),
  1456 => (x"f8",x"27",x"1e",x"d1"),
  1457 => (x"0f",x"00",x"00",x"11"),
  1458 => (x"a6",x"c8",x"86",x"c8"),
  1459 => (x"02",x"66",x"c4",x"58"),
  1460 => (x"c4",x"87",x"d8",x"c0"),
  1461 => (x"e0",x"c0",x"1e",x"66"),
  1462 => (x"3d",x"27",x"1e",x"66"),
  1463 => (x"1e",x"00",x"00",x"17"),
  1464 => (x"00",x"00",x"3f",x"27"),
  1465 => (x"86",x"cc",x"0f",x"00"),
  1466 => (x"c5",x"87",x"c4",x"c1"),
  1467 => (x"4c",x"df",x"cd",x"ee"),
  1468 => (x"6b",x"7b",x"ff",x"c3"),
  1469 => (x"9a",x"ff",x"c3",x"4a"),
  1470 => (x"aa",x"b7",x"fe",x"c3"),
  1471 => (x"87",x"dc",x"c0",x"05"),
  1472 => (x"20",x"27",x"4a",x"c0"),
  1473 => (x"0f",x"00",x"00",x"11"),
  1474 => (x"85",x"c4",x"7d",x"70"),
  1475 => (x"c0",x"c2",x"82",x"c1"),
  1476 => (x"ff",x"04",x"aa",x"b7"),
  1477 => (x"4c",x"c1",x"87",x"ec"),
  1478 => (x"79",x"c1",x"49",x"76"),
  1479 => (x"9c",x"74",x"8c",x"c1"),
  1480 => (x"87",x"cc",x"ff",x"05"),
  1481 => (x"c0",x"7b",x"ff",x"c3"),
  1482 => (x"c4",x"c0",x"e4",x"f6"),
  1483 => (x"6e",x"79",x"c3",x"49"),
  1484 => (x"26",x"86",x"c8",x"48"),
  1485 => (x"26",x"4c",x"26",x"4d"),
  1486 => (x"26",x"4a",x"26",x"4b"),
  1487 => (x"61",x"65",x"52",x"4f"),
  1488 => (x"6f",x"63",x"20",x"64"),
  1489 => (x"6e",x"61",x"6d",x"6d"),
  1490 => (x"61",x"66",x"20",x"64"),
  1491 => (x"64",x"65",x"6c",x"69"),
  1492 => (x"20",x"74",x"61",x"20"),
  1493 => (x"28",x"20",x"64",x"25"),
  1494 => (x"0a",x"29",x"64",x"25"),
  1495 => (x"5f",x"64",x"73",x"00"),
  1496 => (x"64",x"61",x"65",x"72"),
  1497 => (x"63",x"65",x"73",x"5f"),
  1498 => (x"20",x"72",x"6f",x"74"),
  1499 => (x"20",x"2c",x"64",x"25"),
  1500 => (x"00",x"0a",x"64",x"25"),
  1501 => (x"1e",x"1e",x"72",x"1e"),
  1502 => (x"c0",x"e8",x"f6",x"c0"),
  1503 => (x"48",x"6a",x"4a",x"c0"),
  1504 => (x"c4",x"98",x"c0",x"c4"),
  1505 => (x"05",x"6e",x"58",x"a6"),
  1506 => (x"6a",x"87",x"cd",x"c0"),
  1507 => (x"98",x"c0",x"c4",x"48"),
  1508 => (x"6e",x"58",x"a6",x"c4"),
  1509 => (x"87",x"f3",x"ff",x"02"),
  1510 => (x"cc",x"7a",x"66",x"cc"),
  1511 => (x"26",x"26",x"48",x"66"),
  1512 => (x"0e",x"4f",x"26",x"4a"),
  1513 => (x"5c",x"5b",x"5a",x"5e"),
  1514 => (x"4b",x"66",x"d0",x"0e"),
  1515 => (x"4a",x"13",x"4c",x"c0"),
  1516 => (x"c0",x"c0",x"c0",x"c1"),
  1517 => (x"c0",x"c4",x"92",x"c0"),
  1518 => (x"72",x"4a",x"92",x"b7"),
  1519 => (x"17",x"74",x"27",x"1e"),
  1520 => (x"c4",x"0f",x"00",x"00"),
  1521 => (x"72",x"84",x"c1",x"86"),
  1522 => (x"e1",x"ff",x"05",x"9a"),
  1523 => (x"26",x"48",x"74",x"87"),
  1524 => (x"26",x"4b",x"26",x"4c"),
  1525 => (x"0e",x"4f",x"26",x"4a"),
  1526 => (x"5c",x"5b",x"5a",x"5e"),
  1527 => (x"8e",x"c8",x"0e",x"5d"),
  1528 => (x"4c",x"66",x"e0",x"c0"),
  1529 => (x"76",x"4a",x"66",x"dc"),
  1530 => (x"c0",x"79",x"c0",x"49"),
  1531 => (x"c1",x"06",x"ac",x"b7"),
  1532 => (x"4b",x"12",x"87",x"e2"),
  1533 => (x"8c",x"c1",x"33",x"c8"),
  1534 => (x"06",x"ac",x"b7",x"c0"),
  1535 => (x"12",x"87",x"c8",x"c0"),
  1536 => (x"58",x"a6",x"c8",x"48"),
  1537 => (x"c4",x"87",x"c5",x"c0"),
  1538 => (x"79",x"c0",x"49",x"a6"),
  1539 => (x"66",x"c4",x"4b",x"73"),
  1540 => (x"c1",x"33",x"c8",x"b3"),
  1541 => (x"ac",x"b7",x"c0",x"8c"),
  1542 => (x"87",x"c5",x"c0",x"06"),
  1543 => (x"c2",x"c0",x"4d",x"12"),
  1544 => (x"73",x"4d",x"c0",x"87"),
  1545 => (x"c8",x"b3",x"75",x"4b"),
  1546 => (x"c0",x"8c",x"c1",x"33"),
  1547 => (x"c0",x"06",x"ac",x"b7"),
  1548 => (x"48",x"12",x"87",x"c8"),
  1549 => (x"c0",x"58",x"a6",x"c8"),
  1550 => (x"a6",x"c4",x"87",x"c5"),
  1551 => (x"73",x"79",x"c0",x"49"),
  1552 => (x"b3",x"66",x"c4",x"4b"),
  1553 => (x"80",x"6e",x"48",x"73"),
  1554 => (x"c1",x"58",x"a6",x"c4"),
  1555 => (x"ac",x"b7",x"c0",x"8c"),
  1556 => (x"87",x"de",x"fe",x"01"),
  1557 => (x"86",x"c8",x"48",x"6e"),
  1558 => (x"4c",x"26",x"4d",x"26"),
  1559 => (x"4a",x"26",x"4b",x"26"),
  1560 => (x"68",x"43",x"4f",x"26"),
  1561 => (x"73",x"6b",x"63",x"65"),
  1562 => (x"74",x"20",x"6d",x"75"),
  1563 => (x"64",x"25",x"20",x"6f"),
  1564 => (x"64",x"25",x"20",x"3a"),
  1565 => (x"65",x"52",x"00",x"0a"),
  1566 => (x"6f",x"20",x"64",x"61"),
  1567 => (x"42",x"4d",x"20",x"66"),
  1568 => (x"61",x"66",x"20",x"52"),
  1569 => (x"64",x"65",x"6c",x"69"),
  1570 => (x"6f",x"4e",x"00",x"0a"),
  1571 => (x"72",x"61",x"70",x"20"),
  1572 => (x"69",x"74",x"69",x"74"),
  1573 => (x"73",x"20",x"6e",x"6f"),
  1574 => (x"61",x"6e",x"67",x"69"),
  1575 => (x"65",x"72",x"75",x"74"),
  1576 => (x"75",x"6f",x"66",x"20"),
  1577 => (x"00",x"0a",x"64",x"6e"),
  1578 => (x"73",x"52",x"42",x"4d"),
  1579 => (x"3a",x"65",x"7a",x"69"),
  1580 => (x"2c",x"64",x"25",x"20"),
  1581 => (x"72",x"61",x"70",x"20"),
  1582 => (x"69",x"74",x"69",x"74"),
  1583 => (x"69",x"73",x"6e",x"6f"),
  1584 => (x"20",x"3a",x"65",x"7a"),
  1585 => (x"20",x"2c",x"64",x"25"),
  1586 => (x"73",x"66",x"66",x"6f"),
  1587 => (x"6f",x"20",x"74",x"65"),
  1588 => (x"69",x"73",x"20",x"66"),
  1589 => (x"25",x"20",x"3a",x"67"),
  1590 => (x"73",x"20",x"2c",x"64"),
  1591 => (x"30",x"20",x"67",x"69"),
  1592 => (x"0a",x"78",x"25",x"78"),
  1593 => (x"61",x"65",x"52",x"00"),
  1594 => (x"67",x"6e",x"69",x"64"),
  1595 => (x"6f",x"6f",x"62",x"20"),
  1596 => (x"65",x"73",x"20",x"74"),
  1597 => (x"72",x"6f",x"74",x"63"),
  1598 => (x"0a",x"64",x"25",x"20"),
  1599 => (x"61",x"65",x"52",x"00"),
  1600 => (x"6f",x"62",x"20",x"64"),
  1601 => (x"73",x"20",x"74",x"6f"),
  1602 => (x"6f",x"74",x"63",x"65"),
  1603 => (x"72",x"66",x"20",x"72"),
  1604 => (x"66",x"20",x"6d",x"6f"),
  1605 => (x"74",x"73",x"72",x"69"),
  1606 => (x"72",x"61",x"70",x"20"),
  1607 => (x"69",x"74",x"69",x"74"),
  1608 => (x"00",x"0a",x"6e",x"6f"),
  1609 => (x"75",x"73",x"6e",x"55"),
  1610 => (x"72",x"6f",x"70",x"70"),
  1611 => (x"20",x"64",x"65",x"74"),
  1612 => (x"74",x"72",x"61",x"70"),
  1613 => (x"6f",x"69",x"74",x"69"),
  1614 => (x"79",x"74",x"20",x"6e"),
  1615 => (x"0d",x"21",x"65",x"70"),
  1616 => (x"54",x"41",x"46",x"00"),
  1617 => (x"20",x"20",x"32",x"33"),
  1618 => (x"65",x"52",x"00",x"20"),
  1619 => (x"6e",x"69",x"64",x"61"),
  1620 => (x"42",x"4d",x"20",x"67"),
  1621 => (x"4d",x"00",x"0a",x"52"),
  1622 => (x"73",x"20",x"52",x"42"),
  1623 => (x"65",x"63",x"63",x"75"),
  1624 => (x"75",x"66",x"73",x"73"),
  1625 => (x"20",x"79",x"6c",x"6c"),
  1626 => (x"64",x"61",x"65",x"72"),
  1627 => (x"41",x"46",x"00",x"0a"),
  1628 => (x"20",x"36",x"31",x"54"),
  1629 => (x"46",x"00",x"20",x"20"),
  1630 => (x"32",x"33",x"54",x"41"),
  1631 => (x"00",x"20",x"20",x"20"),
  1632 => (x"74",x"72",x"61",x"50"),
  1633 => (x"6f",x"69",x"74",x"69"),
  1634 => (x"75",x"6f",x"63",x"6e"),
  1635 => (x"25",x"20",x"74",x"6e"),
  1636 => (x"48",x"00",x"0a",x"64"),
  1637 => (x"69",x"74",x"6e",x"75"),
  1638 => (x"66",x"20",x"67",x"6e"),
  1639 => (x"66",x"20",x"72",x"6f"),
  1640 => (x"73",x"65",x"6c",x"69"),
  1641 => (x"65",x"74",x"73",x"79"),
  1642 => (x"46",x"00",x"0a",x"6d"),
  1643 => (x"32",x"33",x"54",x"41"),
  1644 => (x"00",x"20",x"20",x"20"),
  1645 => (x"31",x"54",x"41",x"46"),
  1646 => (x"20",x"20",x"20",x"36"),
  1647 => (x"75",x"6c",x"43",x"00"),
  1648 => (x"72",x"65",x"74",x"73"),
  1649 => (x"7a",x"69",x"73",x"20"),
  1650 => (x"25",x"20",x"3a",x"65"),
  1651 => (x"43",x"20",x"2c",x"64"),
  1652 => (x"74",x"73",x"75",x"6c"),
  1653 => (x"6d",x"20",x"72",x"65"),
  1654 => (x"2c",x"6b",x"73",x"61"),
  1655 => (x"0a",x"64",x"25",x"20"),
  1656 => (x"74",x"6f",x"47",x"00"),
  1657 => (x"73",x"65",x"72",x"20"),
  1658 => (x"20",x"74",x"6c",x"75"),
  1659 => (x"0a",x"20",x"64",x"25"),
  1660 => (x"0a",x"20",x"64",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
