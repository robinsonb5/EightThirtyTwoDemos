
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"2c",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"29"),
    10 => (x"87",x"fd",x"00",x"4f"),
    11 => (x"e0",x"f2",x"c3",x"4f"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"e0",x"f2",x"c3"),
    14 => (x"48",x"e8",x"cf",x"c1"),
    15 => (x"03",x"89",x"d0",x"89"),
    16 => (x"40",x"40",x"40",x"c0"),
    17 => (x"d0",x"87",x"f6",x"40"),
    18 => (x"50",x"c0",x"05",x"81"),
    19 => (x"f9",x"05",x"89",x"c1"),
    20 => (x"e6",x"cf",x"c1",x"87"),
    21 => (x"e6",x"cf",x"c1",x"4d"),
    22 => (x"02",x"ad",x"74",x"4c"),
    23 => (x"0f",x"24",x"87",x"c4"),
    24 => (x"ed",x"cd",x"87",x"f7"),
    25 => (x"e6",x"cf",x"c1",x"87"),
    26 => (x"e6",x"cf",x"c1",x"4d"),
    27 => (x"02",x"ad",x"74",x"4c"),
    28 => (x"8c",x"c4",x"87",x"c6"),
    29 => (x"87",x"f5",x"0f",x"6c"),
    30 => (x"0e",x"87",x"fd",x"00"),
    31 => (x"5d",x"5c",x"5b",x"5e"),
    32 => (x"71",x"86",x"fc",x"0e"),
    33 => (x"66",x"e0",x"c0",x"4a"),
    34 => (x"e8",x"cf",x"c1",x"4c"),
    35 => (x"72",x"7e",x"c0",x"4b"),
    36 => (x"87",x"ce",x"05",x"9a"),
    37 => (x"4b",x"e9",x"cf",x"c1"),
    38 => (x"48",x"e8",x"cf",x"c1"),
    39 => (x"c1",x"50",x"f0",x"c0"),
    40 => (x"9a",x"72",x"87",x"d1"),
    41 => (x"87",x"e8",x"c0",x"02"),
    42 => (x"72",x"4d",x"66",x"d4"),
    43 => (x"75",x"49",x"72",x"1e"),
    44 => (x"87",x"f9",x"ca",x"4a"),
    45 => (x"e4",x"c4",x"4a",x"26"),
    46 => (x"71",x"53",x"11",x"81"),
    47 => (x"75",x"49",x"72",x"1e"),
    48 => (x"87",x"e9",x"ca",x"4a"),
    49 => (x"49",x"26",x"4a",x"70"),
    50 => (x"9a",x"72",x"8c",x"c1"),
    51 => (x"87",x"db",x"ff",x"05"),
    52 => (x"06",x"ac",x"b7",x"c0"),
    53 => (x"e4",x"c0",x"87",x"dd"),
    54 => (x"87",x"c5",x"02",x"66"),
    55 => (x"c3",x"4a",x"f0",x"c0"),
    56 => (x"4a",x"e0",x"c0",x"87"),
    57 => (x"7a",x"97",x"0a",x"73"),
    58 => (x"8c",x"83",x"c1",x"0a"),
    59 => (x"01",x"ac",x"b7",x"c0"),
    60 => (x"c1",x"87",x"e3",x"ff"),
    61 => (x"02",x"ab",x"e8",x"cf"),
    62 => (x"66",x"d8",x"87",x"de"),
    63 => (x"1e",x"66",x"dc",x"4c"),
    64 => (x"6b",x"97",x"8b",x"c1"),
    65 => (x"c4",x"0f",x"74",x"49"),
    66 => (x"c1",x"48",x"6e",x"86"),
    67 => (x"58",x"a6",x"c4",x"80"),
    68 => (x"ab",x"e8",x"cf",x"c1"),
    69 => (x"87",x"e5",x"ff",x"05"),
    70 => (x"8e",x"fc",x"48",x"6e"),
    71 => (x"4c",x"26",x"4d",x"26"),
    72 => (x"4f",x"26",x"4b",x"26"),
    73 => (x"33",x"32",x"31",x"30"),
    74 => (x"37",x"36",x"35",x"34"),
    75 => (x"42",x"41",x"39",x"38"),
    76 => (x"46",x"45",x"44",x"43"),
    77 => (x"5b",x"5e",x"0e",x"00"),
    78 => (x"71",x"0e",x"5d",x"5c"),
    79 => (x"13",x"4d",x"ff",x"4b"),
    80 => (x"02",x"9c",x"74",x"4c"),
    81 => (x"85",x"c1",x"87",x"d8"),
    82 => (x"74",x"1e",x"66",x"d4"),
    83 => (x"0f",x"66",x"d4",x"49"),
    84 => (x"a8",x"74",x"86",x"c4"),
    85 => (x"13",x"87",x"c7",x"05"),
    86 => (x"05",x"9c",x"74",x"4c"),
    87 => (x"48",x"75",x"87",x"e8"),
    88 => (x"4c",x"26",x"4d",x"26"),
    89 => (x"4f",x"26",x"4b",x"26"),
    90 => (x"5c",x"5b",x"5e",x"0e"),
    91 => (x"86",x"e8",x"0e",x"5d"),
    92 => (x"c0",x"59",x"a6",x"c4"),
    93 => (x"c0",x"4d",x"66",x"e8"),
    94 => (x"48",x"a6",x"c8",x"4c"),
    95 => (x"97",x"6e",x"78",x"c0"),
    96 => (x"48",x"6e",x"4b",x"bf"),
    97 => (x"a6",x"c4",x"80",x"c1"),
    98 => (x"02",x"9b",x"73",x"58"),
    99 => (x"c8",x"87",x"d3",x"c6"),
   100 => (x"db",x"c5",x"02",x"66"),
   101 => (x"48",x"a6",x"cc",x"87"),
   102 => (x"80",x"fc",x"78",x"c0"),
   103 => (x"4a",x"73",x"78",x"c0"),
   104 => (x"02",x"8a",x"e0",x"c0"),
   105 => (x"c3",x"87",x"c6",x"c3"),
   106 => (x"c0",x"c3",x"02",x"8a"),
   107 => (x"02",x"8a",x"c2",x"87"),
   108 => (x"c2",x"87",x"e8",x"c2"),
   109 => (x"f4",x"c2",x"02",x"8a"),
   110 => (x"02",x"8a",x"c4",x"87"),
   111 => (x"c2",x"87",x"ee",x"c2"),
   112 => (x"e8",x"c2",x"02",x"8a"),
   113 => (x"02",x"8a",x"c3",x"87"),
   114 => (x"d4",x"87",x"ea",x"c2"),
   115 => (x"f6",x"c0",x"02",x"8a"),
   116 => (x"02",x"8a",x"d4",x"87"),
   117 => (x"ca",x"87",x"c0",x"c1"),
   118 => (x"f2",x"c0",x"02",x"8a"),
   119 => (x"02",x"8a",x"c1",x"87"),
   120 => (x"c1",x"87",x"e1",x"c1"),
   121 => (x"87",x"df",x"02",x"8a"),
   122 => (x"c1",x"02",x"8a",x"c8"),
   123 => (x"8a",x"c4",x"87",x"ce"),
   124 => (x"87",x"e3",x"c0",x"02"),
   125 => (x"c0",x"02",x"8a",x"c3"),
   126 => (x"8a",x"c2",x"87",x"e5"),
   127 => (x"c3",x"87",x"c8",x"02"),
   128 => (x"87",x"d3",x"02",x"8a"),
   129 => (x"cc",x"87",x"fa",x"c1"),
   130 => (x"78",x"ca",x"48",x"a6"),
   131 => (x"cc",x"87",x"d2",x"c2"),
   132 => (x"78",x"c2",x"48",x"a6"),
   133 => (x"cc",x"87",x"ca",x"c2"),
   134 => (x"78",x"d0",x"48",x"a6"),
   135 => (x"c0",x"87",x"c2",x"c2"),
   136 => (x"c0",x"1e",x"66",x"f0"),
   137 => (x"c4",x"1e",x"66",x"f0"),
   138 => (x"c4",x"4a",x"75",x"85"),
   139 => (x"fc",x"49",x"6a",x"8a"),
   140 => (x"86",x"c8",x"87",x"c3"),
   141 => (x"a4",x"71",x"49",x"70"),
   142 => (x"87",x"e5",x"c1",x"4c"),
   143 => (x"c1",x"48",x"a6",x"c8"),
   144 => (x"87",x"dd",x"c1",x"78"),
   145 => (x"1e",x"66",x"f0",x"c0"),
   146 => (x"4a",x"75",x"85",x"c4"),
   147 => (x"49",x"6a",x"8a",x"c4"),
   148 => (x"0f",x"66",x"f0",x"c0"),
   149 => (x"84",x"c1",x"86",x"c4"),
   150 => (x"c0",x"87",x"c6",x"c1"),
   151 => (x"c0",x"1e",x"66",x"f0"),
   152 => (x"f0",x"c0",x"49",x"e5"),
   153 => (x"86",x"c4",x"0f",x"66"),
   154 => (x"f4",x"c0",x"84",x"c1"),
   155 => (x"48",x"a6",x"c8",x"87"),
   156 => (x"ec",x"c0",x"78",x"c1"),
   157 => (x"48",x"a6",x"d0",x"87"),
   158 => (x"80",x"f8",x"78",x"c1"),
   159 => (x"e0",x"c0",x"78",x"c1"),
   160 => (x"ab",x"f0",x"c0",x"87"),
   161 => (x"c0",x"87",x"da",x"06"),
   162 => (x"d4",x"03",x"ab",x"f9"),
   163 => (x"49",x"66",x"d4",x"87"),
   164 => (x"4a",x"73",x"91",x"ca"),
   165 => (x"d4",x"8a",x"f0",x"c0"),
   166 => (x"a1",x"72",x"48",x"a6"),
   167 => (x"c1",x"80",x"f4",x"78"),
   168 => (x"02",x"66",x"cc",x"78"),
   169 => (x"c4",x"87",x"ea",x"c1"),
   170 => (x"c4",x"49",x"75",x"85"),
   171 => (x"69",x"48",x"a6",x"89"),
   172 => (x"ab",x"e4",x"c1",x"78"),
   173 => (x"c4",x"87",x"d8",x"05"),
   174 => (x"b7",x"c0",x"48",x"66"),
   175 => (x"87",x"cf",x"03",x"a8"),
   176 => (x"c1",x"49",x"ed",x"c0"),
   177 => (x"66",x"c4",x"87",x"fb"),
   178 => (x"88",x"08",x"c0",x"48"),
   179 => (x"d0",x"58",x"a6",x"c8"),
   180 => (x"66",x"d8",x"1e",x"66"),
   181 => (x"66",x"f8",x"c0",x"1e"),
   182 => (x"66",x"f8",x"c0",x"1e"),
   183 => (x"1e",x"66",x"dc",x"1e"),
   184 => (x"f6",x"49",x"66",x"d8"),
   185 => (x"86",x"d4",x"87",x"d5"),
   186 => (x"a4",x"71",x"49",x"70"),
   187 => (x"87",x"e1",x"c0",x"4c"),
   188 => (x"05",x"ab",x"e5",x"c0"),
   189 => (x"a6",x"d0",x"87",x"cf"),
   190 => (x"c4",x"78",x"c0",x"48"),
   191 => (x"f4",x"78",x"c0",x"80"),
   192 => (x"cc",x"78",x"c1",x"80"),
   193 => (x"66",x"f0",x"c0",x"87"),
   194 => (x"c0",x"49",x"73",x"1e"),
   195 => (x"c4",x"0f",x"66",x"f0"),
   196 => (x"bf",x"97",x"6e",x"86"),
   197 => (x"c1",x"48",x"6e",x"4b"),
   198 => (x"58",x"a6",x"c4",x"80"),
   199 => (x"f9",x"05",x"9b",x"73"),
   200 => (x"48",x"74",x"87",x"ed"),
   201 => (x"4d",x"26",x"8e",x"e8"),
   202 => (x"4b",x"26",x"4c",x"26"),
   203 => (x"c0",x"1e",x"4f",x"26"),
   204 => (x"1e",x"c1",x"cd",x"1e"),
   205 => (x"d0",x"1e",x"a6",x"d0"),
   206 => (x"eb",x"f8",x"49",x"66"),
   207 => (x"26",x"8e",x"f4",x"87"),
   208 => (x"86",x"fc",x"1e",x"4f"),
   209 => (x"c0",x"ff",x"4a",x"71"),
   210 => (x"c4",x"48",x"69",x"49"),
   211 => (x"a6",x"c4",x"98",x"c0"),
   212 => (x"f4",x"02",x"6e",x"58"),
   213 => (x"48",x"79",x"72",x"87"),
   214 => (x"4f",x"26",x"8e",x"fc"),
   215 => (x"12",x"1e",x"72",x"1e"),
   216 => (x"c4",x"02",x"11",x"48"),
   217 => (x"f6",x"02",x"88",x"87"),
   218 => (x"26",x"4a",x"26",x"87"),
   219 => (x"1e",x"73",x"1e",x"4f"),
   220 => (x"c0",x"02",x"9a",x"72"),
   221 => (x"48",x"c0",x"87",x"e7"),
   222 => (x"a9",x"72",x"4b",x"c1"),
   223 => (x"72",x"87",x"d1",x"06"),
   224 => (x"87",x"c9",x"06",x"82"),
   225 => (x"a9",x"72",x"83",x"73"),
   226 => (x"c3",x"87",x"f4",x"01"),
   227 => (x"3a",x"b2",x"c1",x"87"),
   228 => (x"89",x"03",x"a9",x"72"),
   229 => (x"c1",x"07",x"80",x"73"),
   230 => (x"f3",x"05",x"2b",x"2a"),
   231 => (x"26",x"4b",x"26",x"87"),
   232 => (x"1e",x"75",x"1e",x"4f"),
   233 => (x"b7",x"71",x"4d",x"c4"),
   234 => (x"b9",x"ff",x"04",x"a1"),
   235 => (x"bd",x"c3",x"81",x"c1"),
   236 => (x"a2",x"b7",x"72",x"07"),
   237 => (x"c1",x"ba",x"ff",x"04"),
   238 => (x"07",x"bd",x"c1",x"82"),
   239 => (x"c1",x"87",x"ee",x"fe"),
   240 => (x"b8",x"ff",x"04",x"2d"),
   241 => (x"2d",x"07",x"80",x"c1"),
   242 => (x"c1",x"b9",x"ff",x"04"),
   243 => (x"4d",x"26",x"07",x"81"),
   244 => (x"5e",x"0e",x"4f",x"26"),
   245 => (x"0e",x"5d",x"5c",x"5b"),
   246 => (x"c1",x"86",x"dc",x"ff"),
   247 => (x"c3",x"48",x"fc",x"cf"),
   248 => (x"c1",x"78",x"c0",x"f0"),
   249 => (x"c3",x"48",x"f8",x"cf"),
   250 => (x"48",x"78",x"f0",x"f0"),
   251 => (x"78",x"c0",x"f0",x"c3"),
   252 => (x"48",x"f4",x"f0",x"c3"),
   253 => (x"80",x"c4",x"78",x"c0"),
   254 => (x"80",x"c4",x"78",x"c2"),
   255 => (x"71",x"78",x"e8",x"c0"),
   256 => (x"dc",x"ee",x"c0",x"1e"),
   257 => (x"c0",x"f1",x"c3",x"48"),
   258 => (x"20",x"41",x"20",x"49"),
   259 => (x"20",x"41",x"20",x"41"),
   260 => (x"20",x"41",x"20",x"41"),
   261 => (x"10",x"41",x"20",x"41"),
   262 => (x"10",x"51",x"10",x"51"),
   263 => (x"71",x"49",x"26",x"51"),
   264 => (x"fc",x"ee",x"c0",x"1e"),
   265 => (x"e0",x"f1",x"c3",x"48"),
   266 => (x"20",x"41",x"20",x"49"),
   267 => (x"20",x"41",x"20",x"41"),
   268 => (x"20",x"41",x"20",x"41"),
   269 => (x"10",x"41",x"20",x"41"),
   270 => (x"10",x"51",x"10",x"51"),
   271 => (x"c1",x"49",x"26",x"51"),
   272 => (x"ca",x"48",x"f4",x"ec"),
   273 => (x"dc",x"ef",x"c0",x"78"),
   274 => (x"87",x"e2",x"fb",x"1e"),
   275 => (x"1e",x"e0",x"ef",x"c0"),
   276 => (x"c0",x"87",x"db",x"fb"),
   277 => (x"fb",x"1e",x"d0",x"f0"),
   278 => (x"86",x"cc",x"87",x"d4"),
   279 => (x"bf",x"c0",x"e8",x"c0"),
   280 => (x"c0",x"87",x"d2",x"02"),
   281 => (x"fb",x"1e",x"c8",x"e8"),
   282 => (x"e8",x"c0",x"87",x"c4"),
   283 => (x"fd",x"fa",x"1e",x"f4"),
   284 => (x"d0",x"86",x"c8",x"87"),
   285 => (x"f8",x"e8",x"c0",x"87"),
   286 => (x"87",x"f2",x"fa",x"1e"),
   287 => (x"1e",x"e8",x"e9",x"c0"),
   288 => (x"c8",x"87",x"eb",x"fa"),
   289 => (x"c4",x"e8",x"c0",x"86"),
   290 => (x"f0",x"c0",x"1e",x"bf"),
   291 => (x"dd",x"fa",x"1e",x"d4"),
   292 => (x"c3",x"86",x"c8",x"87"),
   293 => (x"ff",x"48",x"e8",x"ef"),
   294 => (x"c4",x"78",x"bf",x"c8"),
   295 => (x"78",x"c1",x"48",x"a6"),
   296 => (x"bf",x"c4",x"e8",x"c0"),
   297 => (x"a8",x"b7",x"c0",x"48"),
   298 => (x"87",x"f7",x"c8",x"06"),
   299 => (x"d0",x"48",x"a6",x"c8"),
   300 => (x"80",x"c8",x"58",x"a6"),
   301 => (x"c8",x"58",x"a6",x"d8"),
   302 => (x"58",x"a6",x"c4",x"80"),
   303 => (x"48",x"c8",x"d0",x"c1"),
   304 => (x"c1",x"50",x"c1",x"c1"),
   305 => (x"c0",x"48",x"c4",x"d0"),
   306 => (x"c8",x"d0",x"c1",x"78"),
   307 => (x"c1",x"49",x"bf",x"97"),
   308 => (x"c0",x"02",x"a9",x"c1"),
   309 => (x"a6",x"dc",x"87",x"c8"),
   310 => (x"c0",x"78",x"c0",x"48"),
   311 => (x"a6",x"dc",x"87",x"c5"),
   312 => (x"c1",x"78",x"c1",x"48"),
   313 => (x"48",x"bf",x"c4",x"d0"),
   314 => (x"c1",x"b0",x"66",x"dc"),
   315 => (x"c1",x"58",x"c8",x"d0"),
   316 => (x"c1",x"48",x"cc",x"d0"),
   317 => (x"a6",x"d8",x"50",x"c2"),
   318 => (x"c8",x"78",x"c2",x"48"),
   319 => (x"c0",x"78",x"c3",x"80"),
   320 => (x"c3",x"48",x"cc",x"ea"),
   321 => (x"20",x"49",x"c0",x"f2"),
   322 => (x"20",x"41",x"20",x"41"),
   323 => (x"20",x"41",x"20",x"41"),
   324 => (x"20",x"41",x"20",x"41"),
   325 => (x"10",x"51",x"10",x"41"),
   326 => (x"d0",x"51",x"10",x"51"),
   327 => (x"78",x"c1",x"48",x"a6"),
   328 => (x"1e",x"c0",x"f2",x"c3"),
   329 => (x"49",x"e0",x"f1",x"c3"),
   330 => (x"87",x"c4",x"f9",x"c0"),
   331 => (x"98",x"70",x"86",x"c4"),
   332 => (x"87",x"c8",x"c0",x"05"),
   333 => (x"c1",x"48",x"a6",x"dc"),
   334 => (x"87",x"c5",x"c0",x"78"),
   335 => (x"c0",x"48",x"a6",x"dc"),
   336 => (x"c4",x"d0",x"c1",x"78"),
   337 => (x"78",x"66",x"dc",x"48"),
   338 => (x"c3",x"48",x"66",x"d8"),
   339 => (x"c0",x"03",x"a8",x"b7"),
   340 => (x"66",x"d8",x"87",x"ed"),
   341 => (x"71",x"91",x"c5",x"49"),
   342 => (x"cc",x"88",x"c3",x"48"),
   343 => (x"66",x"cc",x"58",x"a6"),
   344 => (x"c0",x"1e",x"c3",x"1e"),
   345 => (x"c0",x"49",x"66",x"e0"),
   346 => (x"c8",x"87",x"c9",x"f5"),
   347 => (x"48",x"66",x"d8",x"86"),
   348 => (x"a6",x"dc",x"80",x"c1"),
   349 => (x"48",x"66",x"d8",x"58"),
   350 => (x"04",x"a8",x"b7",x"c3"),
   351 => (x"c8",x"87",x"d3",x"ff"),
   352 => (x"66",x"dc",x"1e",x"66"),
   353 => (x"d8",x"d3",x"c1",x"1e"),
   354 => (x"d0",x"d0",x"c1",x"1e"),
   355 => (x"f6",x"f4",x"c0",x"49"),
   356 => (x"c1",x"86",x"cc",x"87"),
   357 => (x"4c",x"bf",x"f8",x"cf"),
   358 => (x"bf",x"f8",x"cf",x"c1"),
   359 => (x"1e",x"72",x"4b",x"bf"),
   360 => (x"bf",x"f8",x"cf",x"c1"),
   361 => (x"c0",x"49",x"73",x"48"),
   362 => (x"20",x"4a",x"a1",x"f0"),
   363 => (x"05",x"aa",x"71",x"41"),
   364 => (x"26",x"87",x"f8",x"ff"),
   365 => (x"49",x"a4",x"cc",x"4a"),
   366 => (x"a3",x"cc",x"79",x"c5"),
   367 => (x"6c",x"7d",x"69",x"4d"),
   368 => (x"d0",x"49",x"73",x"7b"),
   369 => (x"a3",x"c4",x"87",x"cf"),
   370 => (x"c0",x"05",x"69",x"49"),
   371 => (x"a3",x"c8",x"87",x"e5"),
   372 => (x"71",x"7d",x"c6",x"49"),
   373 => (x"4a",x"a4",x"c8",x"1e"),
   374 => (x"f1",x"c0",x"49",x"6a"),
   375 => (x"cf",x"c1",x"87",x"f5"),
   376 => (x"7b",x"bf",x"bf",x"f8"),
   377 => (x"1e",x"ca",x"1e",x"75"),
   378 => (x"f3",x"c0",x"49",x"6d"),
   379 => (x"86",x"cc",x"87",x"c6"),
   380 => (x"6c",x"87",x"da",x"c0"),
   381 => (x"72",x"1e",x"71",x"49"),
   382 => (x"74",x"48",x"71",x"1e"),
   383 => (x"a1",x"f0",x"c0",x"49"),
   384 => (x"71",x"41",x"20",x"4a"),
   385 => (x"f8",x"ff",x"05",x"aa"),
   386 => (x"26",x"4a",x"26",x"87"),
   387 => (x"48",x"a6",x"dc",x"49"),
   388 => (x"c1",x"50",x"c1",x"c1"),
   389 => (x"bf",x"97",x"cc",x"d0"),
   390 => (x"b7",x"c1",x"c1",x"49"),
   391 => (x"dc",x"c1",x"04",x"a9"),
   392 => (x"66",x"97",x"dc",x"87"),
   393 => (x"1e",x"c3",x"c1",x"4b"),
   394 => (x"f4",x"c0",x"49",x"73"),
   395 => (x"86",x"c4",x"87",x"dd"),
   396 => (x"05",x"a8",x"66",x"d0"),
   397 => (x"d4",x"87",x"f5",x"c0"),
   398 => (x"49",x"c0",x"1e",x"66"),
   399 => (x"87",x"d3",x"f0",x"c0"),
   400 => (x"e9",x"c0",x"86",x"c4"),
   401 => (x"f2",x"c3",x"48",x"ec"),
   402 => (x"41",x"20",x"49",x"c0"),
   403 => (x"41",x"20",x"41",x"20"),
   404 => (x"41",x"20",x"41",x"20"),
   405 => (x"41",x"20",x"41",x"20"),
   406 => (x"51",x"10",x"51",x"10"),
   407 => (x"e0",x"c0",x"51",x"10"),
   408 => (x"66",x"c4",x"48",x"a6"),
   409 => (x"c0",x"d0",x"c1",x"78"),
   410 => (x"78",x"66",x"c4",x"48"),
   411 => (x"4a",x"73",x"83",x"c1"),
   412 => (x"97",x"cc",x"d0",x"c1"),
   413 => (x"b7",x"71",x"49",x"bf"),
   414 => (x"e8",x"fe",x"06",x"aa"),
   415 => (x"66",x"e0",x"c0",x"87"),
   416 => (x"90",x"66",x"d8",x"48"),
   417 => (x"58",x"a6",x"e4",x"c0"),
   418 => (x"1e",x"72",x"1e",x"71"),
   419 => (x"49",x"66",x"e8",x"c0"),
   420 => (x"f4",x"4a",x"66",x"d0"),
   421 => (x"4a",x"26",x"87",x"cb"),
   422 => (x"a6",x"dc",x"49",x"26"),
   423 => (x"66",x"e0",x"c0",x"58"),
   424 => (x"89",x"66",x"c8",x"49"),
   425 => (x"48",x"71",x"91",x"c7"),
   426 => (x"c0",x"88",x"66",x"d8"),
   427 => (x"6e",x"58",x"a6",x"e4"),
   428 => (x"82",x"ca",x"4a",x"bf"),
   429 => (x"97",x"c8",x"d0",x"c1"),
   430 => (x"c1",x"c1",x"49",x"bf"),
   431 => (x"cd",x"c0",x"05",x"a9"),
   432 => (x"72",x"8a",x"c1",x"87"),
   433 => (x"c0",x"d0",x"c1",x"48"),
   434 => (x"08",x"6e",x"88",x"bf"),
   435 => (x"66",x"c4",x"08",x"78"),
   436 => (x"c8",x"80",x"c1",x"48"),
   437 => (x"66",x"c4",x"58",x"a6"),
   438 => (x"c4",x"e8",x"c0",x"48"),
   439 => (x"06",x"a8",x"b7",x"bf"),
   440 => (x"c3",x"87",x"d9",x"f7"),
   441 => (x"ff",x"48",x"ec",x"ef"),
   442 => (x"c0",x"78",x"bf",x"c8"),
   443 => (x"f0",x"1e",x"c4",x"f1"),
   444 => (x"f1",x"c0",x"87",x"fc"),
   445 => (x"f5",x"f0",x"1e",x"d4"),
   446 => (x"d8",x"f1",x"c0",x"87"),
   447 => (x"87",x"ee",x"f0",x"1e"),
   448 => (x"1e",x"d0",x"f2",x"c0"),
   449 => (x"c1",x"87",x"e7",x"f0"),
   450 => (x"1e",x"bf",x"c0",x"d0"),
   451 => (x"1e",x"d4",x"f2",x"c0"),
   452 => (x"c5",x"87",x"db",x"f0"),
   453 => (x"f0",x"f2",x"c0",x"1e"),
   454 => (x"87",x"d2",x"f0",x"1e"),
   455 => (x"bf",x"c4",x"d0",x"c1"),
   456 => (x"cc",x"f3",x"c0",x"1e"),
   457 => (x"87",x"c6",x"f0",x"1e"),
   458 => (x"f3",x"c0",x"1e",x"c1"),
   459 => (x"fd",x"ef",x"1e",x"e8"),
   460 => (x"c8",x"d0",x"c1",x"87"),
   461 => (x"71",x"49",x"bf",x"97"),
   462 => (x"c4",x"f4",x"c0",x"1e"),
   463 => (x"87",x"ee",x"ef",x"1e"),
   464 => (x"c0",x"1e",x"c1",x"c1"),
   465 => (x"ef",x"1e",x"e0",x"f4"),
   466 => (x"d0",x"c1",x"87",x"e4"),
   467 => (x"49",x"bf",x"97",x"cc"),
   468 => (x"f4",x"c0",x"1e",x"71"),
   469 => (x"d5",x"ef",x"1e",x"fc"),
   470 => (x"1e",x"c2",x"c1",x"87"),
   471 => (x"1e",x"d8",x"f5",x"c0"),
   472 => (x"c1",x"87",x"cb",x"ef"),
   473 => (x"1e",x"bf",x"f0",x"d0"),
   474 => (x"1e",x"f4",x"f5",x"c0"),
   475 => (x"c7",x"87",x"ff",x"ee"),
   476 => (x"d0",x"f6",x"c0",x"1e"),
   477 => (x"87",x"f6",x"ee",x"1e"),
   478 => (x"bf",x"f4",x"ec",x"c1"),
   479 => (x"ec",x"f6",x"c0",x"1e"),
   480 => (x"87",x"ea",x"ee",x"1e"),
   481 => (x"1e",x"c8",x"f7",x"c0"),
   482 => (x"c0",x"87",x"e3",x"ee"),
   483 => (x"ee",x"1e",x"f4",x"f7"),
   484 => (x"cf",x"c1",x"87",x"dc"),
   485 => (x"1e",x"bf",x"bf",x"f8"),
   486 => (x"1e",x"c0",x"f8",x"c0"),
   487 => (x"c0",x"87",x"cf",x"ee"),
   488 => (x"ee",x"1e",x"dc",x"f8"),
   489 => (x"cf",x"c1",x"87",x"c8"),
   490 => (x"c4",x"49",x"bf",x"f8"),
   491 => (x"c0",x"1e",x"69",x"81"),
   492 => (x"ed",x"1e",x"d0",x"f9"),
   493 => (x"1e",x"c0",x"87",x"f8"),
   494 => (x"1e",x"ec",x"f9",x"c0"),
   495 => (x"c1",x"87",x"ef",x"ed"),
   496 => (x"49",x"bf",x"f8",x"cf"),
   497 => (x"1e",x"69",x"81",x"c8"),
   498 => (x"1e",x"c8",x"fa",x"c0"),
   499 => (x"c2",x"87",x"df",x"ed"),
   500 => (x"e4",x"fa",x"c0",x"1e"),
   501 => (x"87",x"d6",x"ed",x"1e"),
   502 => (x"bf",x"f8",x"cf",x"c1"),
   503 => (x"69",x"81",x"cc",x"49"),
   504 => (x"c0",x"fb",x"c0",x"1e"),
   505 => (x"87",x"c6",x"ed",x"1e"),
   506 => (x"fb",x"c0",x"1e",x"d1"),
   507 => (x"fd",x"ec",x"1e",x"dc"),
   508 => (x"f8",x"cf",x"c1",x"87"),
   509 => (x"81",x"d0",x"49",x"bf"),
   510 => (x"fb",x"c0",x"1e",x"71"),
   511 => (x"ed",x"ec",x"1e",x"f8"),
   512 => (x"d4",x"fc",x"c0",x"87"),
   513 => (x"87",x"e6",x"ec",x"1e"),
   514 => (x"1e",x"cc",x"fd",x"c0"),
   515 => (x"c1",x"87",x"df",x"ec"),
   516 => (x"bf",x"bf",x"fc",x"cf"),
   517 => (x"e0",x"fd",x"c0",x"1e"),
   518 => (x"87",x"d2",x"ec",x"1e"),
   519 => (x"1e",x"fc",x"fd",x"c0"),
   520 => (x"c1",x"87",x"cb",x"ec"),
   521 => (x"49",x"bf",x"fc",x"cf"),
   522 => (x"1e",x"69",x"81",x"c4"),
   523 => (x"1e",x"fc",x"fe",x"c0"),
   524 => (x"c0",x"87",x"fb",x"eb"),
   525 => (x"d8",x"ff",x"c0",x"1e"),
   526 => (x"87",x"f2",x"eb",x"1e"),
   527 => (x"bf",x"fc",x"cf",x"c1"),
   528 => (x"69",x"81",x"c8",x"49"),
   529 => (x"f4",x"ff",x"c0",x"1e"),
   530 => (x"87",x"e2",x"eb",x"1e"),
   531 => (x"c0",x"c1",x"1e",x"c1"),
   532 => (x"d9",x"eb",x"1e",x"d0"),
   533 => (x"fc",x"cf",x"c1",x"87"),
   534 => (x"81",x"cc",x"49",x"bf"),
   535 => (x"c0",x"c1",x"1e",x"69"),
   536 => (x"c9",x"eb",x"1e",x"ec"),
   537 => (x"c1",x"1e",x"d2",x"87"),
   538 => (x"eb",x"1e",x"c8",x"c1"),
   539 => (x"cf",x"c1",x"87",x"c0"),
   540 => (x"d0",x"49",x"bf",x"fc"),
   541 => (x"c1",x"1e",x"71",x"81"),
   542 => (x"ea",x"1e",x"e4",x"c1"),
   543 => (x"c2",x"c1",x"87",x"f0"),
   544 => (x"e9",x"ea",x"1e",x"c0"),
   545 => (x"66",x"dc",x"c4",x"87"),
   546 => (x"f8",x"c2",x"c1",x"1e"),
   547 => (x"87",x"de",x"ea",x"1e"),
   548 => (x"c3",x"c1",x"1e",x"c5"),
   549 => (x"d5",x"ea",x"1e",x"d4"),
   550 => (x"66",x"f4",x"c4",x"87"),
   551 => (x"f0",x"c3",x"c1",x"1e"),
   552 => (x"87",x"ca",x"ea",x"1e"),
   553 => (x"c4",x"c1",x"1e",x"cd"),
   554 => (x"c1",x"ea",x"1e",x"cc"),
   555 => (x"66",x"ec",x"c4",x"87"),
   556 => (x"e8",x"c4",x"c1",x"1e"),
   557 => (x"87",x"f6",x"e9",x"1e"),
   558 => (x"c5",x"c1",x"1e",x"c7"),
   559 => (x"ed",x"e9",x"1e",x"c4"),
   560 => (x"66",x"c4",x"c5",x"87"),
   561 => (x"e0",x"c5",x"c1",x"1e"),
   562 => (x"87",x"e2",x"e9",x"1e"),
   563 => (x"c5",x"c1",x"1e",x"c1"),
   564 => (x"d9",x"e9",x"1e",x"fc"),
   565 => (x"e0",x"f1",x"c3",x"87"),
   566 => (x"d8",x"c6",x"c1",x"1e"),
   567 => (x"87",x"ce",x"e9",x"1e"),
   568 => (x"1e",x"f4",x"c6",x"c1"),
   569 => (x"c3",x"87",x"c7",x"e9"),
   570 => (x"c1",x"1e",x"c0",x"f2"),
   571 => (x"e8",x"1e",x"ec",x"c7"),
   572 => (x"c8",x"c1",x"87",x"fc"),
   573 => (x"f5",x"e8",x"1e",x"c8"),
   574 => (x"c0",x"c9",x"c1",x"87"),
   575 => (x"87",x"ee",x"e8",x"1e"),
   576 => (x"bf",x"ec",x"ef",x"c3"),
   577 => (x"e8",x"ef",x"c3",x"49"),
   578 => (x"ef",x"c3",x"89",x"bf"),
   579 => (x"1e",x"71",x"59",x"f4"),
   580 => (x"1e",x"c4",x"c9",x"c1"),
   581 => (x"c5",x"87",x"d7",x"e8"),
   582 => (x"ef",x"c3",x"86",x"e8"),
   583 => (x"c1",x"48",x"bf",x"f0"),
   584 => (x"03",x"a8",x"b7",x"f8"),
   585 => (x"c0",x"87",x"d7",x"c0"),
   586 => (x"e8",x"1e",x"ec",x"ea"),
   587 => (x"eb",x"c0",x"87",x"c0"),
   588 => (x"f9",x"e7",x"1e",x"e4"),
   589 => (x"c4",x"ec",x"c0",x"87"),
   590 => (x"87",x"f2",x"e7",x"1e"),
   591 => (x"ef",x"c3",x"86",x"cc"),
   592 => (x"71",x"49",x"bf",x"f0"),
   593 => (x"92",x"e8",x"cf",x"4a"),
   594 => (x"1e",x"72",x"1e",x"71"),
   595 => (x"e8",x"c0",x"49",x"72"),
   596 => (x"e9",x"4a",x"bf",x"c4"),
   597 => (x"4a",x"26",x"87",x"cb"),
   598 => (x"ef",x"c3",x"49",x"26"),
   599 => (x"e8",x"c0",x"58",x"f8"),
   600 => (x"72",x"4a",x"bf",x"c4"),
   601 => (x"93",x"e8",x"cf",x"4b"),
   602 => (x"1e",x"72",x"1e",x"71"),
   603 => (x"e8",x"4a",x"09",x"73"),
   604 => (x"4a",x"26",x"87",x"ef"),
   605 => (x"ef",x"c3",x"49",x"26"),
   606 => (x"f9",x"c8",x"58",x"fc"),
   607 => (x"72",x"1e",x"71",x"92"),
   608 => (x"4a",x"09",x"72",x"1e"),
   609 => (x"26",x"87",x"da",x"e8"),
   610 => (x"c3",x"49",x"26",x"4a"),
   611 => (x"c0",x"58",x"c0",x"f0"),
   612 => (x"e6",x"1e",x"c8",x"ec"),
   613 => (x"ef",x"c3",x"87",x"d8"),
   614 => (x"c0",x"1e",x"bf",x"f4"),
   615 => (x"e6",x"1e",x"f8",x"ec"),
   616 => (x"ed",x"c0",x"87",x"cc"),
   617 => (x"c5",x"e6",x"1e",x"c0"),
   618 => (x"f8",x"ef",x"c3",x"87"),
   619 => (x"ed",x"c0",x"1e",x"bf"),
   620 => (x"f9",x"e5",x"1e",x"f0"),
   621 => (x"fc",x"ef",x"c3",x"87"),
   622 => (x"ed",x"c0",x"1e",x"bf"),
   623 => (x"ed",x"e5",x"1e",x"f8"),
   624 => (x"d8",x"ee",x"c0",x"87"),
   625 => (x"87",x"e6",x"e5",x"1e"),
   626 => (x"f8",x"fe",x"48",x"c0"),
   627 => (x"26",x"4d",x"26",x"8e"),
   628 => (x"26",x"4b",x"26",x"4c"),
   629 => (x"4a",x"71",x"1e",x"4f"),
   630 => (x"bf",x"f8",x"cf",x"c1"),
   631 => (x"c1",x"87",x"c6",x"02"),
   632 => (x"bf",x"bf",x"f8",x"cf"),
   633 => (x"f8",x"cf",x"c1",x"7a"),
   634 => (x"81",x"cc",x"49",x"bf"),
   635 => (x"d0",x"c1",x"1e",x"71"),
   636 => (x"ca",x"1e",x"bf",x"c0"),
   637 => (x"fb",x"e2",x"c0",x"49"),
   638 => (x"26",x"8e",x"f8",x"87"),
   639 => (x"00",x"00",x"00",x"4f"),
   640 => (x"00",x"00",x"00",x"00"),
   641 => (x"00",x"00",x"61",x"a8"),
   642 => (x"67",x"6f",x"72",x"50"),
   643 => (x"20",x"6d",x"61",x"72"),
   644 => (x"70",x"6d",x"6f",x"63"),
   645 => (x"64",x"65",x"6c",x"69"),
   646 => (x"74",x"69",x"77",x"20"),
   647 => (x"72",x"27",x"20",x"68"),
   648 => (x"73",x"69",x"67",x"65"),
   649 => (x"27",x"72",x"65",x"74"),
   650 => (x"74",x"74",x"61",x"20"),
   651 => (x"75",x"62",x"69",x"72"),
   652 => (x"00",x"0a",x"65",x"74"),
   653 => (x"00",x"00",x"00",x"0a"),
   654 => (x"67",x"6f",x"72",x"50"),
   655 => (x"20",x"6d",x"61",x"72"),
   656 => (x"70",x"6d",x"6f",x"63"),
   657 => (x"64",x"65",x"6c",x"69"),
   658 => (x"74",x"69",x"77",x"20"),
   659 => (x"74",x"75",x"6f",x"68"),
   660 => (x"65",x"72",x"27",x"20"),
   661 => (x"74",x"73",x"69",x"67"),
   662 => (x"20",x"27",x"72",x"65"),
   663 => (x"72",x"74",x"74",x"61"),
   664 => (x"74",x"75",x"62",x"69"),
   665 => (x"00",x"00",x"0a",x"65"),
   666 => (x"00",x"00",x"00",x"0a"),
   667 => (x"59",x"52",x"48",x"44"),
   668 => (x"4e",x"4f",x"54",x"53"),
   669 => (x"52",x"50",x"20",x"45"),
   670 => (x"41",x"52",x"47",x"4f"),
   671 => (x"33",x"20",x"2c",x"4d"),
   672 => (x"20",x"44",x"52",x"27"),
   673 => (x"49",x"52",x"54",x"53"),
   674 => (x"00",x"00",x"47",x"4e"),
   675 => (x"59",x"52",x"48",x"44"),
   676 => (x"4e",x"4f",x"54",x"53"),
   677 => (x"52",x"50",x"20",x"45"),
   678 => (x"41",x"52",x"47",x"4f"),
   679 => (x"32",x"20",x"2c",x"4d"),
   680 => (x"20",x"44",x"4e",x"27"),
   681 => (x"49",x"52",x"54",x"53"),
   682 => (x"00",x"00",x"47",x"4e"),
   683 => (x"73",x"61",x"65",x"4d"),
   684 => (x"64",x"65",x"72",x"75"),
   685 => (x"6d",x"69",x"74",x"20"),
   686 => (x"6f",x"74",x"20",x"65"),
   687 => (x"6d",x"73",x"20",x"6f"),
   688 => (x"20",x"6c",x"6c",x"61"),
   689 => (x"6f",x"20",x"6f",x"74"),
   690 => (x"69",x"61",x"74",x"62"),
   691 => (x"65",x"6d",x"20",x"6e"),
   692 => (x"6e",x"69",x"6e",x"61"),
   693 => (x"6c",x"75",x"66",x"67"),
   694 => (x"73",x"65",x"72",x"20"),
   695 => (x"73",x"74",x"6c",x"75"),
   696 => (x"00",x"00",x"00",x"0a"),
   697 => (x"61",x"65",x"6c",x"50"),
   698 => (x"69",x"20",x"65",x"73"),
   699 => (x"65",x"72",x"63",x"6e"),
   700 => (x"20",x"65",x"73",x"61"),
   701 => (x"62",x"6d",x"75",x"6e"),
   702 => (x"6f",x"20",x"72",x"65"),
   703 => (x"75",x"72",x"20",x"66"),
   704 => (x"00",x"0a",x"73",x"6e"),
   705 => (x"00",x"00",x"00",x"0a"),
   706 => (x"72",x"63",x"69",x"4d"),
   707 => (x"63",x"65",x"73",x"6f"),
   708 => (x"73",x"64",x"6e",x"6f"),
   709 => (x"72",x"6f",x"66",x"20"),
   710 => (x"65",x"6e",x"6f",x"20"),
   711 => (x"6e",x"75",x"72",x"20"),
   712 => (x"72",x"68",x"74",x"20"),
   713 => (x"68",x"67",x"75",x"6f"),
   714 => (x"72",x"68",x"44",x"20"),
   715 => (x"6f",x"74",x"73",x"79"),
   716 => (x"20",x"3a",x"65",x"6e"),
   717 => (x"00",x"00",x"00",x"00"),
   718 => (x"0a",x"20",x"64",x"25"),
   719 => (x"00",x"00",x"00",x"00"),
   720 => (x"79",x"72",x"68",x"44"),
   721 => (x"6e",x"6f",x"74",x"73"),
   722 => (x"70",x"20",x"73",x"65"),
   723 => (x"53",x"20",x"72",x"65"),
   724 => (x"6e",x"6f",x"63",x"65"),
   725 => (x"20",x"20",x"3a",x"64"),
   726 => (x"20",x"20",x"20",x"20"),
   727 => (x"20",x"20",x"20",x"20"),
   728 => (x"20",x"20",x"20",x"20"),
   729 => (x"20",x"20",x"20",x"20"),
   730 => (x"20",x"20",x"20",x"20"),
   731 => (x"00",x"00",x"00",x"00"),
   732 => (x"0a",x"20",x"64",x"25"),
   733 => (x"00",x"00",x"00",x"00"),
   734 => (x"20",x"58",x"41",x"56"),
   735 => (x"53",x"50",x"49",x"4d"),
   736 => (x"74",x"61",x"72",x"20"),
   737 => (x"20",x"67",x"6e",x"69"),
   738 => (x"30",x"31",x"20",x"2a"),
   739 => (x"3d",x"20",x"30",x"30"),
   740 => (x"20",x"64",x"25",x"20"),
   741 => (x"00",x"00",x"00",x"0a"),
   742 => (x"00",x"00",x"00",x"0a"),
   743 => (x"59",x"52",x"48",x"44"),
   744 => (x"4e",x"4f",x"54",x"53"),
   745 => (x"52",x"50",x"20",x"45"),
   746 => (x"41",x"52",x"47",x"4f"),
   747 => (x"53",x"20",x"2c",x"4d"),
   748 => (x"20",x"45",x"4d",x"4f"),
   749 => (x"49",x"52",x"54",x"53"),
   750 => (x"00",x"00",x"47",x"4e"),
   751 => (x"59",x"52",x"48",x"44"),
   752 => (x"4e",x"4f",x"54",x"53"),
   753 => (x"52",x"50",x"20",x"45"),
   754 => (x"41",x"52",x"47",x"4f"),
   755 => (x"31",x"20",x"2c",x"4d"),
   756 => (x"20",x"54",x"53",x"27"),
   757 => (x"49",x"52",x"54",x"53"),
   758 => (x"00",x"00",x"47",x"4e"),
   759 => (x"00",x"00",x"00",x"0a"),
   760 => (x"79",x"72",x"68",x"44"),
   761 => (x"6e",x"6f",x"74",x"73"),
   762 => (x"65",x"42",x"20",x"65"),
   763 => (x"6d",x"68",x"63",x"6e"),
   764 => (x"2c",x"6b",x"72",x"61"),
   765 => (x"72",x"65",x"56",x"20"),
   766 => (x"6e",x"6f",x"69",x"73"),
   767 => (x"31",x"2e",x"32",x"20"),
   768 => (x"61",x"4c",x"28",x"20"),
   769 => (x"61",x"75",x"67",x"6e"),
   770 => (x"20",x"3a",x"65",x"67"),
   771 => (x"00",x"0a",x"29",x"43"),
   772 => (x"00",x"00",x"00",x"0a"),
   773 => (x"63",x"65",x"78",x"45"),
   774 => (x"6f",x"69",x"74",x"75"),
   775 => (x"74",x"73",x"20",x"6e"),
   776 => (x"73",x"74",x"72",x"61"),
   777 => (x"64",x"25",x"20",x"2c"),
   778 => (x"6e",x"75",x"72",x"20"),
   779 => (x"68",x"74",x"20",x"73"),
   780 => (x"67",x"75",x"6f",x"72"),
   781 => (x"68",x"44",x"20",x"68"),
   782 => (x"74",x"73",x"79",x"72"),
   783 => (x"0a",x"65",x"6e",x"6f"),
   784 => (x"00",x"00",x"00",x"00"),
   785 => (x"63",x"65",x"78",x"45"),
   786 => (x"6f",x"69",x"74",x"75"),
   787 => (x"6e",x"65",x"20",x"6e"),
   788 => (x"00",x"0a",x"73",x"64"),
   789 => (x"00",x"00",x"00",x"0a"),
   790 => (x"61",x"6e",x"69",x"46"),
   791 => (x"61",x"76",x"20",x"6c"),
   792 => (x"73",x"65",x"75",x"6c"),
   793 => (x"20",x"66",x"6f",x"20"),
   794 => (x"20",x"65",x"68",x"74"),
   795 => (x"69",x"72",x"61",x"76"),
   796 => (x"65",x"6c",x"62",x"61"),
   797 => (x"73",x"75",x"20",x"73"),
   798 => (x"69",x"20",x"64",x"65"),
   799 => (x"68",x"74",x"20",x"6e"),
   800 => (x"65",x"62",x"20",x"65"),
   801 => (x"6d",x"68",x"63",x"6e"),
   802 => (x"3a",x"6b",x"72",x"61"),
   803 => (x"00",x"00",x"00",x"0a"),
   804 => (x"00",x"00",x"00",x"0a"),
   805 => (x"5f",x"74",x"6e",x"49"),
   806 => (x"62",x"6f",x"6c",x"47"),
   807 => (x"20",x"20",x"20",x"3a"),
   808 => (x"20",x"20",x"20",x"20"),
   809 => (x"20",x"20",x"20",x"20"),
   810 => (x"0a",x"64",x"25",x"20"),
   811 => (x"00",x"00",x"00",x"00"),
   812 => (x"20",x"20",x"20",x"20"),
   813 => (x"20",x"20",x"20",x"20"),
   814 => (x"75",x"6f",x"68",x"73"),
   815 => (x"62",x"20",x"64",x"6c"),
   816 => (x"20",x"20",x"3a",x"65"),
   817 => (x"0a",x"64",x"25",x"20"),
   818 => (x"00",x"00",x"00",x"00"),
   819 => (x"6c",x"6f",x"6f",x"42"),
   820 => (x"6f",x"6c",x"47",x"5f"),
   821 => (x"20",x"20",x"3a",x"62"),
   822 => (x"20",x"20",x"20",x"20"),
   823 => (x"20",x"20",x"20",x"20"),
   824 => (x"0a",x"64",x"25",x"20"),
   825 => (x"00",x"00",x"00",x"00"),
   826 => (x"20",x"20",x"20",x"20"),
   827 => (x"20",x"20",x"20",x"20"),
   828 => (x"75",x"6f",x"68",x"73"),
   829 => (x"62",x"20",x"64",x"6c"),
   830 => (x"20",x"20",x"3a",x"65"),
   831 => (x"0a",x"64",x"25",x"20"),
   832 => (x"00",x"00",x"00",x"00"),
   833 => (x"31",x"5f",x"68",x"43"),
   834 => (x"6f",x"6c",x"47",x"5f"),
   835 => (x"20",x"20",x"3a",x"62"),
   836 => (x"20",x"20",x"20",x"20"),
   837 => (x"20",x"20",x"20",x"20"),
   838 => (x"0a",x"63",x"25",x"20"),
   839 => (x"00",x"00",x"00",x"00"),
   840 => (x"20",x"20",x"20",x"20"),
   841 => (x"20",x"20",x"20",x"20"),
   842 => (x"75",x"6f",x"68",x"73"),
   843 => (x"62",x"20",x"64",x"6c"),
   844 => (x"20",x"20",x"3a",x"65"),
   845 => (x"0a",x"63",x"25",x"20"),
   846 => (x"00",x"00",x"00",x"00"),
   847 => (x"32",x"5f",x"68",x"43"),
   848 => (x"6f",x"6c",x"47",x"5f"),
   849 => (x"20",x"20",x"3a",x"62"),
   850 => (x"20",x"20",x"20",x"20"),
   851 => (x"20",x"20",x"20",x"20"),
   852 => (x"0a",x"63",x"25",x"20"),
   853 => (x"00",x"00",x"00",x"00"),
   854 => (x"20",x"20",x"20",x"20"),
   855 => (x"20",x"20",x"20",x"20"),
   856 => (x"75",x"6f",x"68",x"73"),
   857 => (x"62",x"20",x"64",x"6c"),
   858 => (x"20",x"20",x"3a",x"65"),
   859 => (x"0a",x"63",x"25",x"20"),
   860 => (x"00",x"00",x"00",x"00"),
   861 => (x"5f",x"72",x"72",x"41"),
   862 => (x"6c",x"47",x"5f",x"31"),
   863 => (x"38",x"5b",x"62",x"6f"),
   864 => (x"20",x"20",x"3a",x"5d"),
   865 => (x"20",x"20",x"20",x"20"),
   866 => (x"0a",x"64",x"25",x"20"),
   867 => (x"00",x"00",x"00",x"00"),
   868 => (x"20",x"20",x"20",x"20"),
   869 => (x"20",x"20",x"20",x"20"),
   870 => (x"75",x"6f",x"68",x"73"),
   871 => (x"62",x"20",x"64",x"6c"),
   872 => (x"20",x"20",x"3a",x"65"),
   873 => (x"0a",x"64",x"25",x"20"),
   874 => (x"00",x"00",x"00",x"00"),
   875 => (x"5f",x"72",x"72",x"41"),
   876 => (x"6c",x"47",x"5f",x"32"),
   877 => (x"38",x"5b",x"62",x"6f"),
   878 => (x"5d",x"37",x"5b",x"5d"),
   879 => (x"20",x"20",x"20",x"3a"),
   880 => (x"0a",x"64",x"25",x"20"),
   881 => (x"00",x"00",x"00",x"00"),
   882 => (x"20",x"20",x"20",x"20"),
   883 => (x"20",x"20",x"20",x"20"),
   884 => (x"75",x"6f",x"68",x"73"),
   885 => (x"62",x"20",x"64",x"6c"),
   886 => (x"20",x"20",x"3a",x"65"),
   887 => (x"6d",x"75",x"4e",x"20"),
   888 => (x"5f",x"72",x"65",x"62"),
   889 => (x"52",x"5f",x"66",x"4f"),
   890 => (x"20",x"73",x"6e",x"75"),
   891 => (x"30",x"31",x"20",x"2b"),
   892 => (x"00",x"00",x"00",x"0a"),
   893 => (x"5f",x"72",x"74",x"50"),
   894 => (x"62",x"6f",x"6c",x"47"),
   895 => (x"00",x"0a",x"3e",x"2d"),
   896 => (x"74",x"50",x"20",x"20"),
   897 => (x"6f",x"43",x"5f",x"72"),
   898 => (x"20",x"3a",x"70",x"6d"),
   899 => (x"20",x"20",x"20",x"20"),
   900 => (x"20",x"20",x"20",x"20"),
   901 => (x"0a",x"64",x"25",x"20"),
   902 => (x"00",x"00",x"00",x"00"),
   903 => (x"20",x"20",x"20",x"20"),
   904 => (x"20",x"20",x"20",x"20"),
   905 => (x"75",x"6f",x"68",x"73"),
   906 => (x"62",x"20",x"64",x"6c"),
   907 => (x"20",x"20",x"3a",x"65"),
   908 => (x"6d",x"69",x"28",x"20"),
   909 => (x"6d",x"65",x"6c",x"70"),
   910 => (x"61",x"74",x"6e",x"65"),
   911 => (x"6e",x"6f",x"69",x"74"),
   912 => (x"70",x"65",x"64",x"2d"),
   913 => (x"65",x"64",x"6e",x"65"),
   914 => (x"0a",x"29",x"74",x"6e"),
   915 => (x"00",x"00",x"00",x"00"),
   916 => (x"69",x"44",x"20",x"20"),
   917 => (x"3a",x"72",x"63",x"73"),
   918 => (x"20",x"20",x"20",x"20"),
   919 => (x"20",x"20",x"20",x"20"),
   920 => (x"20",x"20",x"20",x"20"),
   921 => (x"0a",x"64",x"25",x"20"),
   922 => (x"00",x"00",x"00",x"00"),
   923 => (x"20",x"20",x"20",x"20"),
   924 => (x"20",x"20",x"20",x"20"),
   925 => (x"75",x"6f",x"68",x"73"),
   926 => (x"62",x"20",x"64",x"6c"),
   927 => (x"20",x"20",x"3a",x"65"),
   928 => (x"0a",x"64",x"25",x"20"),
   929 => (x"00",x"00",x"00",x"00"),
   930 => (x"6e",x"45",x"20",x"20"),
   931 => (x"43",x"5f",x"6d",x"75"),
   932 => (x"3a",x"70",x"6d",x"6f"),
   933 => (x"20",x"20",x"20",x"20"),
   934 => (x"20",x"20",x"20",x"20"),
   935 => (x"0a",x"64",x"25",x"20"),
   936 => (x"00",x"00",x"00",x"00"),
   937 => (x"20",x"20",x"20",x"20"),
   938 => (x"20",x"20",x"20",x"20"),
   939 => (x"75",x"6f",x"68",x"73"),
   940 => (x"62",x"20",x"64",x"6c"),
   941 => (x"20",x"20",x"3a",x"65"),
   942 => (x"0a",x"64",x"25",x"20"),
   943 => (x"00",x"00",x"00",x"00"),
   944 => (x"6e",x"49",x"20",x"20"),
   945 => (x"6f",x"43",x"5f",x"74"),
   946 => (x"20",x"3a",x"70",x"6d"),
   947 => (x"20",x"20",x"20",x"20"),
   948 => (x"20",x"20",x"20",x"20"),
   949 => (x"0a",x"64",x"25",x"20"),
   950 => (x"00",x"00",x"00",x"00"),
   951 => (x"20",x"20",x"20",x"20"),
   952 => (x"20",x"20",x"20",x"20"),
   953 => (x"75",x"6f",x"68",x"73"),
   954 => (x"62",x"20",x"64",x"6c"),
   955 => (x"20",x"20",x"3a",x"65"),
   956 => (x"0a",x"64",x"25",x"20"),
   957 => (x"00",x"00",x"00",x"00"),
   958 => (x"74",x"53",x"20",x"20"),
   959 => (x"6f",x"43",x"5f",x"72"),
   960 => (x"20",x"3a",x"70",x"6d"),
   961 => (x"20",x"20",x"20",x"20"),
   962 => (x"20",x"20",x"20",x"20"),
   963 => (x"0a",x"73",x"25",x"20"),
   964 => (x"00",x"00",x"00",x"00"),
   965 => (x"20",x"20",x"20",x"20"),
   966 => (x"20",x"20",x"20",x"20"),
   967 => (x"75",x"6f",x"68",x"73"),
   968 => (x"62",x"20",x"64",x"6c"),
   969 => (x"20",x"20",x"3a",x"65"),
   970 => (x"52",x"48",x"44",x"20"),
   971 => (x"4f",x"54",x"53",x"59"),
   972 => (x"50",x"20",x"45",x"4e"),
   973 => (x"52",x"47",x"4f",x"52"),
   974 => (x"20",x"2c",x"4d",x"41"),
   975 => (x"45",x"4d",x"4f",x"53"),
   976 => (x"52",x"54",x"53",x"20"),
   977 => (x"0a",x"47",x"4e",x"49"),
   978 => (x"00",x"00",x"00",x"00"),
   979 => (x"74",x"78",x"65",x"4e"),
   980 => (x"72",x"74",x"50",x"5f"),
   981 => (x"6f",x"6c",x"47",x"5f"),
   982 => (x"0a",x"3e",x"2d",x"62"),
   983 => (x"00",x"00",x"00",x"00"),
   984 => (x"74",x"50",x"20",x"20"),
   985 => (x"6f",x"43",x"5f",x"72"),
   986 => (x"20",x"3a",x"70",x"6d"),
   987 => (x"20",x"20",x"20",x"20"),
   988 => (x"20",x"20",x"20",x"20"),
   989 => (x"0a",x"64",x"25",x"20"),
   990 => (x"00",x"00",x"00",x"00"),
   991 => (x"20",x"20",x"20",x"20"),
   992 => (x"20",x"20",x"20",x"20"),
   993 => (x"75",x"6f",x"68",x"73"),
   994 => (x"62",x"20",x"64",x"6c"),
   995 => (x"20",x"20",x"3a",x"65"),
   996 => (x"6d",x"69",x"28",x"20"),
   997 => (x"6d",x"65",x"6c",x"70"),
   998 => (x"61",x"74",x"6e",x"65"),
   999 => (x"6e",x"6f",x"69",x"74"),
  1000 => (x"70",x"65",x"64",x"2d"),
  1001 => (x"65",x"64",x"6e",x"65"),
  1002 => (x"2c",x"29",x"74",x"6e"),
  1003 => (x"6d",x"61",x"73",x"20"),
  1004 => (x"73",x"61",x"20",x"65"),
  1005 => (x"6f",x"62",x"61",x"20"),
  1006 => (x"00",x"0a",x"65",x"76"),
  1007 => (x"69",x"44",x"20",x"20"),
  1008 => (x"3a",x"72",x"63",x"73"),
  1009 => (x"20",x"20",x"20",x"20"),
  1010 => (x"20",x"20",x"20",x"20"),
  1011 => (x"20",x"20",x"20",x"20"),
  1012 => (x"0a",x"64",x"25",x"20"),
  1013 => (x"00",x"00",x"00",x"00"),
  1014 => (x"20",x"20",x"20",x"20"),
  1015 => (x"20",x"20",x"20",x"20"),
  1016 => (x"75",x"6f",x"68",x"73"),
  1017 => (x"62",x"20",x"64",x"6c"),
  1018 => (x"20",x"20",x"3a",x"65"),
  1019 => (x"0a",x"64",x"25",x"20"),
  1020 => (x"00",x"00",x"00",x"00"),
  1021 => (x"6e",x"45",x"20",x"20"),
  1022 => (x"43",x"5f",x"6d",x"75"),
  1023 => (x"3a",x"70",x"6d",x"6f"),
  1024 => (x"20",x"20",x"20",x"20"),
  1025 => (x"20",x"20",x"20",x"20"),
  1026 => (x"0a",x"64",x"25",x"20"),
  1027 => (x"00",x"00",x"00",x"00"),
  1028 => (x"20",x"20",x"20",x"20"),
  1029 => (x"20",x"20",x"20",x"20"),
  1030 => (x"75",x"6f",x"68",x"73"),
  1031 => (x"62",x"20",x"64",x"6c"),
  1032 => (x"20",x"20",x"3a",x"65"),
  1033 => (x"0a",x"64",x"25",x"20"),
  1034 => (x"00",x"00",x"00",x"00"),
  1035 => (x"6e",x"49",x"20",x"20"),
  1036 => (x"6f",x"43",x"5f",x"74"),
  1037 => (x"20",x"3a",x"70",x"6d"),
  1038 => (x"20",x"20",x"20",x"20"),
  1039 => (x"20",x"20",x"20",x"20"),
  1040 => (x"0a",x"64",x"25",x"20"),
  1041 => (x"00",x"00",x"00",x"00"),
  1042 => (x"20",x"20",x"20",x"20"),
  1043 => (x"20",x"20",x"20",x"20"),
  1044 => (x"75",x"6f",x"68",x"73"),
  1045 => (x"62",x"20",x"64",x"6c"),
  1046 => (x"20",x"20",x"3a",x"65"),
  1047 => (x"0a",x"64",x"25",x"20"),
  1048 => (x"00",x"00",x"00",x"00"),
  1049 => (x"74",x"53",x"20",x"20"),
  1050 => (x"6f",x"43",x"5f",x"72"),
  1051 => (x"20",x"3a",x"70",x"6d"),
  1052 => (x"20",x"20",x"20",x"20"),
  1053 => (x"20",x"20",x"20",x"20"),
  1054 => (x"0a",x"73",x"25",x"20"),
  1055 => (x"00",x"00",x"00",x"00"),
  1056 => (x"20",x"20",x"20",x"20"),
  1057 => (x"20",x"20",x"20",x"20"),
  1058 => (x"75",x"6f",x"68",x"73"),
  1059 => (x"62",x"20",x"64",x"6c"),
  1060 => (x"20",x"20",x"3a",x"65"),
  1061 => (x"52",x"48",x"44",x"20"),
  1062 => (x"4f",x"54",x"53",x"59"),
  1063 => (x"50",x"20",x"45",x"4e"),
  1064 => (x"52",x"47",x"4f",x"52"),
  1065 => (x"20",x"2c",x"4d",x"41"),
  1066 => (x"45",x"4d",x"4f",x"53"),
  1067 => (x"52",x"54",x"53",x"20"),
  1068 => (x"0a",x"47",x"4e",x"49"),
  1069 => (x"00",x"00",x"00",x"00"),
  1070 => (x"5f",x"74",x"6e",x"49"),
  1071 => (x"6f",x"4c",x"5f",x"31"),
  1072 => (x"20",x"20",x"3a",x"63"),
  1073 => (x"20",x"20",x"20",x"20"),
  1074 => (x"20",x"20",x"20",x"20"),
  1075 => (x"0a",x"64",x"25",x"20"),
  1076 => (x"00",x"00",x"00",x"00"),
  1077 => (x"20",x"20",x"20",x"20"),
  1078 => (x"20",x"20",x"20",x"20"),
  1079 => (x"75",x"6f",x"68",x"73"),
  1080 => (x"62",x"20",x"64",x"6c"),
  1081 => (x"20",x"20",x"3a",x"65"),
  1082 => (x"0a",x"64",x"25",x"20"),
  1083 => (x"00",x"00",x"00",x"00"),
  1084 => (x"5f",x"74",x"6e",x"49"),
  1085 => (x"6f",x"4c",x"5f",x"32"),
  1086 => (x"20",x"20",x"3a",x"63"),
  1087 => (x"20",x"20",x"20",x"20"),
  1088 => (x"20",x"20",x"20",x"20"),
  1089 => (x"0a",x"64",x"25",x"20"),
  1090 => (x"00",x"00",x"00",x"00"),
  1091 => (x"20",x"20",x"20",x"20"),
  1092 => (x"20",x"20",x"20",x"20"),
  1093 => (x"75",x"6f",x"68",x"73"),
  1094 => (x"62",x"20",x"64",x"6c"),
  1095 => (x"20",x"20",x"3a",x"65"),
  1096 => (x"0a",x"64",x"25",x"20"),
  1097 => (x"00",x"00",x"00",x"00"),
  1098 => (x"5f",x"74",x"6e",x"49"),
  1099 => (x"6f",x"4c",x"5f",x"33"),
  1100 => (x"20",x"20",x"3a",x"63"),
  1101 => (x"20",x"20",x"20",x"20"),
  1102 => (x"20",x"20",x"20",x"20"),
  1103 => (x"0a",x"64",x"25",x"20"),
  1104 => (x"00",x"00",x"00",x"00"),
  1105 => (x"20",x"20",x"20",x"20"),
  1106 => (x"20",x"20",x"20",x"20"),
  1107 => (x"75",x"6f",x"68",x"73"),
  1108 => (x"62",x"20",x"64",x"6c"),
  1109 => (x"20",x"20",x"3a",x"65"),
  1110 => (x"0a",x"64",x"25",x"20"),
  1111 => (x"00",x"00",x"00",x"00"),
  1112 => (x"6d",x"75",x"6e",x"45"),
  1113 => (x"63",x"6f",x"4c",x"5f"),
  1114 => (x"20",x"20",x"20",x"3a"),
  1115 => (x"20",x"20",x"20",x"20"),
  1116 => (x"20",x"20",x"20",x"20"),
  1117 => (x"0a",x"64",x"25",x"20"),
  1118 => (x"00",x"00",x"00",x"00"),
  1119 => (x"20",x"20",x"20",x"20"),
  1120 => (x"20",x"20",x"20",x"20"),
  1121 => (x"75",x"6f",x"68",x"73"),
  1122 => (x"62",x"20",x"64",x"6c"),
  1123 => (x"20",x"20",x"3a",x"65"),
  1124 => (x"0a",x"64",x"25",x"20"),
  1125 => (x"00",x"00",x"00",x"00"),
  1126 => (x"5f",x"72",x"74",x"53"),
  1127 => (x"6f",x"4c",x"5f",x"31"),
  1128 => (x"20",x"20",x"3a",x"63"),
  1129 => (x"20",x"20",x"20",x"20"),
  1130 => (x"20",x"20",x"20",x"20"),
  1131 => (x"0a",x"73",x"25",x"20"),
  1132 => (x"00",x"00",x"00",x"00"),
  1133 => (x"20",x"20",x"20",x"20"),
  1134 => (x"20",x"20",x"20",x"20"),
  1135 => (x"75",x"6f",x"68",x"73"),
  1136 => (x"62",x"20",x"64",x"6c"),
  1137 => (x"20",x"20",x"3a",x"65"),
  1138 => (x"52",x"48",x"44",x"20"),
  1139 => (x"4f",x"54",x"53",x"59"),
  1140 => (x"50",x"20",x"45",x"4e"),
  1141 => (x"52",x"47",x"4f",x"52"),
  1142 => (x"20",x"2c",x"4d",x"41"),
  1143 => (x"54",x"53",x"27",x"31"),
  1144 => (x"52",x"54",x"53",x"20"),
  1145 => (x"0a",x"47",x"4e",x"49"),
  1146 => (x"00",x"00",x"00",x"00"),
  1147 => (x"5f",x"72",x"74",x"53"),
  1148 => (x"6f",x"4c",x"5f",x"32"),
  1149 => (x"20",x"20",x"3a",x"63"),
  1150 => (x"20",x"20",x"20",x"20"),
  1151 => (x"20",x"20",x"20",x"20"),
  1152 => (x"0a",x"73",x"25",x"20"),
  1153 => (x"00",x"00",x"00",x"00"),
  1154 => (x"20",x"20",x"20",x"20"),
  1155 => (x"20",x"20",x"20",x"20"),
  1156 => (x"75",x"6f",x"68",x"73"),
  1157 => (x"62",x"20",x"64",x"6c"),
  1158 => (x"20",x"20",x"3a",x"65"),
  1159 => (x"52",x"48",x"44",x"20"),
  1160 => (x"4f",x"54",x"53",x"59"),
  1161 => (x"50",x"20",x"45",x"4e"),
  1162 => (x"52",x"47",x"4f",x"52"),
  1163 => (x"20",x"2c",x"4d",x"41"),
  1164 => (x"44",x"4e",x"27",x"32"),
  1165 => (x"52",x"54",x"53",x"20"),
  1166 => (x"0a",x"47",x"4e",x"49"),
  1167 => (x"00",x"00",x"00",x"00"),
  1168 => (x"00",x"00",x"00",x"0a"),
  1169 => (x"72",x"65",x"73",x"55"),
  1170 => (x"6d",x"69",x"74",x"20"),
  1171 => (x"25",x"20",x"3a",x"65"),
  1172 => (x"1e",x"00",x"0a",x"64"),
  1173 => (x"1e",x"74",x"1e",x"73"),
  1174 => (x"66",x"cc",x"4b",x"71"),
  1175 => (x"c2",x"7a",x"73",x"4a"),
  1176 => (x"87",x"c4",x"05",x"ab"),
  1177 => (x"87",x"c2",x"4c",x"c1"),
  1178 => (x"9c",x"74",x"4c",x"c0"),
  1179 => (x"c3",x"87",x"c2",x"05"),
  1180 => (x"02",x"9b",x"73",x"7a"),
  1181 => (x"49",x"73",x"87",x"da"),
  1182 => (x"d7",x"02",x"89",x"c1"),
  1183 => (x"02",x"89",x"c1",x"87"),
  1184 => (x"c1",x"87",x"e5",x"c0"),
  1185 => (x"e5",x"c0",x"02",x"89"),
  1186 => (x"02",x"89",x"c1",x"87"),
  1187 => (x"87",x"de",x"87",x"de"),
  1188 => (x"87",x"da",x"7a",x"c0"),
  1189 => (x"bf",x"c0",x"d0",x"c1"),
  1190 => (x"b7",x"e4",x"c1",x"48"),
  1191 => (x"87",x"c4",x"06",x"a8"),
  1192 => (x"87",x"ca",x"7a",x"c0"),
  1193 => (x"87",x"c6",x"7a",x"c3"),
  1194 => (x"87",x"c2",x"7a",x"c1"),
  1195 => (x"4c",x"26",x"7a",x"c2"),
  1196 => (x"4f",x"26",x"4b",x"26"),
  1197 => (x"72",x"4a",x"71",x"1e"),
  1198 => (x"c4",x"81",x"c2",x"49"),
  1199 => (x"80",x"71",x"48",x"66"),
  1200 => (x"78",x"08",x"66",x"c8"),
  1201 => (x"0e",x"4f",x"26",x"08"),
  1202 => (x"5d",x"5c",x"5b",x"5e"),
  1203 => (x"c4",x"86",x"f4",x"0e"),
  1204 => (x"e0",x"c0",x"59",x"a6"),
  1205 => (x"84",x"c5",x"4c",x"66"),
  1206 => (x"90",x"c4",x"48",x"74"),
  1207 => (x"6e",x"58",x"a6",x"c8"),
  1208 => (x"85",x"66",x"c4",x"4d"),
  1209 => (x"7d",x"66",x"e4",x"c0"),
  1210 => (x"c0",x"49",x"a5",x"c4"),
  1211 => (x"c1",x"79",x"66",x"e4"),
  1212 => (x"74",x"49",x"a5",x"f8"),
  1213 => (x"48",x"a6",x"c8",x"79"),
  1214 => (x"b7",x"78",x"a4",x"c1"),
  1215 => (x"87",x"dd",x"01",x"ac"),
  1216 => (x"c8",x"c3",x"49",x"74"),
  1217 => (x"4a",x"66",x"dc",x"91"),
  1218 => (x"66",x"c4",x"82",x"71"),
  1219 => (x"4b",x"66",x"c8",x"82"),
  1220 => (x"83",x"c1",x"8b",x"74"),
  1221 => (x"82",x"c4",x"7a",x"74"),
  1222 => (x"f7",x"01",x"8b",x"c1"),
  1223 => (x"c3",x"49",x"74",x"87"),
  1224 => (x"66",x"dc",x"91",x"c8"),
  1225 => (x"c4",x"4a",x"71",x"81"),
  1226 => (x"8a",x"c4",x"82",x"66"),
  1227 => (x"80",x"c1",x"48",x"6a"),
  1228 => (x"fe",x"c0",x"7a",x"70"),
  1229 => (x"66",x"c4",x"81",x"e0"),
  1230 => (x"c1",x"79",x"6d",x"81"),
  1231 => (x"c5",x"48",x"c0",x"d0"),
  1232 => (x"26",x"8e",x"f4",x"78"),
  1233 => (x"26",x"4c",x"26",x"4d"),
  1234 => (x"1e",x"4f",x"26",x"4b"),
  1235 => (x"1e",x"74",x"1e",x"73"),
  1236 => (x"4c",x"73",x"4b",x"71"),
  1237 => (x"66",x"cc",x"4a",x"74"),
  1238 => (x"aa",x"b7",x"71",x"49"),
  1239 => (x"c0",x"87",x"c4",x"02"),
  1240 => (x"c1",x"87",x"c7",x"48"),
  1241 => (x"5c",x"97",x"cc",x"d0"),
  1242 => (x"4c",x"26",x"48",x"c1"),
  1243 => (x"4f",x"26",x"4b",x"26"),
  1244 => (x"5c",x"5b",x"5e",x"0e"),
  1245 => (x"86",x"f4",x"0e",x"5d"),
  1246 => (x"c2",x"59",x"a6",x"c4"),
  1247 => (x"49",x"66",x"dc",x"4d"),
  1248 => (x"4c",x"6e",x"81",x"c1"),
  1249 => (x"4b",x"a1",x"84",x"c2"),
  1250 => (x"ff",x"c3",x"49",x"6b"),
  1251 => (x"48",x"a6",x"c4",x"99"),
  1252 => (x"97",x"c4",x"50",x"6c"),
  1253 => (x"b7",x"71",x"4a",x"66"),
  1254 => (x"87",x"c7",x"02",x"aa"),
  1255 => (x"c0",x"48",x"a6",x"c8"),
  1256 => (x"c1",x"87",x"cd",x"78"),
  1257 => (x"c4",x"48",x"c8",x"d0"),
  1258 => (x"c8",x"50",x"66",x"97"),
  1259 => (x"78",x"c1",x"48",x"a6"),
  1260 => (x"c4",x"05",x"66",x"c8"),
  1261 => (x"83",x"85",x"c1",x"87"),
  1262 => (x"ad",x"b7",x"c2",x"84"),
  1263 => (x"87",x"c8",x"ff",x"06"),
  1264 => (x"66",x"dc",x"4a",x"6e"),
  1265 => (x"d3",x"fe",x"fe",x"49"),
  1266 => (x"a8",x"b7",x"c0",x"87"),
  1267 => (x"c1",x"87",x"cb",x"06"),
  1268 => (x"c7",x"48",x"c0",x"d0"),
  1269 => (x"48",x"c1",x"78",x"a5"),
  1270 => (x"48",x"c0",x"87",x"c2"),
  1271 => (x"4d",x"26",x"8e",x"f4"),
  1272 => (x"4b",x"26",x"4c",x"26"),
  1273 => (x"4b",x"26",x"4f",x"26"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
