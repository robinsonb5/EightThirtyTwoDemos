
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"2c",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"29"),
    10 => (x"87",x"fd",x"00",x"4f"),
    11 => (x"cc",x"df",x"c1",x"4f"),
    12 => (x"c0",x"c0",x"c1",x"4e"),
    13 => (x"cc",x"df",x"c1",x"86"),
    14 => (x"f4",x"d4",x"c1",x"49"),
    15 => (x"89",x"d0",x"89",x"48"),
    16 => (x"40",x"40",x"c0",x"03"),
    17 => (x"87",x"f6",x"40",x"40"),
    18 => (x"c0",x"05",x"81",x"d0"),
    19 => (x"05",x"89",x"c1",x"50"),
    20 => (x"d4",x"c1",x"87",x"f9"),
    21 => (x"d4",x"c1",x"4d",x"f4"),
    22 => (x"ad",x"74",x"4c",x"f4"),
    23 => (x"24",x"87",x"c4",x"02"),
    24 => (x"d8",x"87",x"f7",x"0f"),
    25 => (x"d4",x"c1",x"87",x"ea"),
    26 => (x"d4",x"c1",x"4d",x"f4"),
    27 => (x"ad",x"74",x"4c",x"f4"),
    28 => (x"c4",x"87",x"c6",x"02"),
    29 => (x"f5",x"0f",x"6c",x"8c"),
    30 => (x"87",x"fd",x"00",x"87"),
    31 => (x"5c",x"5b",x"5e",x"0e"),
    32 => (x"86",x"fc",x"0e",x"5d"),
    33 => (x"e0",x"c0",x"4a",x"71"),
    34 => (x"d4",x"c1",x"4c",x"66"),
    35 => (x"7e",x"c0",x"4b",x"f4"),
    36 => (x"ce",x"05",x"9a",x"72"),
    37 => (x"f5",x"d4",x"c1",x"87"),
    38 => (x"f4",x"d4",x"c1",x"4b"),
    39 => (x"50",x"f0",x"c0",x"48"),
    40 => (x"72",x"87",x"d1",x"c1"),
    41 => (x"e8",x"c0",x"02",x"9a"),
    42 => (x"4d",x"66",x"d4",x"87"),
    43 => (x"49",x"72",x"1e",x"72"),
    44 => (x"ce",x"cb",x"4a",x"75"),
    45 => (x"c4",x"4a",x"26",x"87"),
    46 => (x"53",x"11",x"81",x"e5"),
    47 => (x"49",x"72",x"1e",x"71"),
    48 => (x"fe",x"ca",x"4a",x"75"),
    49 => (x"26",x"4a",x"70",x"87"),
    50 => (x"72",x"8c",x"c1",x"49"),
    51 => (x"db",x"ff",x"05",x"9a"),
    52 => (x"ac",x"b7",x"c0",x"87"),
    53 => (x"c0",x"87",x"dd",x"06"),
    54 => (x"c5",x"02",x"66",x"e4"),
    55 => (x"4a",x"f0",x"c0",x"87"),
    56 => (x"e0",x"c0",x"87",x"c3"),
    57 => (x"97",x"0a",x"73",x"4a"),
    58 => (x"83",x"c1",x"0a",x"7a"),
    59 => (x"ac",x"b7",x"c0",x"8c"),
    60 => (x"87",x"e3",x"ff",x"01"),
    61 => (x"ab",x"f4",x"d4",x"c1"),
    62 => (x"d8",x"87",x"de",x"02"),
    63 => (x"66",x"dc",x"4c",x"66"),
    64 => (x"97",x"8b",x"c1",x"1e"),
    65 => (x"0f",x"74",x"49",x"6b"),
    66 => (x"48",x"6e",x"86",x"c4"),
    67 => (x"a6",x"c4",x"80",x"c1"),
    68 => (x"f4",x"d4",x"c1",x"58"),
    69 => (x"e5",x"ff",x"05",x"ab"),
    70 => (x"fc",x"48",x"6e",x"87"),
    71 => (x"26",x"4d",x"26",x"8e"),
    72 => (x"26",x"4b",x"26",x"4c"),
    73 => (x"32",x"31",x"30",x"4f"),
    74 => (x"36",x"35",x"34",x"33"),
    75 => (x"41",x"39",x"38",x"37"),
    76 => (x"45",x"44",x"43",x"42"),
    77 => (x"5e",x"0e",x"00",x"46"),
    78 => (x"0e",x"5d",x"5c",x"5b"),
    79 => (x"4d",x"ff",x"4b",x"71"),
    80 => (x"9c",x"74",x"4c",x"13"),
    81 => (x"c1",x"87",x"d8",x"02"),
    82 => (x"1e",x"66",x"d4",x"85"),
    83 => (x"66",x"d4",x"49",x"74"),
    84 => (x"74",x"86",x"c4",x"0f"),
    85 => (x"87",x"c7",x"05",x"a8"),
    86 => (x"9c",x"74",x"4c",x"13"),
    87 => (x"75",x"87",x"e8",x"05"),
    88 => (x"26",x"4d",x"26",x"48"),
    89 => (x"26",x"4b",x"26",x"4c"),
    90 => (x"5b",x"5e",x"0e",x"4f"),
    91 => (x"e8",x"0e",x"5d",x"5c"),
    92 => (x"59",x"a6",x"c4",x"86"),
    93 => (x"4d",x"66",x"e8",x"c0"),
    94 => (x"a6",x"c8",x"4c",x"c0"),
    95 => (x"6e",x"78",x"c0",x"48"),
    96 => (x"6e",x"4b",x"bf",x"97"),
    97 => (x"c4",x"80",x"c1",x"48"),
    98 => (x"9b",x"73",x"58",x"a6"),
    99 => (x"87",x"d3",x"c6",x"02"),
   100 => (x"c5",x"02",x"66",x"c8"),
   101 => (x"a6",x"cc",x"87",x"db"),
   102 => (x"fc",x"78",x"c0",x"48"),
   103 => (x"73",x"78",x"c0",x"80"),
   104 => (x"8a",x"e0",x"c0",x"4a"),
   105 => (x"87",x"c6",x"c3",x"02"),
   106 => (x"c3",x"02",x"8a",x"c3"),
   107 => (x"8a",x"c2",x"87",x"c0"),
   108 => (x"87",x"e8",x"c2",x"02"),
   109 => (x"c2",x"02",x"8a",x"c2"),
   110 => (x"8a",x"c4",x"87",x"f4"),
   111 => (x"87",x"ee",x"c2",x"02"),
   112 => (x"c2",x"02",x"8a",x"c2"),
   113 => (x"8a",x"c3",x"87",x"e8"),
   114 => (x"87",x"ea",x"c2",x"02"),
   115 => (x"c0",x"02",x"8a",x"d4"),
   116 => (x"8a",x"d4",x"87",x"f6"),
   117 => (x"87",x"c0",x"c1",x"02"),
   118 => (x"c0",x"02",x"8a",x"ca"),
   119 => (x"8a",x"c1",x"87",x"f2"),
   120 => (x"87",x"e1",x"c1",x"02"),
   121 => (x"df",x"02",x"8a",x"c1"),
   122 => (x"02",x"8a",x"c8",x"87"),
   123 => (x"c4",x"87",x"ce",x"c1"),
   124 => (x"e3",x"c0",x"02",x"8a"),
   125 => (x"02",x"8a",x"c3",x"87"),
   126 => (x"c2",x"87",x"e5",x"c0"),
   127 => (x"87",x"c8",x"02",x"8a"),
   128 => (x"d3",x"02",x"8a",x"c3"),
   129 => (x"87",x"fa",x"c1",x"87"),
   130 => (x"ca",x"48",x"a6",x"cc"),
   131 => (x"87",x"d2",x"c2",x"78"),
   132 => (x"c2",x"48",x"a6",x"cc"),
   133 => (x"87",x"ca",x"c2",x"78"),
   134 => (x"d0",x"48",x"a6",x"cc"),
   135 => (x"87",x"c2",x"c2",x"78"),
   136 => (x"1e",x"66",x"f0",x"c0"),
   137 => (x"1e",x"66",x"f0",x"c0"),
   138 => (x"4a",x"75",x"85",x"c4"),
   139 => (x"49",x"6a",x"8a",x"c4"),
   140 => (x"c8",x"87",x"c3",x"fc"),
   141 => (x"71",x"49",x"70",x"86"),
   142 => (x"e5",x"c1",x"4c",x"a4"),
   143 => (x"48",x"a6",x"c8",x"87"),
   144 => (x"dd",x"c1",x"78",x"c1"),
   145 => (x"66",x"f0",x"c0",x"87"),
   146 => (x"75",x"85",x"c4",x"1e"),
   147 => (x"6a",x"8a",x"c4",x"4a"),
   148 => (x"66",x"f0",x"c0",x"49"),
   149 => (x"c1",x"86",x"c4",x"0f"),
   150 => (x"87",x"c6",x"c1",x"84"),
   151 => (x"1e",x"66",x"f0",x"c0"),
   152 => (x"c0",x"49",x"e5",x"c0"),
   153 => (x"c4",x"0f",x"66",x"f0"),
   154 => (x"c0",x"84",x"c1",x"86"),
   155 => (x"a6",x"c8",x"87",x"f4"),
   156 => (x"c0",x"78",x"c1",x"48"),
   157 => (x"a6",x"d0",x"87",x"ec"),
   158 => (x"f8",x"78",x"c1",x"48"),
   159 => (x"c0",x"78",x"c1",x"80"),
   160 => (x"f0",x"c0",x"87",x"e0"),
   161 => (x"87",x"da",x"06",x"ab"),
   162 => (x"03",x"ab",x"f9",x"c0"),
   163 => (x"66",x"d4",x"87",x"d4"),
   164 => (x"73",x"91",x"ca",x"49"),
   165 => (x"8a",x"f0",x"c0",x"4a"),
   166 => (x"72",x"48",x"a6",x"d4"),
   167 => (x"80",x"f4",x"78",x"a1"),
   168 => (x"66",x"cc",x"78",x"c1"),
   169 => (x"87",x"ea",x"c1",x"02"),
   170 => (x"49",x"75",x"85",x"c4"),
   171 => (x"48",x"a6",x"89",x"c4"),
   172 => (x"e4",x"c1",x"78",x"69"),
   173 => (x"87",x"d8",x"05",x"ab"),
   174 => (x"c0",x"48",x"66",x"c4"),
   175 => (x"cf",x"03",x"a8",x"b7"),
   176 => (x"49",x"ed",x"c0",x"87"),
   177 => (x"c4",x"87",x"fb",x"c1"),
   178 => (x"08",x"c0",x"48",x"66"),
   179 => (x"58",x"a6",x"c8",x"88"),
   180 => (x"d8",x"1e",x"66",x"d0"),
   181 => (x"f8",x"c0",x"1e",x"66"),
   182 => (x"f8",x"c0",x"1e",x"66"),
   183 => (x"66",x"dc",x"1e",x"66"),
   184 => (x"49",x"66",x"d8",x"1e"),
   185 => (x"d4",x"87",x"d5",x"f6"),
   186 => (x"71",x"49",x"70",x"86"),
   187 => (x"e1",x"c0",x"4c",x"a4"),
   188 => (x"ab",x"e5",x"c0",x"87"),
   189 => (x"d0",x"87",x"cf",x"05"),
   190 => (x"78",x"c0",x"48",x"a6"),
   191 => (x"78",x"c0",x"80",x"c4"),
   192 => (x"78",x"c1",x"80",x"f4"),
   193 => (x"f0",x"c0",x"87",x"cc"),
   194 => (x"49",x"73",x"1e",x"66"),
   195 => (x"0f",x"66",x"f0",x"c0"),
   196 => (x"97",x"6e",x"86",x"c4"),
   197 => (x"48",x"6e",x"4b",x"bf"),
   198 => (x"a6",x"c4",x"80",x"c1"),
   199 => (x"05",x"9b",x"73",x"58"),
   200 => (x"74",x"87",x"ed",x"f9"),
   201 => (x"26",x"8e",x"e8",x"48"),
   202 => (x"26",x"4c",x"26",x"4d"),
   203 => (x"1e",x"4f",x"26",x"4b"),
   204 => (x"c2",x"cd",x"1e",x"c0"),
   205 => (x"1e",x"a6",x"d0",x"1e"),
   206 => (x"f8",x"49",x"66",x"d0"),
   207 => (x"8e",x"f4",x"87",x"eb"),
   208 => (x"fc",x"1e",x"4f",x"26"),
   209 => (x"ff",x"4a",x"71",x"86"),
   210 => (x"48",x"69",x"49",x"c0"),
   211 => (x"c4",x"98",x"c0",x"c4"),
   212 => (x"02",x"6e",x"58",x"a6"),
   213 => (x"79",x"72",x"87",x"f4"),
   214 => (x"26",x"8e",x"fc",x"48"),
   215 => (x"5b",x"5e",x"0e",x"4f"),
   216 => (x"4b",x"71",x"0e",x"5c"),
   217 => (x"4a",x"13",x"4c",x"c0"),
   218 => (x"ce",x"02",x"9a",x"72"),
   219 => (x"ff",x"49",x"72",x"87"),
   220 => (x"84",x"c1",x"87",x"d0"),
   221 => (x"9a",x"72",x"4a",x"13"),
   222 => (x"74",x"87",x"f2",x"05"),
   223 => (x"26",x"4c",x"26",x"48"),
   224 => (x"1e",x"4f",x"26",x"4b"),
   225 => (x"9a",x"72",x"1e",x"73"),
   226 => (x"87",x"e7",x"c0",x"02"),
   227 => (x"4b",x"c1",x"48",x"c0"),
   228 => (x"d1",x"06",x"a9",x"72"),
   229 => (x"06",x"82",x"72",x"87"),
   230 => (x"83",x"73",x"87",x"c9"),
   231 => (x"f4",x"01",x"a9",x"72"),
   232 => (x"c1",x"87",x"c3",x"87"),
   233 => (x"a9",x"72",x"3a",x"b2"),
   234 => (x"80",x"73",x"89",x"03"),
   235 => (x"2b",x"2a",x"c1",x"07"),
   236 => (x"26",x"87",x"f3",x"05"),
   237 => (x"1e",x"4f",x"26",x"4b"),
   238 => (x"4d",x"c4",x"1e",x"75"),
   239 => (x"04",x"a1",x"b7",x"71"),
   240 => (x"81",x"c1",x"b9",x"ff"),
   241 => (x"72",x"07",x"bd",x"c3"),
   242 => (x"ff",x"04",x"a2",x"b7"),
   243 => (x"c1",x"82",x"c1",x"ba"),
   244 => (x"ee",x"fe",x"07",x"bd"),
   245 => (x"04",x"2d",x"c1",x"87"),
   246 => (x"80",x"c1",x"b8",x"ff"),
   247 => (x"ff",x"04",x"2d",x"07"),
   248 => (x"07",x"81",x"c1",x"b9"),
   249 => (x"4f",x"26",x"4d",x"26"),
   250 => (x"d0",x"1e",x"73",x"1e"),
   251 => (x"c0",x"c0",x"c0",x"c0"),
   252 => (x"fe",x"0f",x"73",x"4b"),
   253 => (x"26",x"87",x"c4",x"87"),
   254 => (x"26",x"4c",x"26",x"4d"),
   255 => (x"1e",x"4f",x"26",x"4b"),
   256 => (x"c3",x"4a",x"66",x"c4"),
   257 => (x"f7",x"c0",x"9a",x"df"),
   258 => (x"aa",x"b7",x"c0",x"8a"),
   259 => (x"c0",x"87",x"c3",x"03"),
   260 => (x"31",x"c4",x"82",x"e7"),
   261 => (x"48",x"71",x"b1",x"72"),
   262 => (x"5e",x"0e",x"4f",x"26"),
   263 => (x"0e",x"5d",x"5c",x"5b"),
   264 => (x"c0",x"d0",x"4a",x"71"),
   265 => (x"4d",x"c0",x"c0",x"c0"),
   266 => (x"bf",x"c4",x"d5",x"c1"),
   267 => (x"c1",x"80",x"c1",x"48"),
   268 => (x"72",x"58",x"c8",x"d5"),
   269 => (x"81",x"c0",x"fe",x"49"),
   270 => (x"a9",x"d3",x"c1",x"b9"),
   271 => (x"c1",x"87",x"db",x"05"),
   272 => (x"c0",x"48",x"c4",x"d5"),
   273 => (x"c8",x"d5",x"c1",x"78"),
   274 => (x"c1",x"78",x"c0",x"48"),
   275 => (x"c0",x"48",x"d0",x"d5"),
   276 => (x"d4",x"d5",x"c1",x"78"),
   277 => (x"c6",x"78",x"c0",x"48"),
   278 => (x"d5",x"c1",x"87",x"ea"),
   279 => (x"c1",x"48",x"bf",x"c4"),
   280 => (x"f6",x"c0",x"05",x"a8"),
   281 => (x"fe",x"49",x"72",x"87"),
   282 => (x"71",x"b9",x"81",x"c0"),
   283 => (x"d4",x"d5",x"c1",x"1e"),
   284 => (x"ca",x"fe",x"49",x"bf"),
   285 => (x"c1",x"86",x"c4",x"87"),
   286 => (x"c1",x"58",x"d8",x"d5"),
   287 => (x"4b",x"bf",x"d4",x"d5"),
   288 => (x"06",x"ab",x"b7",x"c3"),
   289 => (x"48",x"ca",x"87",x"c6"),
   290 => (x"4b",x"70",x"88",x"73"),
   291 => (x"81",x"c1",x"49",x"73"),
   292 => (x"30",x"c1",x"48",x"71"),
   293 => (x"58",x"d0",x"d5",x"c1"),
   294 => (x"c1",x"87",x"e9",x"c5"),
   295 => (x"48",x"bf",x"d4",x"d5"),
   296 => (x"01",x"a8",x"b7",x"c9"),
   297 => (x"c1",x"87",x"dd",x"c5"),
   298 => (x"48",x"bf",x"d4",x"d5"),
   299 => (x"06",x"a8",x"b7",x"c0"),
   300 => (x"c1",x"87",x"d1",x"c5"),
   301 => (x"48",x"bf",x"c4",x"d5"),
   302 => (x"01",x"a8",x"b7",x"c3"),
   303 => (x"49",x"72",x"87",x"d9"),
   304 => (x"b9",x"81",x"c0",x"fe"),
   305 => (x"d5",x"c1",x"1e",x"71"),
   306 => (x"fc",x"49",x"bf",x"d0"),
   307 => (x"86",x"c4",x"87",x"f1"),
   308 => (x"58",x"d4",x"d5",x"c1"),
   309 => (x"c1",x"87",x"ed",x"c4"),
   310 => (x"49",x"bf",x"cc",x"d5"),
   311 => (x"d5",x"c1",x"81",x"c3"),
   312 => (x"a9",x"b7",x"bf",x"c4"),
   313 => (x"72",x"87",x"df",x"04"),
   314 => (x"81",x"c0",x"fe",x"49"),
   315 => (x"c1",x"1e",x"71",x"b9"),
   316 => (x"49",x"bf",x"c8",x"d5"),
   317 => (x"c4",x"87",x"c8",x"fc"),
   318 => (x"cc",x"d5",x"c1",x"86"),
   319 => (x"d8",x"d5",x"c1",x"58"),
   320 => (x"c3",x"78",x"c1",x"48"),
   321 => (x"d5",x"c1",x"87",x"fe"),
   322 => (x"c0",x"48",x"bf",x"d4"),
   323 => (x"c2",x"06",x"a8",x"b7"),
   324 => (x"d5",x"c1",x"87",x"d5"),
   325 => (x"c3",x"48",x"bf",x"d4"),
   326 => (x"c2",x"01",x"a8",x"b7"),
   327 => (x"d5",x"c1",x"87",x"c9"),
   328 => (x"c1",x"49",x"bf",x"d0"),
   329 => (x"d5",x"c1",x"81",x"31"),
   330 => (x"a9",x"b7",x"bf",x"c4"),
   331 => (x"87",x"d9",x"c1",x"04"),
   332 => (x"c0",x"fe",x"49",x"72"),
   333 => (x"1e",x"71",x"b9",x"81"),
   334 => (x"bf",x"dc",x"d5",x"c1"),
   335 => (x"87",x"ff",x"fa",x"49"),
   336 => (x"d5",x"c1",x"86",x"c4"),
   337 => (x"d5",x"c1",x"58",x"e0"),
   338 => (x"c1",x"49",x"bf",x"d8"),
   339 => (x"dc",x"d5",x"c1",x"89"),
   340 => (x"a9",x"b7",x"c0",x"59"),
   341 => (x"87",x"ec",x"c2",x"03"),
   342 => (x"bf",x"c8",x"d5",x"c1"),
   343 => (x"dc",x"d5",x"c1",x"49"),
   344 => (x"d5",x"c1",x"51",x"bf"),
   345 => (x"c1",x"49",x"bf",x"c8"),
   346 => (x"cc",x"d5",x"c1",x"81"),
   347 => (x"e0",x"d5",x"c1",x"59"),
   348 => (x"06",x"a9",x"b7",x"bf"),
   349 => (x"c1",x"87",x"c9",x"c0"),
   350 => (x"c1",x"48",x"e0",x"d5"),
   351 => (x"78",x"bf",x"c8",x"d5"),
   352 => (x"48",x"d8",x"d5",x"c1"),
   353 => (x"fb",x"c1",x"78",x"c1"),
   354 => (x"d8",x"d5",x"c1",x"87"),
   355 => (x"f3",x"c1",x"05",x"bf"),
   356 => (x"dc",x"d5",x"c1",x"87"),
   357 => (x"31",x"c4",x"49",x"bf"),
   358 => (x"59",x"e0",x"d5",x"c1"),
   359 => (x"bf",x"c8",x"d5",x"c1"),
   360 => (x"09",x"79",x"97",x"09"),
   361 => (x"c1",x"87",x"dd",x"c1"),
   362 => (x"48",x"bf",x"d4",x"d5"),
   363 => (x"04",x"a8",x"b7",x"c7"),
   364 => (x"c0",x"87",x"d1",x"c1"),
   365 => (x"48",x"f4",x"fe",x"4c"),
   366 => (x"d5",x"c1",x"78",x"c1"),
   367 => (x"75",x"1e",x"bf",x"e0"),
   368 => (x"1e",x"c7",x"d8",x"1e"),
   369 => (x"cc",x"87",x"e8",x"f5"),
   370 => (x"cc",x"d5",x"c1",x"86"),
   371 => (x"c8",x"d5",x"c1",x"5d"),
   372 => (x"d5",x"c1",x"48",x"bf"),
   373 => (x"a8",x"b7",x"bf",x"e0"),
   374 => (x"87",x"db",x"c0",x"03"),
   375 => (x"bf",x"c8",x"d5",x"c1"),
   376 => (x"d5",x"c1",x"84",x"bf"),
   377 => (x"c4",x"49",x"bf",x"c8"),
   378 => (x"cc",x"d5",x"c1",x"81"),
   379 => (x"e0",x"d5",x"c1",x"59"),
   380 => (x"04",x"a9",x"b7",x"bf"),
   381 => (x"74",x"87",x"e5",x"ff"),
   382 => (x"1e",x"e6",x"d8",x"1e"),
   383 => (x"c8",x"87",x"f0",x"f4"),
   384 => (x"87",x"e4",x"f7",x"86"),
   385 => (x"43",x"87",x"f0",x"f7"),
   386 => (x"6b",x"63",x"65",x"68"),
   387 => (x"6d",x"6d",x"75",x"73"),
   388 => (x"20",x"67",x"6e",x"69"),
   389 => (x"6d",x"6f",x"72",x"66"),
   390 => (x"20",x"64",x"25",x"20"),
   391 => (x"25",x"20",x"6f",x"74"),
   392 => (x"2e",x"2e",x"2e",x"64"),
   393 => (x"64",x"25",x"00",x"20"),
   394 => (x"6f",x"42",x"00",x"0a"),
   395 => (x"6e",x"69",x"74",x"6f"),
   396 => (x"2e",x"2e",x"2e",x"67"),
   397 => (x"4f",x"42",x"00",x"0a"),
   398 => (x"33",x"38",x"54",x"4f"),
   399 => (x"49",x"42",x"20",x"32"),
   400 => (x"44",x"53",x"00",x"4e"),
   401 => (x"6f",x"6f",x"62",x"20"),
   402 => (x"61",x"66",x"20",x"74"),
   403 => (x"64",x"65",x"6c",x"69"),
   404 => (x"6e",x"49",x"00",x"0a"),
   405 => (x"61",x"69",x"74",x"69"),
   406 => (x"69",x"7a",x"69",x"6c"),
   407 => (x"53",x"20",x"67",x"6e"),
   408 => (x"61",x"63",x"20",x"44"),
   409 => (x"00",x"0a",x"64",x"72"),
   410 => (x"33",x"32",x"53",x"52"),
   411 => (x"6f",x"62",x"20",x"32"),
   412 => (x"2d",x"20",x"74",x"6f"),
   413 => (x"65",x"72",x"70",x"20"),
   414 => (x"45",x"20",x"73",x"73"),
   415 => (x"74",x"20",x"43",x"53"),
   416 => (x"6f",x"62",x"20",x"6f"),
   417 => (x"66",x"20",x"74",x"6f"),
   418 => (x"20",x"6d",x"6f",x"72"),
   419 => (x"00",x"2e",x"44",x"53"),
   420 => (x"5c",x"5b",x"5e",x"0e"),
   421 => (x"d9",x"1e",x"0e",x"5d"),
   422 => (x"c0",x"f3",x"49",x"d2"),
   423 => (x"d5",x"ed",x"c0",x"87"),
   424 => (x"02",x"98",x"70",x"87"),
   425 => (x"ca",x"c3",x"87",x"cc"),
   426 => (x"02",x"98",x"70",x"87"),
   427 => (x"4b",x"c1",x"87",x"c4"),
   428 => (x"4b",x"c0",x"87",x"c2"),
   429 => (x"d9",x"5b",x"a6",x"c4"),
   430 => (x"e0",x"f2",x"49",x"e8"),
   431 => (x"e0",x"d5",x"c1",x"87"),
   432 => (x"c0",x"78",x"c0",x"48"),
   433 => (x"f9",x"f1",x"49",x"ee"),
   434 => (x"c8",x"f4",x"c3",x"87"),
   435 => (x"c0",x"ff",x"4a",x"ff"),
   436 => (x"49",x"73",x"4b",x"bf"),
   437 => (x"02",x"99",x"c0",x"c8"),
   438 => (x"73",x"87",x"fd",x"c0"),
   439 => (x"9c",x"ff",x"c3",x"4c"),
   440 => (x"c0",x"05",x"ac",x"db"),
   441 => (x"02",x"6e",x"87",x"e8"),
   442 => (x"c0",x"d0",x"87",x"de"),
   443 => (x"1e",x"c0",x"c0",x"c0"),
   444 => (x"db",x"49",x"f6",x"d8"),
   445 => (x"86",x"c4",x"87",x"f7"),
   446 => (x"cb",x"02",x"98",x"70"),
   447 => (x"49",x"ea",x"d8",x"87"),
   448 => (x"f3",x"87",x"da",x"f1"),
   449 => (x"87",x"c6",x"87",x"e2"),
   450 => (x"f1",x"49",x"c2",x"d9"),
   451 => (x"49",x"74",x"87",x"cf"),
   452 => (x"c3",x"87",x"c7",x"f4"),
   453 => (x"4a",x"c0",x"c9",x"f4"),
   454 => (x"8a",x"c1",x"49",x"72"),
   455 => (x"fe",x"05",x"99",x"71"),
   456 => (x"de",x"fe",x"87",x"ec"),
   457 => (x"ce",x"f3",x"26",x"87"),
   458 => (x"5b",x"5e",x"0e",x"87"),
   459 => (x"4b",x"71",x"0e",x"5c"),
   460 => (x"66",x"d0",x"4c",x"c0"),
   461 => (x"a8",x"b7",x"c0",x"48"),
   462 => (x"87",x"eb",x"c0",x"06"),
   463 => (x"c0",x"fe",x"4a",x"13"),
   464 => (x"66",x"cc",x"ba",x"82"),
   465 => (x"fe",x"49",x"bf",x"97"),
   466 => (x"cc",x"b9",x"81",x"c0"),
   467 => (x"80",x"c1",x"48",x"66"),
   468 => (x"71",x"58",x"a6",x"d0"),
   469 => (x"c4",x"02",x"aa",x"b7"),
   470 => (x"cc",x"48",x"c1",x"87"),
   471 => (x"d0",x"84",x"c1",x"87"),
   472 => (x"04",x"ac",x"b7",x"66"),
   473 => (x"c0",x"87",x"d5",x"ff"),
   474 => (x"26",x"87",x"c2",x"48"),
   475 => (x"26",x"4c",x"26",x"4d"),
   476 => (x"0e",x"4f",x"26",x"4b"),
   477 => (x"5d",x"5c",x"5b",x"5e"),
   478 => (x"ec",x"dd",x"c1",x"0e"),
   479 => (x"c0",x"78",x"c0",x"48"),
   480 => (x"ef",x"49",x"c1",x"ed"),
   481 => (x"d5",x"c1",x"87",x"d7"),
   482 => (x"49",x"c0",x"1e",x"e4"),
   483 => (x"87",x"cb",x"ef",x"c0"),
   484 => (x"98",x"70",x"86",x"c4"),
   485 => (x"c0",x"87",x"cc",x"05"),
   486 => (x"ee",x"49",x"ed",x"e9"),
   487 => (x"48",x"c0",x"87",x"ff"),
   488 => (x"c0",x"87",x"c7",x"cb"),
   489 => (x"ee",x"49",x"ce",x"ed"),
   490 => (x"4b",x"c0",x"87",x"f3"),
   491 => (x"48",x"d8",x"de",x"c1"),
   492 => (x"1e",x"c8",x"78",x"c1"),
   493 => (x"1e",x"e5",x"ed",x"c0"),
   494 => (x"49",x"da",x"d6",x"c1"),
   495 => (x"c8",x"87",x"ea",x"fd"),
   496 => (x"05",x"98",x"70",x"86"),
   497 => (x"de",x"c1",x"87",x"c6"),
   498 => (x"78",x"c0",x"48",x"d8"),
   499 => (x"ed",x"c0",x"1e",x"c8"),
   500 => (x"d6",x"c1",x"1e",x"ee"),
   501 => (x"d0",x"fd",x"49",x"f6"),
   502 => (x"70",x"86",x"c8",x"87"),
   503 => (x"87",x"c6",x"05",x"98"),
   504 => (x"48",x"d8",x"de",x"c1"),
   505 => (x"de",x"c1",x"78",x"c0"),
   506 => (x"c0",x"1e",x"bf",x"d8"),
   507 => (x"ec",x"1e",x"f7",x"ed"),
   508 => (x"86",x"c8",x"87",x"fd"),
   509 => (x"bf",x"d8",x"de",x"c1"),
   510 => (x"87",x"cd",x"c2",x"02"),
   511 => (x"4d",x"e4",x"d5",x"c1"),
   512 => (x"a0",x"fe",x"c6",x"48"),
   513 => (x"e2",x"dd",x"c1",x"4c"),
   514 => (x"71",x"49",x"bf",x"9f"),
   515 => (x"80",x"fe",x"c7",x"1e"),
   516 => (x"f8",x"48",x"49",x"70"),
   517 => (x"71",x"89",x"a0",x"c2"),
   518 => (x"c8",x"1e",x"d0",x"1e"),
   519 => (x"ea",x"c0",x"1e",x"c0"),
   520 => (x"ca",x"ec",x"1e",x"df"),
   521 => (x"c8",x"86",x"d4",x"87"),
   522 => (x"4b",x"69",x"49",x"a4"),
   523 => (x"9f",x"e2",x"dd",x"c1"),
   524 => (x"d6",x"c5",x"49",x"bf"),
   525 => (x"c0",x"05",x"a9",x"ea"),
   526 => (x"a4",x"c8",x"87",x"cd"),
   527 => (x"c0",x"49",x"6a",x"4a"),
   528 => (x"70",x"87",x"fd",x"f2"),
   529 => (x"c7",x"87",x"db",x"4b"),
   530 => (x"9f",x"49",x"a5",x"fe"),
   531 => (x"e9",x"ca",x"49",x"69"),
   532 => (x"c0",x"02",x"a9",x"d5"),
   533 => (x"ea",x"c0",x"87",x"cc"),
   534 => (x"c0",x"ec",x"49",x"c1"),
   535 => (x"c8",x"48",x"c0",x"87"),
   536 => (x"1e",x"73",x"87",x"c8"),
   537 => (x"1e",x"dc",x"eb",x"c0"),
   538 => (x"c1",x"87",x"c4",x"eb"),
   539 => (x"73",x"1e",x"e4",x"d5"),
   540 => (x"e6",x"eb",x"c0",x"49"),
   541 => (x"70",x"86",x"cc",x"87"),
   542 => (x"c5",x"c0",x"05",x"98"),
   543 => (x"c7",x"48",x"c0",x"87"),
   544 => (x"eb",x"c0",x"87",x"e8"),
   545 => (x"d4",x"eb",x"49",x"f4"),
   546 => (x"ca",x"ee",x"c0",x"87"),
   547 => (x"87",x"df",x"ea",x"1e"),
   548 => (x"ee",x"c0",x"1e",x"c8"),
   549 => (x"d6",x"c1",x"1e",x"e2"),
   550 => (x"cc",x"fa",x"49",x"f6"),
   551 => (x"70",x"86",x"cc",x"87"),
   552 => (x"c9",x"c0",x"05",x"98"),
   553 => (x"ec",x"dd",x"c1",x"87"),
   554 => (x"c0",x"78",x"c1",x"48"),
   555 => (x"1e",x"c8",x"87",x"e3"),
   556 => (x"1e",x"eb",x"ee",x"c0"),
   557 => (x"49",x"da",x"d6",x"c1"),
   558 => (x"c8",x"87",x"ee",x"f9"),
   559 => (x"02",x"98",x"70",x"86"),
   560 => (x"c0",x"87",x"ce",x"c0"),
   561 => (x"e9",x"1e",x"db",x"ec"),
   562 => (x"86",x"c4",x"87",x"e5"),
   563 => (x"d9",x"c6",x"48",x"c0"),
   564 => (x"e2",x"dd",x"c1",x"87"),
   565 => (x"c1",x"49",x"bf",x"97"),
   566 => (x"c0",x"05",x"a9",x"d5"),
   567 => (x"dd",x"c1",x"87",x"cd"),
   568 => (x"49",x"bf",x"97",x"e3"),
   569 => (x"02",x"a9",x"ea",x"c2"),
   570 => (x"c0",x"87",x"c5",x"c0"),
   571 => (x"87",x"fa",x"c5",x"48"),
   572 => (x"97",x"e4",x"d5",x"c1"),
   573 => (x"e9",x"c3",x"49",x"bf"),
   574 => (x"d2",x"c0",x"02",x"a9"),
   575 => (x"e4",x"d5",x"c1",x"87"),
   576 => (x"c3",x"49",x"bf",x"97"),
   577 => (x"c0",x"02",x"a9",x"eb"),
   578 => (x"48",x"c0",x"87",x"c5"),
   579 => (x"c1",x"87",x"db",x"c5"),
   580 => (x"bf",x"97",x"ef",x"d5"),
   581 => (x"05",x"99",x"71",x"49"),
   582 => (x"c1",x"87",x"cc",x"c0"),
   583 => (x"bf",x"97",x"f0",x"d5"),
   584 => (x"02",x"a9",x"c2",x"49"),
   585 => (x"c0",x"87",x"c5",x"c0"),
   586 => (x"87",x"fe",x"c4",x"48"),
   587 => (x"97",x"f1",x"d5",x"c1"),
   588 => (x"dd",x"c1",x"48",x"bf"),
   589 => (x"dd",x"c1",x"58",x"e8"),
   590 => (x"71",x"49",x"bf",x"e4"),
   591 => (x"c1",x"8a",x"c1",x"4a"),
   592 => (x"72",x"5a",x"ec",x"dd"),
   593 => (x"c0",x"1e",x"71",x"1e"),
   594 => (x"e7",x"1e",x"f4",x"ee"),
   595 => (x"86",x"cc",x"87",x"e1"),
   596 => (x"97",x"f2",x"d5",x"c1"),
   597 => (x"81",x"73",x"49",x"bf"),
   598 => (x"97",x"f3",x"d5",x"c1"),
   599 => (x"32",x"c8",x"4a",x"bf"),
   600 => (x"48",x"f8",x"dd",x"c1"),
   601 => (x"c1",x"78",x"a1",x"72"),
   602 => (x"bf",x"97",x"f4",x"d5"),
   603 => (x"d0",x"de",x"c1",x"48"),
   604 => (x"ec",x"dd",x"c1",x"58"),
   605 => (x"df",x"c2",x"02",x"bf"),
   606 => (x"c0",x"1e",x"c8",x"87"),
   607 => (x"c1",x"1e",x"f8",x"ec"),
   608 => (x"f6",x"49",x"f6",x"d6"),
   609 => (x"86",x"c8",x"87",x"e3"),
   610 => (x"c0",x"02",x"98",x"70"),
   611 => (x"48",x"c0",x"87",x"c5"),
   612 => (x"c1",x"87",x"d7",x"c3"),
   613 => (x"4a",x"bf",x"e4",x"dd"),
   614 => (x"30",x"c4",x"48",x"72"),
   615 => (x"58",x"d4",x"de",x"c1"),
   616 => (x"5a",x"cc",x"de",x"c1"),
   617 => (x"97",x"c9",x"d6",x"c1"),
   618 => (x"31",x"c8",x"49",x"bf"),
   619 => (x"97",x"c8",x"d6",x"c1"),
   620 => (x"a1",x"73",x"4b",x"bf"),
   621 => (x"ca",x"d6",x"c1",x"49"),
   622 => (x"d0",x"4b",x"bf",x"97"),
   623 => (x"49",x"a1",x"73",x"33"),
   624 => (x"97",x"cb",x"d6",x"c1"),
   625 => (x"33",x"d8",x"4b",x"bf"),
   626 => (x"c1",x"49",x"a1",x"73"),
   627 => (x"c1",x"59",x"d8",x"de"),
   628 => (x"91",x"bf",x"cc",x"de"),
   629 => (x"bf",x"f8",x"dd",x"c1"),
   630 => (x"c0",x"de",x"c1",x"81"),
   631 => (x"d1",x"d6",x"c1",x"59"),
   632 => (x"c8",x"4b",x"bf",x"97"),
   633 => (x"d0",x"d6",x"c1",x"33"),
   634 => (x"74",x"4c",x"bf",x"97"),
   635 => (x"d6",x"c1",x"4b",x"a3"),
   636 => (x"4c",x"bf",x"97",x"d2"),
   637 => (x"a3",x"74",x"34",x"d0"),
   638 => (x"d3",x"d6",x"c1",x"4b"),
   639 => (x"cf",x"4c",x"bf",x"97"),
   640 => (x"74",x"34",x"d8",x"9c"),
   641 => (x"de",x"c1",x"4b",x"a3"),
   642 => (x"8b",x"c2",x"5b",x"c4"),
   643 => (x"de",x"c1",x"92",x"73"),
   644 => (x"a1",x"72",x"48",x"c4"),
   645 => (x"87",x"d0",x"c1",x"78"),
   646 => (x"97",x"f6",x"d5",x"c1"),
   647 => (x"31",x"c8",x"49",x"bf"),
   648 => (x"97",x"f5",x"d5",x"c1"),
   649 => (x"a1",x"72",x"4a",x"bf"),
   650 => (x"d4",x"de",x"c1",x"49"),
   651 => (x"c7",x"31",x"c5",x"59"),
   652 => (x"29",x"c9",x"81",x"ff"),
   653 => (x"59",x"cc",x"de",x"c1"),
   654 => (x"97",x"fb",x"d5",x"c1"),
   655 => (x"32",x"c8",x"4a",x"bf"),
   656 => (x"97",x"fa",x"d5",x"c1"),
   657 => (x"a2",x"73",x"4b",x"bf"),
   658 => (x"d8",x"de",x"c1",x"4a"),
   659 => (x"cc",x"de",x"c1",x"5a"),
   660 => (x"dd",x"c1",x"92",x"bf"),
   661 => (x"c1",x"82",x"bf",x"f8"),
   662 => (x"c1",x"5a",x"c8",x"de"),
   663 => (x"c0",x"48",x"c0",x"de"),
   664 => (x"fc",x"dd",x"c1",x"78"),
   665 => (x"78",x"a1",x"72",x"48"),
   666 => (x"fe",x"f3",x"48",x"c1"),
   667 => (x"61",x"65",x"52",x"87"),
   668 => (x"66",x"6f",x"20",x"64"),
   669 => (x"52",x"42",x"4d",x"20"),
   670 => (x"69",x"61",x"66",x"20"),
   671 => (x"0a",x"64",x"65",x"6c"),
   672 => (x"20",x"6f",x"4e",x"00"),
   673 => (x"74",x"72",x"61",x"70"),
   674 => (x"6f",x"69",x"74",x"69"),
   675 => (x"69",x"73",x"20",x"6e"),
   676 => (x"74",x"61",x"6e",x"67"),
   677 => (x"20",x"65",x"72",x"75"),
   678 => (x"6e",x"75",x"6f",x"66"),
   679 => (x"4d",x"00",x"0a",x"64"),
   680 => (x"69",x"73",x"52",x"42"),
   681 => (x"20",x"3a",x"65",x"7a"),
   682 => (x"20",x"2c",x"64",x"25"),
   683 => (x"74",x"72",x"61",x"70"),
   684 => (x"6f",x"69",x"74",x"69"),
   685 => (x"7a",x"69",x"73",x"6e"),
   686 => (x"25",x"20",x"3a",x"65"),
   687 => (x"6f",x"20",x"2c",x"64"),
   688 => (x"65",x"73",x"66",x"66"),
   689 => (x"66",x"6f",x"20",x"74"),
   690 => (x"67",x"69",x"73",x"20"),
   691 => (x"64",x"25",x"20",x"3a"),
   692 => (x"69",x"73",x"20",x"2c"),
   693 => (x"78",x"30",x"20",x"67"),
   694 => (x"00",x"0a",x"78",x"25"),
   695 => (x"64",x"61",x"65",x"52"),
   696 => (x"20",x"67",x"6e",x"69"),
   697 => (x"74",x"6f",x"6f",x"62"),
   698 => (x"63",x"65",x"73",x"20"),
   699 => (x"20",x"72",x"6f",x"74"),
   700 => (x"00",x"0a",x"64",x"25"),
   701 => (x"64",x"61",x"65",x"52"),
   702 => (x"6f",x"6f",x"62",x"20"),
   703 => (x"65",x"73",x"20",x"74"),
   704 => (x"72",x"6f",x"74",x"63"),
   705 => (x"6f",x"72",x"66",x"20"),
   706 => (x"69",x"66",x"20",x"6d"),
   707 => (x"20",x"74",x"73",x"72"),
   708 => (x"74",x"72",x"61",x"70"),
   709 => (x"6f",x"69",x"74",x"69"),
   710 => (x"55",x"00",x"0a",x"6e"),
   711 => (x"70",x"75",x"73",x"6e"),
   712 => (x"74",x"72",x"6f",x"70"),
   713 => (x"70",x"20",x"64",x"65"),
   714 => (x"69",x"74",x"72",x"61"),
   715 => (x"6e",x"6f",x"69",x"74"),
   716 => (x"70",x"79",x"74",x"20"),
   717 => (x"00",x"0d",x"21",x"65"),
   718 => (x"33",x"54",x"41",x"46"),
   719 => (x"20",x"20",x"20",x"32"),
   720 => (x"61",x"65",x"52",x"00"),
   721 => (x"67",x"6e",x"69",x"64"),
   722 => (x"52",x"42",x"4d",x"20"),
   723 => (x"42",x"4d",x"00",x"0a"),
   724 => (x"75",x"73",x"20",x"52"),
   725 => (x"73",x"65",x"63",x"63"),
   726 => (x"6c",x"75",x"66",x"73"),
   727 => (x"72",x"20",x"79",x"6c"),
   728 => (x"0a",x"64",x"61",x"65"),
   729 => (x"54",x"41",x"46",x"00"),
   730 => (x"20",x"20",x"36",x"31"),
   731 => (x"41",x"46",x"00",x"20"),
   732 => (x"20",x"32",x"33",x"54"),
   733 => (x"50",x"00",x"20",x"20"),
   734 => (x"69",x"74",x"72",x"61"),
   735 => (x"6e",x"6f",x"69",x"74"),
   736 => (x"6e",x"75",x"6f",x"63"),
   737 => (x"64",x"25",x"20",x"74"),
   738 => (x"75",x"48",x"00",x"0a"),
   739 => (x"6e",x"69",x"74",x"6e"),
   740 => (x"6f",x"66",x"20",x"67"),
   741 => (x"69",x"66",x"20",x"72"),
   742 => (x"79",x"73",x"65",x"6c"),
   743 => (x"6d",x"65",x"74",x"73"),
   744 => (x"41",x"46",x"00",x"0a"),
   745 => (x"20",x"32",x"33",x"54"),
   746 => (x"46",x"00",x"20",x"20"),
   747 => (x"36",x"31",x"54",x"41"),
   748 => (x"00",x"20",x"20",x"20"),
   749 => (x"73",x"75",x"6c",x"43"),
   750 => (x"20",x"72",x"65",x"74"),
   751 => (x"65",x"7a",x"69",x"73"),
   752 => (x"64",x"25",x"20",x"3a"),
   753 => (x"6c",x"43",x"20",x"2c"),
   754 => (x"65",x"74",x"73",x"75"),
   755 => (x"61",x"6d",x"20",x"72"),
   756 => (x"20",x"2c",x"6b",x"73"),
   757 => (x"00",x"0a",x"64",x"25"),
   758 => (x"6e",x"65",x"70",x"4f"),
   759 => (x"66",x"20",x"64",x"65"),
   760 => (x"2c",x"65",x"6c",x"69"),
   761 => (x"61",x"6f",x"6c",x"20"),
   762 => (x"67",x"6e",x"69",x"64"),
   763 => (x"0a",x"2e",x"2e",x"2e"),
   764 => (x"6e",x"61",x"43",x"00"),
   765 => (x"6f",x"20",x"74",x"27"),
   766 => (x"20",x"6e",x"65",x"70"),
   767 => (x"00",x"0a",x"73",x"25"),
   768 => (x"5c",x"5b",x"5e",x"0e"),
   769 => (x"4a",x"71",x"0e",x"5d"),
   770 => (x"bf",x"ec",x"dd",x"c1"),
   771 => (x"72",x"87",x"cc",x"02"),
   772 => (x"2b",x"b7",x"c7",x"4b"),
   773 => (x"ff",x"c1",x"4d",x"72"),
   774 => (x"72",x"87",x"ca",x"9d"),
   775 => (x"2b",x"b7",x"c8",x"4b"),
   776 => (x"ff",x"c3",x"4d",x"72"),
   777 => (x"e4",x"d5",x"c1",x"9d"),
   778 => (x"f8",x"dd",x"c1",x"1e"),
   779 => (x"81",x"73",x"49",x"bf"),
   780 => (x"e6",x"dc",x"49",x"71"),
   781 => (x"70",x"86",x"c4",x"87"),
   782 => (x"87",x"c5",x"05",x"98"),
   783 => (x"e6",x"c0",x"48",x"c0"),
   784 => (x"ec",x"dd",x"c1",x"87"),
   785 => (x"87",x"d2",x"02",x"bf"),
   786 => (x"91",x"c4",x"49",x"75"),
   787 => (x"81",x"e4",x"d5",x"c1"),
   788 => (x"ff",x"cf",x"4c",x"69"),
   789 => (x"9c",x"ff",x"ff",x"ff"),
   790 => (x"49",x"75",x"87",x"cb"),
   791 => (x"d5",x"c1",x"91",x"c2"),
   792 => (x"69",x"9f",x"81",x"e4"),
   793 => (x"ec",x"48",x"74",x"4c"),
   794 => (x"5e",x"0e",x"87",x"c1"),
   795 => (x"0e",x"5d",x"5c",x"5b"),
   796 => (x"4c",x"71",x"86",x"f4"),
   797 => (x"de",x"c1",x"4b",x"c0"),
   798 => (x"c1",x"4d",x"bf",x"c0"),
   799 => (x"7e",x"bf",x"c4",x"de"),
   800 => (x"bf",x"ec",x"dd",x"c1"),
   801 => (x"c1",x"87",x"c9",x"02"),
   802 => (x"4a",x"bf",x"e4",x"dd"),
   803 => (x"87",x"c7",x"32",x"c4"),
   804 => (x"bf",x"c8",x"de",x"c1"),
   805 => (x"c8",x"32",x"c4",x"4a"),
   806 => (x"a6",x"c8",x"5a",x"a6"),
   807 => (x"c4",x"78",x"c0",x"48"),
   808 => (x"a8",x"c0",x"48",x"66"),
   809 => (x"87",x"ee",x"c2",x"06"),
   810 => (x"cf",x"49",x"66",x"c8"),
   811 => (x"87",x"da",x"05",x"99"),
   812 => (x"1e",x"e4",x"d5",x"c1"),
   813 => (x"48",x"49",x"66",x"c4"),
   814 => (x"a6",x"c8",x"80",x"c1"),
   815 => (x"da",x"49",x"71",x"58"),
   816 => (x"86",x"c4",x"87",x"d9"),
   817 => (x"4b",x"e4",x"d5",x"c1"),
   818 => (x"e0",x"c0",x"87",x"c3"),
   819 => (x"49",x"6b",x"97",x"83"),
   820 => (x"c1",x"02",x"99",x"71"),
   821 => (x"6b",x"97",x"87",x"ee"),
   822 => (x"a9",x"e5",x"c3",x"49"),
   823 => (x"87",x"e4",x"c1",x"02"),
   824 => (x"97",x"49",x"a3",x"cb"),
   825 => (x"99",x"d8",x"49",x"69"),
   826 => (x"87",x"d8",x"c1",x"05"),
   827 => (x"d9",x"ff",x"49",x"73"),
   828 => (x"1e",x"cb",x"87",x"eb"),
   829 => (x"1e",x"66",x"e0",x"c0"),
   830 => (x"ec",x"e8",x"49",x"73"),
   831 => (x"70",x"86",x"c8",x"87"),
   832 => (x"ff",x"c0",x"05",x"98"),
   833 => (x"4a",x"a3",x"dc",x"87"),
   834 => (x"6a",x"49",x"a4",x"c4"),
   835 => (x"4a",x"a3",x"da",x"79"),
   836 => (x"9f",x"49",x"a4",x"c8"),
   837 => (x"79",x"70",x"48",x"6a"),
   838 => (x"c1",x"59",x"a6",x"c4"),
   839 => (x"02",x"bf",x"ec",x"dd"),
   840 => (x"a3",x"d4",x"87",x"d0"),
   841 => (x"49",x"69",x"9f",x"49"),
   842 => (x"ff",x"c0",x"4a",x"71"),
   843 => (x"32",x"d0",x"9a",x"ff"),
   844 => (x"4a",x"c0",x"87",x"c2"),
   845 => (x"bf",x"6e",x"48",x"72"),
   846 => (x"78",x"08",x"6e",x"80"),
   847 => (x"c1",x"7c",x"c0",x"08"),
   848 => (x"87",x"c5",x"c1",x"48"),
   849 => (x"c1",x"48",x"66",x"c8"),
   850 => (x"58",x"a6",x"cc",x"80"),
   851 => (x"c4",x"48",x"66",x"c8"),
   852 => (x"fd",x"04",x"a8",x"66"),
   853 => (x"dd",x"c1",x"87",x"d2"),
   854 => (x"c0",x"02",x"bf",x"ec"),
   855 => (x"49",x"75",x"87",x"e9"),
   856 => (x"70",x"87",x"dd",x"fa"),
   857 => (x"cf",x"49",x"75",x"4d"),
   858 => (x"f8",x"ff",x"ff",x"ff"),
   859 => (x"d6",x"02",x"a9",x"99"),
   860 => (x"c2",x"49",x"75",x"87"),
   861 => (x"e4",x"dd",x"c1",x"89"),
   862 => (x"dd",x"c1",x"91",x"bf"),
   863 => (x"71",x"48",x"bf",x"fc"),
   864 => (x"58",x"a6",x"c4",x"80"),
   865 => (x"c0",x"87",x"d3",x"fc"),
   866 => (x"e7",x"8e",x"f4",x"48"),
   867 => (x"73",x"1e",x"87",x"dd"),
   868 => (x"6a",x"4a",x"71",x"1e"),
   869 => (x"71",x"81",x"c1",x"49"),
   870 => (x"e8",x"dd",x"c1",x"7a"),
   871 => (x"cc",x"05",x"99",x"bf"),
   872 => (x"4b",x"a2",x"c8",x"87"),
   873 => (x"d7",x"f9",x"49",x"6b"),
   874 => (x"71",x"49",x"70",x"87"),
   875 => (x"e6",x"48",x"c1",x"7b"),
   876 => (x"73",x"1e",x"87",x"fd"),
   877 => (x"c1",x"4b",x"71",x"1e"),
   878 => (x"49",x"bf",x"fc",x"dd"),
   879 => (x"6a",x"4a",x"a3",x"c8"),
   880 => (x"c1",x"8a",x"c2",x"4a"),
   881 => (x"92",x"bf",x"e4",x"dd"),
   882 => (x"c1",x"49",x"a1",x"72"),
   883 => (x"4a",x"bf",x"e8",x"dd"),
   884 => (x"a1",x"72",x"9a",x"6b"),
   885 => (x"1e",x"66",x"c8",x"49"),
   886 => (x"fe",x"d5",x"49",x"71"),
   887 => (x"70",x"86",x"c4",x"87"),
   888 => (x"87",x"c4",x"05",x"98"),
   889 => (x"87",x"c2",x"48",x"c0"),
   890 => (x"c2",x"e6",x"48",x"c1"),
   891 => (x"5b",x"5e",x"0e",x"87"),
   892 => (x"71",x"0e",x"5d",x"5c"),
   893 => (x"c1",x"1e",x"73",x"4b"),
   894 => (x"f9",x"49",x"dc",x"de"),
   895 => (x"86",x"c4",x"87",x"ec"),
   896 => (x"c1",x"02",x"98",x"70"),
   897 => (x"de",x"c1",x"87",x"ce"),
   898 => (x"c7",x"49",x"bf",x"e0"),
   899 => (x"29",x"c9",x"81",x"ff"),
   900 => (x"4c",x"c0",x"4d",x"71"),
   901 => (x"49",x"d8",x"ef",x"c0"),
   902 => (x"87",x"c1",x"d5",x"ff"),
   903 => (x"06",x"ad",x"b7",x"c0"),
   904 => (x"d0",x"87",x"c1",x"c1"),
   905 => (x"de",x"c1",x"1e",x"66"),
   906 => (x"c5",x"fe",x"49",x"dc"),
   907 => (x"70",x"86",x"c4",x"87"),
   908 => (x"87",x"c5",x"05",x"98"),
   909 => (x"ed",x"c0",x"48",x"c0"),
   910 => (x"dc",x"de",x"c1",x"87"),
   911 => (x"87",x"ce",x"fd",x"49"),
   912 => (x"c8",x"48",x"66",x"d0"),
   913 => (x"a6",x"d4",x"80",x"c0"),
   914 => (x"75",x"84",x"c1",x"58"),
   915 => (x"ff",x"04",x"ac",x"b7"),
   916 => (x"87",x"d0",x"87",x"d1"),
   917 => (x"ef",x"c0",x"1e",x"73"),
   918 => (x"d3",x"ff",x"1e",x"f1"),
   919 => (x"86",x"c8",x"87",x"d1"),
   920 => (x"87",x"c2",x"48",x"c0"),
   921 => (x"c2",x"e4",x"48",x"c1"),
   922 => (x"86",x"e8",x"1e",x"87"),
   923 => (x"c3",x"4a",x"d4",x"ff"),
   924 => (x"49",x"6a",x"7a",x"ff"),
   925 => (x"6a",x"7a",x"ff",x"c3"),
   926 => (x"c4",x"30",x"c8",x"48"),
   927 => (x"a6",x"c8",x"58",x"a6"),
   928 => (x"c3",x"b1",x"6e",x"59"),
   929 => (x"48",x"6a",x"7a",x"ff"),
   930 => (x"a6",x"cc",x"30",x"d0"),
   931 => (x"59",x"a6",x"d0",x"58"),
   932 => (x"c3",x"b1",x"66",x"c8"),
   933 => (x"48",x"6a",x"7a",x"ff"),
   934 => (x"a6",x"d4",x"30",x"d8"),
   935 => (x"59",x"a6",x"d8",x"58"),
   936 => (x"71",x"b1",x"66",x"d0"),
   937 => (x"26",x"8e",x"e8",x"48"),
   938 => (x"86",x"f4",x"1e",x"4f"),
   939 => (x"c3",x"4a",x"d4",x"ff"),
   940 => (x"49",x"6a",x"7a",x"ff"),
   941 => (x"71",x"7a",x"ff",x"c3"),
   942 => (x"c4",x"30",x"c8",x"48"),
   943 => (x"49",x"6a",x"58",x"a6"),
   944 => (x"ff",x"c3",x"b1",x"6e"),
   945 => (x"c8",x"48",x"71",x"7a"),
   946 => (x"6a",x"58",x"a6",x"30"),
   947 => (x"b1",x"66",x"c4",x"49"),
   948 => (x"71",x"7a",x"ff",x"c3"),
   949 => (x"cc",x"30",x"c8",x"48"),
   950 => (x"49",x"6a",x"58",x"a6"),
   951 => (x"71",x"b1",x"66",x"c8"),
   952 => (x"26",x"8e",x"f4",x"48"),
   953 => (x"5b",x"5e",x"0e",x"4f"),
   954 => (x"71",x"0e",x"5d",x"5c"),
   955 => (x"4c",x"d4",x"ff",x"4d"),
   956 => (x"ff",x"c3",x"48",x"75"),
   957 => (x"c1",x"7c",x"70",x"98"),
   958 => (x"05",x"bf",x"ec",x"de"),
   959 => (x"66",x"d0",x"87",x"c8"),
   960 => (x"d4",x"30",x"c9",x"48"),
   961 => (x"66",x"d0",x"58",x"a6"),
   962 => (x"71",x"29",x"d8",x"49"),
   963 => (x"98",x"ff",x"c3",x"48"),
   964 => (x"66",x"d0",x"7c",x"70"),
   965 => (x"71",x"29",x"d0",x"49"),
   966 => (x"98",x"ff",x"c3",x"48"),
   967 => (x"66",x"d0",x"7c",x"70"),
   968 => (x"71",x"29",x"c8",x"49"),
   969 => (x"98",x"ff",x"c3",x"48"),
   970 => (x"66",x"d0",x"7c",x"70"),
   971 => (x"98",x"ff",x"c3",x"48"),
   972 => (x"49",x"75",x"7c",x"70"),
   973 => (x"48",x"71",x"29",x"d0"),
   974 => (x"70",x"98",x"ff",x"c3"),
   975 => (x"c9",x"4b",x"6c",x"7c"),
   976 => (x"c3",x"4a",x"ff",x"f0"),
   977 => (x"d1",x"05",x"ab",x"ff"),
   978 => (x"49",x"ff",x"c3",x"87"),
   979 => (x"4b",x"6c",x"7c",x"71"),
   980 => (x"c5",x"02",x"8a",x"c1"),
   981 => (x"02",x"ab",x"71",x"87"),
   982 => (x"48",x"73",x"87",x"f2"),
   983 => (x"4c",x"26",x"4d",x"26"),
   984 => (x"4f",x"26",x"4b",x"26"),
   985 => (x"ff",x"49",x"c0",x"1e"),
   986 => (x"ff",x"c3",x"48",x"d4"),
   987 => (x"c3",x"81",x"c1",x"78"),
   988 => (x"04",x"a9",x"b7",x"c8"),
   989 => (x"4f",x"26",x"87",x"f1"),
   990 => (x"5c",x"5b",x"5e",x"0e"),
   991 => (x"ff",x"c0",x"0e",x"5d"),
   992 => (x"4d",x"f7",x"c1",x"f0"),
   993 => (x"c0",x"c0",x"c0",x"c1"),
   994 => (x"ff",x"4b",x"c0",x"c0"),
   995 => (x"f8",x"c4",x"87",x"d6"),
   996 => (x"1e",x"c0",x"4c",x"df"),
   997 => (x"cc",x"fd",x"49",x"75"),
   998 => (x"c1",x"86",x"c4",x"87"),
   999 => (x"e5",x"c0",x"05",x"a8"),
  1000 => (x"48",x"d4",x"ff",x"87"),
  1001 => (x"73",x"78",x"ff",x"c3"),
  1002 => (x"f0",x"e1",x"c0",x"1e"),
  1003 => (x"fc",x"49",x"e9",x"c1"),
  1004 => (x"86",x"c4",x"87",x"f3"),
  1005 => (x"ca",x"05",x"98",x"70"),
  1006 => (x"48",x"d4",x"ff",x"87"),
  1007 => (x"c1",x"78",x"ff",x"c3"),
  1008 => (x"fe",x"87",x"cb",x"48"),
  1009 => (x"8c",x"c1",x"87",x"de"),
  1010 => (x"87",x"c6",x"ff",x"05"),
  1011 => (x"4d",x"26",x"48",x"c0"),
  1012 => (x"4b",x"26",x"4c",x"26"),
  1013 => (x"5e",x"0e",x"4f",x"26"),
  1014 => (x"c0",x"0e",x"5c",x"5b"),
  1015 => (x"c1",x"c1",x"f0",x"ff"),
  1016 => (x"48",x"d4",x"ff",x"4c"),
  1017 => (x"c1",x"78",x"ff",x"c3"),
  1018 => (x"ff",x"49",x"da",x"c0"),
  1019 => (x"d3",x"87",x"ee",x"cd"),
  1020 => (x"74",x"1e",x"c0",x"4b"),
  1021 => (x"87",x"ed",x"fb",x"49"),
  1022 => (x"98",x"70",x"86",x"c4"),
  1023 => (x"ff",x"87",x"ca",x"05"),
  1024 => (x"ff",x"c3",x"48",x"d4"),
  1025 => (x"cb",x"48",x"c1",x"78"),
  1026 => (x"87",x"d8",x"fd",x"87"),
  1027 => (x"ff",x"05",x"8b",x"c1"),
  1028 => (x"48",x"c0",x"87",x"df"),
  1029 => (x"4b",x"26",x"4c",x"26"),
  1030 => (x"4d",x"43",x"4f",x"26"),
  1031 => (x"4d",x"43",x"00",x"44"),
  1032 => (x"20",x"38",x"35",x"44"),
  1033 => (x"20",x"0a",x"64",x"25"),
  1034 => (x"4d",x"43",x"00",x"20"),
  1035 => (x"5f",x"38",x"35",x"44"),
  1036 => (x"64",x"25",x"20",x"32"),
  1037 => (x"00",x"20",x"20",x"0a"),
  1038 => (x"35",x"44",x"4d",x"43"),
  1039 => (x"64",x"25",x"20",x"38"),
  1040 => (x"00",x"20",x"20",x"0a"),
  1041 => (x"43",x"48",x"44",x"53"),
  1042 => (x"69",x"6e",x"49",x"20"),
  1043 => (x"6c",x"61",x"69",x"74"),
  1044 => (x"74",x"61",x"7a",x"69"),
  1045 => (x"20",x"6e",x"6f",x"69"),
  1046 => (x"6f",x"72",x"72",x"65"),
  1047 => (x"00",x"0a",x"21",x"72"),
  1048 => (x"5f",x"64",x"6d",x"63"),
  1049 => (x"38",x"44",x"4d",x"43"),
  1050 => (x"73",x"65",x"72",x"20"),
  1051 => (x"73",x"6e",x"6f",x"70"),
  1052 => (x"25",x"20",x"3a",x"65"),
  1053 => (x"49",x"00",x"0a",x"64"),
  1054 => (x"00",x"52",x"52",x"45"),
  1055 => (x"00",x"49",x"50",x"53"),
  1056 => (x"63",x"20",x"44",x"53"),
  1057 => (x"20",x"64",x"72",x"61"),
  1058 => (x"65",x"7a",x"69",x"73"),
  1059 => (x"20",x"73",x"69",x"20"),
  1060 => (x"00",x"0a",x"64",x"25"),
  1061 => (x"74",x"69",x"72",x"57"),
  1062 => (x"61",x"66",x"20",x"65"),
  1063 => (x"64",x"65",x"6c",x"69"),
  1064 => (x"65",x"52",x"00",x"0a"),
  1065 => (x"63",x"20",x"64",x"61"),
  1066 => (x"61",x"6d",x"6d",x"6f"),
  1067 => (x"66",x"20",x"64",x"6e"),
  1068 => (x"65",x"6c",x"69",x"61"),
  1069 => (x"74",x"61",x"20",x"64"),
  1070 => (x"20",x"64",x"25",x"20"),
  1071 => (x"29",x"64",x"25",x"28"),
  1072 => (x"5f",x"63",x"00",x"0a"),
  1073 => (x"65",x"7a",x"69",x"73"),
  1074 => (x"6c",x"75",x"6d",x"5f"),
  1075 => (x"25",x"20",x"3a",x"74"),
  1076 => (x"72",x"20",x"2c",x"64"),
  1077 => (x"5f",x"64",x"61",x"65"),
  1078 => (x"6c",x"5f",x"6c",x"62"),
  1079 => (x"20",x"3a",x"6e",x"65"),
  1080 => (x"20",x"2c",x"64",x"25"),
  1081 => (x"7a",x"69",x"73",x"63"),
  1082 => (x"25",x"20",x"3a",x"65"),
  1083 => (x"4d",x"00",x"0a",x"64"),
  1084 => (x"20",x"74",x"6c",x"75"),
  1085 => (x"00",x"0a",x"64",x"25"),
  1086 => (x"62",x"20",x"64",x"25"),
  1087 => (x"6b",x"63",x"6f",x"6c"),
  1088 => (x"66",x"6f",x"20",x"73"),
  1089 => (x"7a",x"69",x"73",x"20"),
  1090 => (x"64",x"25",x"20",x"65"),
  1091 => (x"64",x"25",x"00",x"0a"),
  1092 => (x"6f",x"6c",x"62",x"20"),
  1093 => (x"20",x"73",x"6b",x"63"),
  1094 => (x"35",x"20",x"66",x"6f"),
  1095 => (x"62",x"20",x"32",x"31"),
  1096 => (x"73",x"65",x"74",x"79"),
  1097 => (x"5e",x"0e",x"00",x"0a"),
  1098 => (x"0e",x"5d",x"5c",x"5b"),
  1099 => (x"f8",x"4c",x"d4",x"ff"),
  1100 => (x"ea",x"c6",x"87",x"f2"),
  1101 => (x"f0",x"e1",x"c0",x"1e"),
  1102 => (x"f6",x"49",x"c8",x"c1"),
  1103 => (x"4b",x"70",x"87",x"e7"),
  1104 => (x"c1",x"c1",x"1e",x"73"),
  1105 => (x"c7",x"ff",x"1e",x"e0"),
  1106 => (x"86",x"cc",x"87",x"e5"),
  1107 => (x"c8",x"02",x"ab",x"c1"),
  1108 => (x"87",x"c2",x"fa",x"87"),
  1109 => (x"d5",x"c2",x"48",x"c0"),
  1110 => (x"87",x"cd",x"f5",x"87"),
  1111 => (x"ff",x"cf",x"49",x"70"),
  1112 => (x"ea",x"c6",x"99",x"ff"),
  1113 => (x"87",x"c8",x"02",x"a9"),
  1114 => (x"c0",x"87",x"eb",x"f9"),
  1115 => (x"87",x"fe",x"c1",x"48"),
  1116 => (x"c0",x"7c",x"ff",x"c3"),
  1117 => (x"ff",x"f7",x"4d",x"f1"),
  1118 => (x"02",x"98",x"70",x"87"),
  1119 => (x"c0",x"87",x"d4",x"c1"),
  1120 => (x"f0",x"ff",x"c0",x"1e"),
  1121 => (x"f5",x"49",x"fa",x"c1"),
  1122 => (x"86",x"c4",x"87",x"db"),
  1123 => (x"9b",x"73",x"4b",x"70"),
  1124 => (x"87",x"f3",x"c0",x"05"),
  1125 => (x"c0",x"c1",x"1e",x"73"),
  1126 => (x"c6",x"ff",x"1e",x"de"),
  1127 => (x"ff",x"c3",x"87",x"d1"),
  1128 => (x"73",x"4b",x"6c",x"7c"),
  1129 => (x"ea",x"c0",x"c1",x"1e"),
  1130 => (x"c2",x"c6",x"ff",x"1e"),
  1131 => (x"c3",x"86",x"d0",x"87"),
  1132 => (x"7c",x"7c",x"7c",x"ff"),
  1133 => (x"c1",x"49",x"73",x"7c"),
  1134 => (x"c5",x"02",x"99",x"c0"),
  1135 => (x"c0",x"48",x"c1",x"87"),
  1136 => (x"48",x"c0",x"87",x"ec"),
  1137 => (x"73",x"87",x"e7",x"c0"),
  1138 => (x"f8",x"c0",x"c1",x"1e"),
  1139 => (x"de",x"c5",x"ff",x"1e"),
  1140 => (x"c2",x"86",x"c8",x"87"),
  1141 => (x"87",x"ce",x"05",x"ad"),
  1142 => (x"1e",x"c4",x"c1",x"c1"),
  1143 => (x"87",x"cf",x"c5",x"ff"),
  1144 => (x"48",x"c0",x"86",x"c4"),
  1145 => (x"8d",x"c1",x"87",x"c8"),
  1146 => (x"87",x"ca",x"fe",x"05"),
  1147 => (x"4d",x"26",x"48",x"c0"),
  1148 => (x"4b",x"26",x"4c",x"26"),
  1149 => (x"5e",x"0e",x"4f",x"26"),
  1150 => (x"0e",x"5d",x"5c",x"5b"),
  1151 => (x"d0",x"ff",x"86",x"fc"),
  1152 => (x"c0",x"c0",x"c8",x"4c"),
  1153 => (x"ec",x"de",x"c1",x"4b"),
  1154 => (x"c1",x"78",x"c1",x"48"),
  1155 => (x"ff",x"49",x"fc",x"c1"),
  1156 => (x"c7",x"87",x"ca",x"c5"),
  1157 => (x"73",x"48",x"6c",x"4d"),
  1158 => (x"58",x"a6",x"c4",x"98"),
  1159 => (x"87",x"cb",x"02",x"6e"),
  1160 => (x"98",x"73",x"48",x"6c"),
  1161 => (x"6e",x"58",x"a6",x"c4"),
  1162 => (x"c0",x"87",x"f5",x"05"),
  1163 => (x"87",x"f4",x"f4",x"7c"),
  1164 => (x"98",x"73",x"48",x"6c"),
  1165 => (x"6e",x"58",x"a6",x"c4"),
  1166 => (x"6c",x"87",x"cb",x"02"),
  1167 => (x"c4",x"98",x"73",x"48"),
  1168 => (x"05",x"6e",x"58",x"a6"),
  1169 => (x"7c",x"c1",x"87",x"f5"),
  1170 => (x"e5",x"c0",x"1e",x"c0"),
  1171 => (x"49",x"c0",x"c1",x"d0"),
  1172 => (x"c4",x"87",x"d2",x"f2"),
  1173 => (x"05",x"a8",x"c1",x"86"),
  1174 => (x"4d",x"c1",x"87",x"c2"),
  1175 => (x"cd",x"05",x"ad",x"c2"),
  1176 => (x"f7",x"c1",x"c1",x"87"),
  1177 => (x"f4",x"c3",x"ff",x"49"),
  1178 => (x"c1",x"48",x"c0",x"87"),
  1179 => (x"8d",x"c1",x"87",x"de"),
  1180 => (x"87",x"e1",x"fe",x"05"),
  1181 => (x"c1",x"87",x"ef",x"fa"),
  1182 => (x"c1",x"58",x"f0",x"de"),
  1183 => (x"05",x"bf",x"ec",x"de"),
  1184 => (x"1e",x"c1",x"87",x"cd"),
  1185 => (x"c1",x"f0",x"ff",x"c0"),
  1186 => (x"d8",x"f1",x"49",x"d0"),
  1187 => (x"ff",x"86",x"c4",x"87"),
  1188 => (x"ff",x"c3",x"48",x"d4"),
  1189 => (x"87",x"d6",x"c5",x"78"),
  1190 => (x"58",x"f4",x"de",x"c1"),
  1191 => (x"bf",x"f0",x"de",x"c1"),
  1192 => (x"c0",x"c2",x"c1",x"1e"),
  1193 => (x"c6",x"c2",x"ff",x"1e"),
  1194 => (x"6c",x"86",x"c8",x"87"),
  1195 => (x"c4",x"98",x"73",x"48"),
  1196 => (x"02",x"6e",x"58",x"a6"),
  1197 => (x"48",x"6c",x"87",x"cc"),
  1198 => (x"a6",x"c4",x"98",x"73"),
  1199 => (x"ff",x"05",x"6e",x"58"),
  1200 => (x"7c",x"c0",x"87",x"f4"),
  1201 => (x"c3",x"48",x"d4",x"ff"),
  1202 => (x"48",x"c1",x"78",x"ff"),
  1203 => (x"4d",x"26",x"8e",x"fc"),
  1204 => (x"4b",x"26",x"4c",x"26"),
  1205 => (x"5e",x"0e",x"4f",x"26"),
  1206 => (x"0e",x"5d",x"5c",x"5b"),
  1207 => (x"d4",x"ff",x"4b",x"71"),
  1208 => (x"4c",x"66",x"d0",x"4d"),
  1209 => (x"ee",x"c5",x"4a",x"c0"),
  1210 => (x"c3",x"49",x"df",x"cd"),
  1211 => (x"48",x"6d",x"7d",x"ff"),
  1212 => (x"05",x"a8",x"fe",x"c3"),
  1213 => (x"c1",x"87",x"d1",x"c1"),
  1214 => (x"c0",x"48",x"e8",x"de"),
  1215 => (x"ac",x"b7",x"c4",x"78"),
  1216 => (x"ed",x"87",x"db",x"04"),
  1217 => (x"49",x"70",x"87",x"e3"),
  1218 => (x"83",x"c4",x"7b",x"71"),
  1219 => (x"bf",x"e8",x"de",x"c1"),
  1220 => (x"c1",x"80",x"71",x"48"),
  1221 => (x"c4",x"58",x"ec",x"de"),
  1222 => (x"03",x"ac",x"b7",x"8c"),
  1223 => (x"b7",x"c0",x"87",x"e5"),
  1224 => (x"e0",x"c0",x"06",x"ac"),
  1225 => (x"7d",x"ff",x"c3",x"87"),
  1226 => (x"09",x"73",x"49",x"6d"),
  1227 => (x"c1",x"09",x"79",x"97"),
  1228 => (x"e8",x"de",x"c1",x"83"),
  1229 => (x"80",x"71",x"48",x"bf"),
  1230 => (x"58",x"ec",x"de",x"c1"),
  1231 => (x"b7",x"c0",x"8c",x"c1"),
  1232 => (x"e0",x"ff",x"01",x"ac"),
  1233 => (x"4a",x"49",x"c1",x"87"),
  1234 => (x"fe",x"05",x"89",x"c1"),
  1235 => (x"ff",x"c3",x"87",x"dd"),
  1236 => (x"26",x"48",x"72",x"7d"),
  1237 => (x"26",x"4c",x"26",x"4d"),
  1238 => (x"0e",x"4f",x"26",x"4b"),
  1239 => (x"5d",x"5c",x"5b",x"5e"),
  1240 => (x"71",x"86",x"f8",x"0e"),
  1241 => (x"4c",x"d0",x"ff",x"4d"),
  1242 => (x"4b",x"c0",x"c0",x"c8"),
  1243 => (x"d4",x"ff",x"7e",x"c0"),
  1244 => (x"78",x"ff",x"c3",x"48"),
  1245 => (x"98",x"73",x"48",x"6c"),
  1246 => (x"c4",x"58",x"a6",x"c8"),
  1247 => (x"87",x"cc",x"02",x"66"),
  1248 => (x"98",x"73",x"48",x"6c"),
  1249 => (x"c4",x"58",x"a6",x"c8"),
  1250 => (x"87",x"f4",x"05",x"66"),
  1251 => (x"ff",x"7c",x"c1",x"c4"),
  1252 => (x"ff",x"c3",x"48",x"d4"),
  1253 => (x"c0",x"1e",x"75",x"78"),
  1254 => (x"d1",x"c1",x"f0",x"ff"),
  1255 => (x"87",x"c5",x"ed",x"49"),
  1256 => (x"4a",x"70",x"86",x"c4"),
  1257 => (x"d1",x"02",x"9a",x"72"),
  1258 => (x"75",x"1e",x"72",x"87"),
  1259 => (x"e2",x"c2",x"c1",x"1e"),
  1260 => (x"fa",x"fd",x"fe",x"1e"),
  1261 => (x"c0",x"86",x"cc",x"87"),
  1262 => (x"c0",x"c8",x"87",x"e8"),
  1263 => (x"49",x"66",x"dc",x"1e"),
  1264 => (x"c4",x"87",x"d3",x"fc"),
  1265 => (x"58",x"a6",x"c4",x"86"),
  1266 => (x"98",x"73",x"48",x"6c"),
  1267 => (x"c4",x"58",x"a6",x"c8"),
  1268 => (x"87",x"cc",x"02",x"66"),
  1269 => (x"98",x"73",x"48",x"6c"),
  1270 => (x"c4",x"58",x"a6",x"c8"),
  1271 => (x"87",x"f4",x"05",x"66"),
  1272 => (x"48",x"6e",x"7c",x"c0"),
  1273 => (x"4d",x"26",x"8e",x"f8"),
  1274 => (x"4b",x"26",x"4c",x"26"),
  1275 => (x"5e",x"0e",x"4f",x"26"),
  1276 => (x"0e",x"5d",x"5c",x"5b"),
  1277 => (x"1e",x"c0",x"86",x"fc"),
  1278 => (x"c1",x"f0",x"ff",x"c0"),
  1279 => (x"e4",x"eb",x"49",x"c9"),
  1280 => (x"c1",x"1e",x"d2",x"87"),
  1281 => (x"fb",x"49",x"fa",x"de"),
  1282 => (x"86",x"c8",x"87",x"cc"),
  1283 => (x"85",x"c1",x"4d",x"c0"),
  1284 => (x"04",x"ad",x"b7",x"d2"),
  1285 => (x"de",x"c1",x"87",x"f8"),
  1286 => (x"49",x"bf",x"97",x"fa"),
  1287 => (x"c1",x"99",x"c0",x"c3"),
  1288 => (x"c0",x"05",x"a9",x"c0"),
  1289 => (x"df",x"c1",x"87",x"e8"),
  1290 => (x"49",x"bf",x"97",x"c1"),
  1291 => (x"df",x"c1",x"31",x"d0"),
  1292 => (x"4a",x"bf",x"97",x"c2"),
  1293 => (x"b1",x"72",x"32",x"c8"),
  1294 => (x"97",x"c3",x"df",x"c1"),
  1295 => (x"b1",x"72",x"4a",x"bf"),
  1296 => (x"ff",x"cf",x"4d",x"71"),
  1297 => (x"c1",x"9d",x"ff",x"ff"),
  1298 => (x"c2",x"35",x"ca",x"85"),
  1299 => (x"df",x"c1",x"87",x"e6"),
  1300 => (x"4b",x"bf",x"97",x"c3"),
  1301 => (x"9b",x"c6",x"33",x"c1"),
  1302 => (x"97",x"c4",x"df",x"c1"),
  1303 => (x"b7",x"c7",x"49",x"bf"),
  1304 => (x"c1",x"b3",x"71",x"29"),
  1305 => (x"bf",x"97",x"ff",x"de"),
  1306 => (x"cf",x"48",x"71",x"49"),
  1307 => (x"58",x"a6",x"c4",x"98"),
  1308 => (x"97",x"c0",x"df",x"c1"),
  1309 => (x"9c",x"c3",x"4c",x"bf"),
  1310 => (x"df",x"c1",x"34",x"ca"),
  1311 => (x"49",x"bf",x"97",x"c1"),
  1312 => (x"b4",x"71",x"31",x"c2"),
  1313 => (x"97",x"c2",x"df",x"c1"),
  1314 => (x"c0",x"c3",x"49",x"bf"),
  1315 => (x"29",x"b7",x"c6",x"99"),
  1316 => (x"1e",x"74",x"b4",x"71"),
  1317 => (x"73",x"1e",x"66",x"c4"),
  1318 => (x"c2",x"c3",x"c1",x"1e"),
  1319 => (x"ce",x"fa",x"fe",x"1e"),
  1320 => (x"c1",x"83",x"c2",x"87"),
  1321 => (x"70",x"30",x"73",x"48"),
  1322 => (x"c1",x"1e",x"73",x"4b"),
  1323 => (x"fe",x"1e",x"ef",x"c3"),
  1324 => (x"c1",x"87",x"fc",x"f9"),
  1325 => (x"30",x"66",x"d8",x"48"),
  1326 => (x"c1",x"58",x"a6",x"dc"),
  1327 => (x"73",x"4d",x"49",x"a4"),
  1328 => (x"1e",x"66",x"d8",x"95"),
  1329 => (x"c3",x"c1",x"1e",x"75"),
  1330 => (x"f9",x"fe",x"1e",x"f8"),
  1331 => (x"e4",x"c0",x"87",x"e1"),
  1332 => (x"c8",x"48",x"6e",x"86"),
  1333 => (x"06",x"a8",x"b7",x"c0"),
  1334 => (x"4b",x"6e",x"87",x"ce"),
  1335 => (x"2b",x"b7",x"35",x"c1"),
  1336 => (x"ab",x"b7",x"c0",x"c8"),
  1337 => (x"87",x"f4",x"ff",x"01"),
  1338 => (x"c4",x"c1",x"1e",x"75"),
  1339 => (x"f8",x"fe",x"1e",x"ce"),
  1340 => (x"86",x"c8",x"87",x"fd"),
  1341 => (x"8e",x"fc",x"48",x"75"),
  1342 => (x"4c",x"26",x"4d",x"26"),
  1343 => (x"4f",x"26",x"4b",x"26"),
  1344 => (x"71",x"1e",x"73",x"1e"),
  1345 => (x"d8",x"49",x"73",x"4b"),
  1346 => (x"99",x"ff",x"c3",x"29"),
  1347 => (x"2a",x"c8",x"4a",x"73"),
  1348 => (x"9a",x"c0",x"fc",x"cf"),
  1349 => (x"4a",x"73",x"b1",x"72"),
  1350 => (x"ff",x"c0",x"32",x"c8"),
  1351 => (x"9a",x"c0",x"c0",x"f0"),
  1352 => (x"4a",x"73",x"b1",x"72"),
  1353 => (x"c0",x"ff",x"32",x"d8"),
  1354 => (x"9a",x"c0",x"c0",x"c0"),
  1355 => (x"48",x"71",x"b1",x"72"),
  1356 => (x"4f",x"26",x"4b",x"26"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
