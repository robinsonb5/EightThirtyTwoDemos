library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;
use work.DMACache_pkg.ALL;
use work.DMACache_config.ALL;
use work.SoC_Peripheral_config.all;
use work.SoC_Peripheral_pkg.all;


entity VirtualToplevel is
	generic (
		sdram_rows : integer := 12;
		sdram_cols : integer := 8;
		sysclk_frequency : integer := 1000; -- Sysclk frequency * 10
		jtag_uart : boolean := false;
		debug : boolean := false
	);
	port (
		clk 			: in std_logic;
		slowclk		: in std_logic;
		videoclk	: in std_logic;
		reset_in 	: in std_logic;

		-- VGA
		vga_red 		: out unsigned(7 downto 0);
		vga_green 	: out unsigned(7 downto 0);
		vga_blue 	: out unsigned(7 downto 0);
		vga_hsync 	: out std_logic;
		vga_vsync 	: buffer std_logic;
		vga_window	: out std_logic;
		vga_pixel	: out std_logic;

		-- SDRAM
		sdr_drive_data  : out std_logic;
		sdr_data_in		: in std_logic_vector(31 downto 0) := (others => '0');
		sdr_data_out	: inout std_logic_vector(31 downto 0);
		sdr_addr		: out std_logic_vector((sdram_rows-1) downto 0);
		sdr_dqm 		: out std_logic_vector(3 downto 0);
		sdr_we 		: out std_logic;
		sdr_cas 		: out std_logic;
		sdr_ras 		: out std_logic;
		sdr_cs		: out std_logic;
		sdr_ba		: out std_logic_vector(1 downto 0);
--		sdr_clk		: out std_logic;
		sdr_cke		: out std_logic;

		-- SPI signals
		spi_miso		: in std_logic := '1'; -- Allow the SPI interface not to be plumbed in.
		spi_mosi		: out std_logic;
		spi_clk		: out std_logic;
		spi_cs 		: out std_logic;
		
		-- PS/2 signals
		ps2k_clk_in : in std_logic := '1';
		ps2k_dat_in : in std_logic := '1';
		ps2k_clk_out : out std_logic;
		ps2k_dat_out : out std_logic;
		ps2m_clk_in : in std_logic := '1';
		ps2m_dat_in : in std_logic := '1';
		ps2m_clk_out : out std_logic;
		ps2m_dat_out : out std_logic;

		-- UARTs
		rxd	: in std_logic := '1';
		txd	: out std_logic;
		rxd2	: in std_logic := '1';
		txd2	: out std_logic;
		
		-- Audio
		AUDIO_L : out signed(15 downto 0);
		AUDIO_R : out signed(15 downto 0)
);
end entity;

architecture rtl of VirtualToplevel is

	constant Peripheral_Blocks : integer := 4;

	component debug_bridge_jtag is
	generic (
		id : natural := 16#832D#
	);
	port (
		clk : in std_logic;
		reset_n : in std_logic;
		d : in std_logic_vector(31 downto 0);
		q : out std_logic_vector(31 downto 0);
		req : in std_logic;
		wr : in std_logic;
		ack : buffer std_logic
	);
	end component;

	constant sysclk_hz : integer := sysclk_frequency*1000;
	constant maxAddrBit : integer := 31;

	signal reset_n : std_logic := '0';
	signal reset : std_logic := '0';
	signal reset_counter : unsigned(15 downto 0) := X"FFFF";

	-- Interrupt signals

	constant int_max : integer := 2;
	signal int_triggers : std_logic_vector(int_max downto 0);

	-- Timer register block signals

	signal timer_reg_req : std_logic;
	signal timer_tick : std_logic;


	-- Plumbing between DMA controller and SDRAM

	signal video_addr : std_logic_vector(31 downto 0);
	signal video_data_in : std_logic_vector(31 downto 0);
	signal video_req : std_logic;
	signal video_pri : std_logic;
	signal video_ack : std_logic;
	signal video_fill : std_logic;

	signal dma_addr : std_logic_vector(31 downto 0);
	signal dma_data_in : std_logic_vector(31 downto 0);
	signal dma_req : std_logic;
	signal dma_ack : std_logic;
	signal dma_fill : std_logic;

	signal dma_data : std_logic_vector(31 downto 0);

	-- Plumbing between VGA controller and DMA controller

	signal vgachannel_fromhost : DMAChannel_FromHost;
	signal vgachannel_tohost : DMAChannel_ToHost;
	signal spr0channel_fromhost : DMAChannel_FromHost;
	signal spr0channel_tohost : DMAChannel_ToHost;

	-- Audio channel plumbing

	signal aud0_fromhost : DMAChannel_FromHost;
	signal aud0_tohost : DMAChannel_ToHost;
	signal aud1_fromhost : DMAChannel_FromHost;
	signal aud1_tohost : DMAChannel_ToHost;
	signal aud2_fromhost : DMAChannel_FromHost;
	signal aud2_tohost : DMAChannel_ToHost;
	signal aud3_fromhost : DMAChannel_FromHost;
	signal aud3_tohost : DMAChannel_ToHost;

	signal audio_reg_req : std_logic;
	signal audio_ints : std_logic_vector(3 downto 0);
	signal audio_int : std_logic;
	
	signal audio_l_i : signed(23 downto 0);
	signal audio_r_i : signed(23 downto 0);

	-- VGA register block signals

	signal vga_reg_addr : std_logic_vector(11 downto 0);
	signal vga_reg_dataout : std_logic_vector(15 downto 0);
	signal vga_reg_datain : std_logic_vector(15 downto 0);
	signal vga_reg_rw : std_logic;
	signal vga_reg_req : std_logic;
	signal vga_reg_dtack : std_logic;
	signal vga_ack : std_logic;
	signal vblank_int : std_logic;
	signal vga_vsync_i : std_logic;


	-- SDRAM signals

	signal sdr_ready : std_logic;
	signal sdram_write : std_logic_vector(31 downto 0); -- 32-bit width for ZPU
	signal sdram_req : std_logic;
	signal sdram_wr : std_logic;
	signal sdram_read : std_logic_vector(31 downto 0);
	signal sdram_ack : std_logic;
	signal sdram_bytesel : std_logic_vector(3 downto 0);

	type sdram_states is (idle, waiting, pause);
	signal sdram_state : sdram_states;


	-- CPU signals
	signal cpu_reset : std_logic;
	signal cpu_int : std_logic;
	signal soft_reset_n : std_logic;
	
	signal mem_peripherals : std_logic;
	signal peripherals_ack : std_logic;
	signal from_peripherals : std_logic_vector(31 downto 0);

	signal mem_ram : std_logic;
	signal ram_ack : std_logic;
	signal from_ram : std_logic_vector(31 downto 0);

	signal mem_rom : std_logic;
	signal rom_ack : std_logic;
	signal from_rom : std_logic_vector(31 downto 0);

	signal cpu_addr : std_logic_vector(31 downto 0);
	signal to_cpu : std_logic_vector(31 downto 0);
	signal from_cpu : std_logic_vector(31 downto 0);
	signal cpu_req : std_logic; 
	signal cpu_ack : std_logic; 
	signal cpu_wr : std_logic; 
	signal cpu_bytesel : std_logic_vector(3 downto 0);
	signal bytesel_rev : std_logic_vector(3 downto 0);
	signal cache_valid : std_logic;
	signal flushcaches : std_logic;

	-- CPU Debug signals
	signal debug_req : std_logic;
	signal debug_ack : std_logic;
	signal debug_fromcpu : std_logic_vector(31 downto 0);
	signal debug_tocpu : std_logic_vector(31 downto 0);
	signal debug_wr : std_logic;

	signal peripheral_block : std_logic_vector(3 downto 0);

begin

	sdr_cke <='1';

	-- Reset counter.

	process(clk,reset_in,sdr_ready)
	begin
		if reset_in='0' or sdr_ready='0' then
			reset_counter<=X"FFFF";
			reset_n<='0';
		elsif rising_edge(clk) then
			reset_counter<=reset_counter-1;
			if reset_counter=X"0000" then
				reset_n<='1';
			end if;
		end if;
	end process;

	reset <= not reset_n;

	
	-- SDRAM
	bytesel_rev <= cpu_bytesel(0)&cpu_bytesel(1)&cpu_bytesel(2)&cpu_bytesel(3);

	mysdram : entity work.sdram_cached_wide
		generic map
		(
			rows => sdram_rows,
			cols => sdram_cols,
			cache => true,
			dqwidth => 32,
			dqmwidth => 4
		)
		port map
		(
		-- Physical connections to the SDRAM
			drive_sdata => sdr_drive_data,
			sdata_in => sdr_data_in,
			sdata_out => sdr_data_out,
			sdaddr => sdr_addr,
			sd_we	=> sdr_we,
			sd_ras => sdr_ras,
			sd_cas => sdr_cas,
			sd_cs	=> sdr_cs,
			dqm => sdr_dqm,
			ba	=> sdr_ba,

		-- Housekeeping
			sysclk => clk,
			reset => reset_in,  -- Contributes to reset, so have to use reset_in here.
			reset_out => sdr_ready,

			vga_addr => video_addr,
			vga_data => video_data_in,
			vga_fill => video_fill,
			vga_req => video_req,
			vga_pri => video_pri,
			vga_ack => video_ack,

			datawr1(31 downto 24) => sdram_write(7 downto 0),
			datawr1(23 downto 16) => sdram_write(15 downto 8),
			datawr1(15 downto 8) => sdram_write(23 downto 16),
			datawr1(7 downto 0) => sdram_write(31 downto 24),
			addr1 => cpu_addr,
			req1 => sdram_req,
			cachevalid => cache_valid,
			wr1 => sdram_wr, -- active low
			bytesel => sdram_bytesel, -- cpu_bytesel,
			dataout1 => sdram_read,
			ack1 => sdram_ack,

			addr2 => dma_addr,
			dataout2 => dma_data_in,
			fill2 => dma_fill,
			req2 => dma_req,
			ack2 => dma_ack,
			
			flushcaches => flushcaches
		);

-- DMA controller

	mydmacache : entity work.DMACache
		port map(
			clk => clk,
			reset_n => cpu_reset,

--			channels_from_host(0) => vgachannel_fromhost,
			channels_from_host(0) => spr0channel_fromhost,
			channels_from_host(1) => aud0_fromhost,
			channels_from_host(2) => aud1_fromhost,
			channels_from_host(3) => aud2_fromhost,
			channels_from_host(4) => aud3_fromhost,

--			channels_to_host(0) => vgachannel_tohost,
			channels_to_host(0) => spr0channel_tohost,
			channels_to_host(1) => aud0_tohost,
			channels_to_host(2) => aud1_tohost,
			channels_to_host(3) => aud2_tohost,
			channels_to_host(4) => aud3_tohost,

			data_out => dma_data,

			-- SDRAM interface
			sdram_addr=> dma_addr,
			sdram_req => dma_req,
			sdram_ack => dma_ack,
			sdram_fill => dma_fill,
			sdram_data => dma_data_in
		);


	-- Main CPU

	mem_peripherals <= '1' when cpu_addr(31)='1' else '0';
	mem_rom <='1' when cpu_addr(31 downto 26)=X"0"&"00" else '0';
	mem_ram <='1' when mem_peripherals='0' and mem_rom='0' else '0';
		
	process(clk)
	begin
		if rising_edge(clk) then

			if mem_rom='1' then
				to_cpu<=from_rom;
			elsif mem_peripherals='1' then
				to_cpu<=from_peripherals;
			else
				to_cpu<=from_ram;
			end if;

			if (ram_ack='1' or rom_ack='1' or peripherals_ack='1') and cpu_ack='0' then
				cpu_ack<='1';
			else
				cpu_ack<='0';
			end if;
	
		end if;	
	end process;
	
	cpu_reset<=reset_n and soft_reset_n;
	
	cpu : entity work.eightthirtytwo_cpu
	generic map
	(
		multiplier => true,
		littleendian => true,
		dualthread => true,
		prefetch => true,
		interrupts => true,
		debug => debug
	)
	port map
	(
		clk => clk,
		reset_n => cpu_reset,
		interrupt => cpu_int,

		-- cpu fetch interface

		addr => cpu_addr(31 downto 2),
		d => to_cpu,
		q => from_cpu,
		bytesel => cpu_bytesel,
		wr => cpu_wr,
		req => cpu_req,
		ack => cpu_ack,
		-- Debug signals
		debug_d=>debug_tocpu,
		debug_q=>debug_fromcpu,
		debug_req=>debug_req,
		debug_wr=>debug_wr,
		debug_ack=>debug_ack		
	);
	cpu_addr(1 downto 0) <= (others => '0'); -- Ensure the low order bits are clear
	
	gendebug:
	if debug = true generate
		debugbridge : component debug_bridge_jtag
		port map
		(
			clk => slowclk,
			reset_n => reset_n,
			d => debug_fromcpu,
			q => debug_tocpu,
			req => debug_req,
			ack => debug_ack,
			wr => debug_wr
		);
	end generate;

	gennodebug:
	if debug = false generate
		debug_ack <= '0';
	end generate;


	-- Standard peripheral block
	peripheralblock : block
		signal peripheral_req : SoC_Peripheral_Request;
		type responses_t is array (0 to Peripheral_Blocks-1) of SoC_Peripheral_Response;
		signal peripheral_responses : responses_t;
	begin

		audio_int <= '0' when audio_ints="0000" else '1';
		int_triggers<=(0=>timer_tick, 1=>vblank_int, 2=>audio_int, others => '0');

		standardperipherals : entity work.Peripheral_Standard
			generic map (
				BlockAddress => X"F",
				sysclk_frequency => sysclk_frequency,
				external_interrupts => 3
			)
			port map (
				clk => clk,
				reset_n => cpu_reset,
				request => peripheral_req,
				response => peripheral_responses(0),

				-- CPU / system signals		
				soft_reset_n => soft_reset_n,
				flush_caches => flushcaches,

				-- Interupt signals
				interrupt_triggers => int_triggers,
				interrupt => cpu_int,

				-- SPI signals
				spi_miso => spi_miso,
				spi_mosi => spi_mosi,
				spi_clk => spi_clk,
				spi_cs => spi_cs,
				
				-- PS/2 signals
				ps2k_clk_in => ps2k_clk_in,
				ps2k_dat_in => ps2k_dat_in,
				ps2k_clk_out => ps2k_clk_out,
				ps2k_dat_out => ps2k_dat_out,
				ps2m_clk_in => ps2m_clk_in,
				ps2m_dat_in => ps2m_dat_in,
				ps2m_clk_out => ps2m_clk_out,
				ps2m_dat_out => ps2m_dat_out,

				-- UARTs
				rxd => rxd,
				txd => txd,
				rxd2 => rxd2,
				txd2 => txd2
			);

		-- Video
		
		video : entity work.vga_controller_new
			generic map (
				BlockAddress => X"E",
				dmawidth => 32
			)
			port map (
			clk_sys => clk,
			reset_n => reset_in,

			request => peripheral_req,
			response => peripheral_responses(1),

			-- Sprite
			sprite0_sys => spr0channel_fromhost,
			sprite0_status => spr0channel_tohost,
			spritedata => dma_data,

			-- Video
			
			clk_video => videoclk,
			video_req => video_req,
			video_pri => video_pri,
			video_ack => video_ack,
			video_fill => video_fill,
			video_addr => video_addr,
			video_data_in => video_data_in,		

			vblank_int => vblank_int,
			hsync => vga_hsync,
			vsync => vga_vsync_i,
			red => vga_red,
			green => vga_green,
			blue => vga_blue,
			vga_window => vga_window,
			vga_pixel => vga_pixel
		);

		vga_vsync<=vga_vsync_i;


		-- Audio controller
			
		audio : entity work.sound_wrapper_new
			generic map(
				BlockAddress => X"D",
				dmawidth => 32,
				clk_frequency => sysclk_frequency -- Prescale incoming clock
			)
		port map (
			clk => clk,
			reset => cpu_reset,

			request => peripheral_req,
			response => peripheral_responses(2),

			dma_data => dma_data,
			channel0_fromhost => aud0_fromhost,
			channel0_tohost => aud0_tohost,
			channel1_fromhost => aud1_fromhost,
			channel1_tohost => aud1_tohost,
			channel2_fromhost => aud2_fromhost,
			channel2_tohost => aud2_tohost,
			channel3_fromhost => aud3_fromhost,
			channel3_tohost => aud3_tohost,

			audio_l => audio_l_i,
			audio_r => audio_r_i,
			audio_ints => audio_ints
		);

		audio_l<=audio_l_i(23 downto 8);
		audio_r<=audio_r_i(23 downto 8);

		-- Timer
			
		timer : entity work.timer_controller_new
		generic map(
			BlockAddress => X"C",
			prescale => sysclk_frequency, -- Prescale incoming clock
			timers => 0
		)
		port map (
			clk => clk,
			reset => reset_n,

			request => peripheral_req,
			response => peripheral_responses(3),

			ticks(0) => timer_tick -- Tick signal is used to trigger an interrupt
		);

		
		-- Peripherals

		process(clk,reset_n) begin
			if rising_edge(clk) then
				
				peripheral_req.addr<=cpu_addr;
				peripheral_req.wr<=cpu_wr;
				peripheral_req.d<=from_cpu;
				peripheral_req.req<=mem_peripherals and cpu_req;

				peripherals_ack<='0';
				for I in 0 to Peripheral_Blocks-1 loop
					if peripheral_responses(I).ack='1' then
						peripherals_ack<='1';
						from_peripherals<=peripheral_responses(i).q;
					end if;
				end loop;
			end if;
		end process;
	end block;
	
	-- SDRAM state machine
	
	-- Combinational to take effect one cycle sooner.
	ram_ack <= '1' when sdram_state=waiting and (sdram_ack='1' or cache_valid='1') else '0';
	-- Endian byte mangling
	from_ram(7 downto 0)<=sdram_read(31 downto 24);
	from_ram(15 downto 8)<=sdram_read(23 downto 16);
	from_ram(23 downto 16)<=sdram_read(15 downto 8);
	from_ram(31 downto 24)<=sdram_read(7 downto 0);

	process(clk,reset_n) begin
		if reset_n='0' then
			sdram_state<=idle;
		elsif rising_edge(clk) then

			case sdram_state is
				when idle =>
					if cpu_req='1' and mem_ram='1' then
						sdram_bytesel<=bytesel_rev;
						sdram_wr<=cpu_wr;
						sdram_req<='1';
						sdram_write<=from_cpu;
						sdram_state<=waiting;
					end if;

				when waiting =>	
					if sdram_ack='1' or cache_valid='1' then
						sdram_req<='0';
						sdram_state<=pause;
					end if;

				when pause =>
					sdram_state<=idle;

				when others =>
					null;
			end case;

		end if; -- rising-edge(clk)

	end process;

	-- ROM

	romblock : block
		signal rom_wr : std_logic;
	begin
		process(clk) begin
			if rising_edge(clk) then
				if mem_rom='1' then
					rom_wr<=(cpu_wr and cpu_req);
				else
					rom_wr<='0';
				end if;
				rom_ack<=cpu_req and mem_rom;
			end if;
		end process;

		-- ROM

		rom : entity work.SoCWide_rom
		generic map(
			ADDR_WIDTH => 13
		)
		port map(
			clk => clk,		
			addr => cpu_addr(14 downto 2),
			d => from_cpu,
			q => from_rom,
			we => rom_wr,
			bytesel => cpu_bytesel
		);
		
	end block;

end architecture;
