
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"44",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"36"),
    10 => (x"c0",x"c0",x"c2",x"4f"),
    11 => (x"15",x"0c",x"27",x"4e"),
    12 => (x"00",x"0f",x"00",x"00"),
    13 => (x"f0",x"c1",x"87",x"fd"),
    14 => (x"43",x"27",x"4e",x"c0"),
    15 => (x"0f",x"00",x"00",x"00"),
    16 => (x"4f",x"87",x"fd",x"00"),
    17 => (x"ff",x"1e",x"1e",x"4f"),
    18 => (x"48",x"69",x"49",x"c0"),
    19 => (x"c4",x"98",x"c0",x"c4"),
    20 => (x"02",x"6e",x"58",x"a6"),
    21 => (x"c8",x"87",x"f3",x"ff"),
    22 => (x"26",x"48",x"79",x"66"),
    23 => (x"87",x"c6",x"c0",x"c0"),
    24 => (x"4c",x"26",x"4d",x"26"),
    25 => (x"4f",x"26",x"4b",x"26"),
    26 => (x"5c",x"5b",x"5e",x"0e"),
    27 => (x"4c",x"66",x"cc",x"0e"),
    28 => (x"4a",x"14",x"4b",x"c0"),
    29 => (x"72",x"9a",x"ff",x"c3"),
    30 => (x"d9",x"c0",x"02",x"9a"),
    31 => (x"71",x"49",x"72",x"87"),
    32 => (x"00",x"45",x"27",x"1e"),
    33 => (x"c4",x"0f",x"00",x"00"),
    34 => (x"14",x"83",x"c1",x"86"),
    35 => (x"9a",x"ff",x"c3",x"4a"),
    36 => (x"ff",x"05",x"9a",x"72"),
    37 => (x"48",x"73",x"87",x"e7"),
    38 => (x"87",x"c6",x"ff",x"ff"),
    39 => (x"5c",x"5b",x"5e",x"0e"),
    40 => (x"86",x"f0",x"0e",x"5d"),
    41 => (x"a6",x"c4",x"4b",x"c0"),
    42 => (x"c0",x"78",x"c0",x"48"),
    43 => (x"c0",x"4c",x"a6",x"e4"),
    44 => (x"48",x"49",x"66",x"e0"),
    45 => (x"e4",x"c0",x"80",x"c1"),
    46 => (x"4a",x"11",x"58",x"a6"),
    47 => (x"ba",x"82",x"c0",x"fe"),
    48 => (x"c4",x"02",x"9a",x"72"),
    49 => (x"66",x"c4",x"87",x"ef"),
    50 => (x"87",x"f9",x"c3",x"02"),
    51 => (x"c0",x"48",x"a6",x"c4"),
    52 => (x"c0",x"49",x"72",x"78"),
    53 => (x"c3",x"02",x"aa",x"f0"),
    54 => (x"e3",x"c1",x"87",x"c1"),
    55 => (x"c2",x"c3",x"02",x"a9"),
    56 => (x"a9",x"e4",x"c1",x"87"),
    57 => (x"87",x"e3",x"c0",x"02"),
    58 => (x"02",x"a9",x"ec",x"c1"),
    59 => (x"c1",x"87",x"ec",x"c2"),
    60 => (x"c0",x"02",x"a9",x"f0"),
    61 => (x"f3",x"c1",x"87",x"d5"),
    62 => (x"c7",x"c2",x"02",x"a9"),
    63 => (x"a9",x"f5",x"c1",x"87"),
    64 => (x"87",x"c7",x"c0",x"02"),
    65 => (x"05",x"a9",x"f8",x"c1"),
    66 => (x"c4",x"87",x"ed",x"c2"),
    67 => (x"c4",x"49",x"74",x"84"),
    68 => (x"69",x"48",x"76",x"89"),
    69 => (x"c1",x"02",x"6e",x"78"),
    70 => (x"80",x"c8",x"87",x"da"),
    71 => (x"a6",x"cc",x"78",x"c0"),
    72 => (x"6e",x"78",x"c0",x"48"),
    73 => (x"29",x"b7",x"dc",x"49"),
    74 => (x"9a",x"cf",x"4a",x"71"),
    75 => (x"30",x"c4",x"48",x"6e"),
    76 => (x"72",x"58",x"a6",x"c4"),
    77 => (x"c5",x"c0",x"02",x"9a"),
    78 => (x"48",x"a6",x"c8",x"87"),
    79 => (x"aa",x"c9",x"78",x"c1"),
    80 => (x"87",x"c6",x"c0",x"06"),
    81 => (x"c0",x"82",x"f7",x"c0"),
    82 => (x"f0",x"c0",x"87",x"c3"),
    83 => (x"02",x"66",x"c8",x"82"),
    84 => (x"72",x"87",x"cc",x"c0"),
    85 => (x"00",x"45",x"27",x"1e"),
    86 => (x"c4",x"0f",x"00",x"00"),
    87 => (x"cc",x"83",x"c1",x"86"),
    88 => (x"80",x"c1",x"48",x"66"),
    89 => (x"cc",x"58",x"a6",x"d0"),
    90 => (x"b7",x"c8",x"48",x"66"),
    91 => (x"f2",x"fe",x"04",x"a8"),
    92 => (x"87",x"ea",x"c1",x"87"),
    93 => (x"27",x"1e",x"f0",x"c0"),
    94 => (x"00",x"00",x"00",x"45"),
    95 => (x"c1",x"86",x"c4",x"0f"),
    96 => (x"87",x"da",x"c1",x"83"),
    97 => (x"49",x"74",x"84",x"c4"),
    98 => (x"1e",x"69",x"89",x"c4"),
    99 => (x"00",x"00",x"68",x"27"),
   100 => (x"86",x"c4",x"0f",x"00"),
   101 => (x"83",x"71",x"49",x"70"),
   102 => (x"c4",x"87",x"c3",x"c1"),
   103 => (x"78",x"c1",x"48",x"a6"),
   104 => (x"c4",x"87",x"fb",x"c0"),
   105 => (x"c4",x"49",x"74",x"84"),
   106 => (x"27",x"1e",x"69",x"89"),
   107 => (x"00",x"00",x"00",x"45"),
   108 => (x"c1",x"86",x"c4",x"0f"),
   109 => (x"87",x"e6",x"c0",x"83"),
   110 => (x"45",x"27",x"1e",x"72"),
   111 => (x"0f",x"00",x"00",x"00"),
   112 => (x"d9",x"c0",x"86",x"c4"),
   113 => (x"aa",x"e5",x"c0",x"87"),
   114 => (x"87",x"c8",x"c0",x"05"),
   115 => (x"c1",x"48",x"a6",x"c4"),
   116 => (x"87",x"ca",x"c0",x"78"),
   117 => (x"45",x"27",x"1e",x"72"),
   118 => (x"0f",x"00",x"00",x"00"),
   119 => (x"e0",x"c0",x"86",x"c4"),
   120 => (x"c1",x"48",x"49",x"66"),
   121 => (x"a6",x"e4",x"c0",x"80"),
   122 => (x"fe",x"4a",x"11",x"58"),
   123 => (x"72",x"ba",x"82",x"c0"),
   124 => (x"d1",x"fb",x"05",x"9a"),
   125 => (x"f0",x"48",x"73",x"87"),
   126 => (x"26",x"4d",x"26",x"8e"),
   127 => (x"26",x"4b",x"26",x"4c"),
   128 => (x"00",x"00",x"00",x"4f"),
   129 => (x"1e",x"75",x"1e",x"00"),
   130 => (x"c3",x"4d",x"d4",x"ff"),
   131 => (x"6d",x"7d",x"49",x"ff"),
   132 => (x"71",x"38",x"c8",x"48"),
   133 => (x"c8",x"b0",x"6d",x"7d"),
   134 => (x"6d",x"7d",x"71",x"38"),
   135 => (x"71",x"38",x"c8",x"b0"),
   136 => (x"c8",x"b0",x"6d",x"7d"),
   137 => (x"26",x"4d",x"26",x"38"),
   138 => (x"1e",x"75",x"1e",x"4f"),
   139 => (x"c3",x"4d",x"d4",x"ff"),
   140 => (x"6d",x"7d",x"49",x"ff"),
   141 => (x"71",x"30",x"c8",x"48"),
   142 => (x"c8",x"b0",x"6d",x"7d"),
   143 => (x"6d",x"7d",x"71",x"30"),
   144 => (x"71",x"30",x"c8",x"b0"),
   145 => (x"26",x"b0",x"6d",x"7d"),
   146 => (x"1e",x"4f",x"26",x"4d"),
   147 => (x"d4",x"ff",x"1e",x"75"),
   148 => (x"49",x"66",x"cc",x"4d"),
   149 => (x"7d",x"48",x"66",x"c8"),
   150 => (x"02",x"67",x"e6",x"fe"),
   151 => (x"d8",x"07",x"31",x"c9"),
   152 => (x"09",x"7d",x"09",x"39"),
   153 => (x"09",x"7d",x"09",x"39"),
   154 => (x"09",x"7d",x"09",x"39"),
   155 => (x"d0",x"7d",x"09",x"39"),
   156 => (x"c9",x"7d",x"70",x"38"),
   157 => (x"c3",x"49",x"c0",x"f1"),
   158 => (x"08",x"6d",x"48",x"ff"),
   159 => (x"87",x"c7",x"05",x"a8"),
   160 => (x"89",x"c1",x"7d",x"08"),
   161 => (x"26",x"87",x"f3",x"05"),
   162 => (x"1e",x"4f",x"26",x"4d"),
   163 => (x"c3",x"49",x"d4",x"ff"),
   164 => (x"79",x"ff",x"48",x"c8"),
   165 => (x"87",x"fa",x"05",x"80"),
   166 => (x"5e",x"0e",x"4f",x"26"),
   167 => (x"5d",x"5c",x"5b",x"5a"),
   168 => (x"f0",x"ff",x"c0",x"0e"),
   169 => (x"c1",x"4d",x"f7",x"c1"),
   170 => (x"c0",x"c0",x"c0",x"c0"),
   171 => (x"8b",x"27",x"4b",x"c0"),
   172 => (x"0f",x"00",x"00",x"02"),
   173 => (x"4c",x"df",x"f8",x"c4"),
   174 => (x"1e",x"75",x"1e",x"c0"),
   175 => (x"00",x"02",x"4b",x"27"),
   176 => (x"86",x"c8",x"0f",x"00"),
   177 => (x"b7",x"c1",x"4a",x"70"),
   178 => (x"ef",x"c0",x"05",x"aa"),
   179 => (x"49",x"d4",x"ff",x"87"),
   180 => (x"73",x"79",x"ff",x"c3"),
   181 => (x"f0",x"e1",x"c0",x"1e"),
   182 => (x"27",x"1e",x"e9",x"c1"),
   183 => (x"00",x"00",x"02",x"4b"),
   184 => (x"70",x"86",x"c8",x"0f"),
   185 => (x"05",x"9a",x"72",x"4a"),
   186 => (x"ff",x"87",x"cb",x"c0"),
   187 => (x"ff",x"c3",x"49",x"d4"),
   188 => (x"c0",x"48",x"c1",x"79"),
   189 => (x"8b",x"27",x"87",x"d0"),
   190 => (x"0f",x"00",x"00",x"02"),
   191 => (x"9c",x"74",x"8c",x"c1"),
   192 => (x"87",x"f4",x"fe",x"05"),
   193 => (x"4d",x"26",x"48",x"c0"),
   194 => (x"4b",x"26",x"4c",x"26"),
   195 => (x"4f",x"26",x"4a",x"26"),
   196 => (x"5b",x"5a",x"5e",x"0e"),
   197 => (x"ff",x"c0",x"0e",x"5c"),
   198 => (x"4c",x"c1",x"c1",x"f0"),
   199 => (x"c3",x"49",x"d4",x"ff"),
   200 => (x"4c",x"27",x"79",x"ff"),
   201 => (x"1e",x"00",x"00",x"16"),
   202 => (x"00",x"00",x"68",x"27"),
   203 => (x"86",x"c4",x"0f",x"00"),
   204 => (x"1e",x"c0",x"4b",x"d3"),
   205 => (x"4b",x"27",x"1e",x"74"),
   206 => (x"0f",x"00",x"00",x"02"),
   207 => (x"4a",x"70",x"86",x"c8"),
   208 => (x"c0",x"05",x"9a",x"72"),
   209 => (x"d4",x"ff",x"87",x"cb"),
   210 => (x"79",x"ff",x"c3",x"49"),
   211 => (x"d0",x"c0",x"48",x"c1"),
   212 => (x"02",x"8b",x"27",x"87"),
   213 => (x"c1",x"0f",x"00",x"00"),
   214 => (x"05",x"9b",x"73",x"8b"),
   215 => (x"c0",x"87",x"d3",x"ff"),
   216 => (x"26",x"4c",x"26",x"48"),
   217 => (x"26",x"4a",x"26",x"4b"),
   218 => (x"5a",x"5e",x"0e",x"4f"),
   219 => (x"0e",x"5d",x"5c",x"5b"),
   220 => (x"4d",x"ff",x"c3",x"1e"),
   221 => (x"27",x"4c",x"d4",x"ff"),
   222 => (x"00",x"00",x"02",x"8b"),
   223 => (x"1e",x"ea",x"c6",x"0f"),
   224 => (x"c1",x"f0",x"e1",x"c0"),
   225 => (x"4b",x"27",x"1e",x"c8"),
   226 => (x"0f",x"00",x"00",x"02"),
   227 => (x"4a",x"70",x"86",x"c8"),
   228 => (x"c8",x"27",x"1e",x"72"),
   229 => (x"1e",x"00",x"00",x"04"),
   230 => (x"00",x"00",x"9c",x"27"),
   231 => (x"86",x"c8",x"0f",x"00"),
   232 => (x"02",x"aa",x"b7",x"c1"),
   233 => (x"27",x"87",x"cb",x"c0"),
   234 => (x"00",x"00",x"03",x"10"),
   235 => (x"c3",x"48",x"c0",x"0f"),
   236 => (x"29",x"27",x"87",x"c9"),
   237 => (x"0f",x"00",x"00",x"02"),
   238 => (x"ff",x"cf",x"4a",x"70"),
   239 => (x"ea",x"c6",x"9a",x"ff"),
   240 => (x"c0",x"02",x"aa",x"b7"),
   241 => (x"10",x"27",x"87",x"cb"),
   242 => (x"0f",x"00",x"00",x"03"),
   243 => (x"ea",x"c2",x"48",x"c0"),
   244 => (x"76",x"7c",x"75",x"87"),
   245 => (x"79",x"f1",x"c0",x"49"),
   246 => (x"00",x"02",x"9a",x"27"),
   247 => (x"4a",x"70",x"0f",x"00"),
   248 => (x"c1",x"02",x"9a",x"72"),
   249 => (x"1e",x"c0",x"87",x"eb"),
   250 => (x"c1",x"f0",x"ff",x"c0"),
   251 => (x"4b",x"27",x"1e",x"fa"),
   252 => (x"0f",x"00",x"00",x"02"),
   253 => (x"4b",x"70",x"86",x"c8"),
   254 => (x"c1",x"05",x"9b",x"73"),
   255 => (x"1e",x"73",x"87",x"c3"),
   256 => (x"00",x"04",x"86",x"27"),
   257 => (x"9c",x"27",x"1e",x"00"),
   258 => (x"0f",x"00",x"00",x"00"),
   259 => (x"7c",x"75",x"86",x"c8"),
   260 => (x"9b",x"75",x"4b",x"6c"),
   261 => (x"92",x"27",x"1e",x"73"),
   262 => (x"1e",x"00",x"00",x"04"),
   263 => (x"00",x"00",x"9c",x"27"),
   264 => (x"86",x"c8",x"0f",x"00"),
   265 => (x"7c",x"75",x"7c",x"75"),
   266 => (x"7c",x"75",x"7c",x"75"),
   267 => (x"c0",x"c1",x"4a",x"73"),
   268 => (x"02",x"9a",x"72",x"9a"),
   269 => (x"c1",x"87",x"c5",x"c0"),
   270 => (x"87",x"ff",x"c0",x"48"),
   271 => (x"fa",x"c0",x"48",x"c0"),
   272 => (x"27",x"1e",x"73",x"87"),
   273 => (x"00",x"00",x"04",x"a0"),
   274 => (x"00",x"9c",x"27",x"1e"),
   275 => (x"c8",x"0f",x"00",x"00"),
   276 => (x"c2",x"49",x"6e",x"86"),
   277 => (x"c0",x"05",x"a9",x"b7"),
   278 => (x"ac",x"27",x"87",x"d3"),
   279 => (x"1e",x"00",x"00",x"04"),
   280 => (x"00",x"00",x"9c",x"27"),
   281 => (x"86",x"c4",x"0f",x"00"),
   282 => (x"ce",x"c0",x"48",x"c0"),
   283 => (x"c1",x"48",x"6e",x"87"),
   284 => (x"58",x"a6",x"c4",x"88"),
   285 => (x"df",x"fd",x"05",x"6e"),
   286 => (x"26",x"48",x"c0",x"87"),
   287 => (x"4c",x"26",x"4d",x"26"),
   288 => (x"4a",x"26",x"4b",x"26"),
   289 => (x"4d",x"43",x"4f",x"26"),
   290 => (x"20",x"38",x"35",x"44"),
   291 => (x"20",x"0a",x"64",x"25"),
   292 => (x"4d",x"43",x"00",x"20"),
   293 => (x"5f",x"38",x"35",x"44"),
   294 => (x"64",x"25",x"20",x"32"),
   295 => (x"00",x"20",x"20",x"0a"),
   296 => (x"35",x"44",x"4d",x"43"),
   297 => (x"64",x"25",x"20",x"38"),
   298 => (x"00",x"20",x"20",x"0a"),
   299 => (x"43",x"48",x"44",x"53"),
   300 => (x"69",x"6e",x"49",x"20"),
   301 => (x"6c",x"61",x"69",x"74"),
   302 => (x"74",x"61",x"7a",x"69"),
   303 => (x"20",x"6e",x"6f",x"69"),
   304 => (x"6f",x"72",x"72",x"65"),
   305 => (x"00",x"0a",x"21",x"72"),
   306 => (x"5f",x"64",x"6d",x"63"),
   307 => (x"38",x"44",x"4d",x"43"),
   308 => (x"73",x"65",x"72",x"20"),
   309 => (x"73",x"6e",x"6f",x"70"),
   310 => (x"25",x"20",x"3a",x"65"),
   311 => (x"0e",x"00",x"0a",x"64"),
   312 => (x"5c",x"5b",x"5a",x"5e"),
   313 => (x"ff",x"1e",x"0e",x"5d"),
   314 => (x"c0",x"c8",x"4c",x"d0"),
   315 => (x"01",x"27",x"4b",x"c0"),
   316 => (x"49",x"00",x"00",x"02"),
   317 => (x"fc",x"27",x"79",x"c1"),
   318 => (x"1e",x"00",x"00",x"05"),
   319 => (x"00",x"00",x"68",x"27"),
   320 => (x"86",x"c4",x"0f",x"00"),
   321 => (x"48",x"6c",x"4d",x"c7"),
   322 => (x"a6",x"c4",x"98",x"73"),
   323 => (x"c0",x"02",x"6e",x"58"),
   324 => (x"48",x"6c",x"87",x"cc"),
   325 => (x"a6",x"c4",x"98",x"73"),
   326 => (x"ff",x"05",x"6e",x"58"),
   327 => (x"7c",x"c0",x"87",x"f4"),
   328 => (x"00",x"02",x"8b",x"27"),
   329 => (x"48",x"6c",x"0f",x"00"),
   330 => (x"a6",x"c4",x"98",x"73"),
   331 => (x"c0",x"02",x"6e",x"58"),
   332 => (x"48",x"6c",x"87",x"cc"),
   333 => (x"a6",x"c4",x"98",x"73"),
   334 => (x"ff",x"05",x"6e",x"58"),
   335 => (x"7c",x"c1",x"87",x"f4"),
   336 => (x"e5",x"c0",x"1e",x"c0"),
   337 => (x"1e",x"c0",x"c1",x"d0"),
   338 => (x"00",x"02",x"4b",x"27"),
   339 => (x"86",x"c8",x"0f",x"00"),
   340 => (x"b7",x"c1",x"4a",x"70"),
   341 => (x"c2",x"c0",x"05",x"aa"),
   342 => (x"c2",x"4d",x"c1",x"87"),
   343 => (x"c0",x"05",x"ad",x"b7"),
   344 => (x"f7",x"27",x"87",x"d3"),
   345 => (x"1e",x"00",x"00",x"05"),
   346 => (x"00",x"00",x"68",x"27"),
   347 => (x"86",x"c4",x"0f",x"00"),
   348 => (x"f7",x"c1",x"48",x"c0"),
   349 => (x"75",x"8d",x"c1",x"87"),
   350 => (x"c9",x"fe",x"05",x"9d"),
   351 => (x"03",x"69",x"27",x"87"),
   352 => (x"27",x"0f",x"00",x"00"),
   353 => (x"00",x"00",x"02",x"05"),
   354 => (x"02",x"01",x"27",x"58"),
   355 => (x"05",x"bf",x"00",x"00"),
   356 => (x"c1",x"87",x"d0",x"c0"),
   357 => (x"f0",x"ff",x"c0",x"1e"),
   358 => (x"27",x"1e",x"d0",x"c1"),
   359 => (x"00",x"00",x"02",x"4b"),
   360 => (x"ff",x"86",x"c8",x"0f"),
   361 => (x"ff",x"c3",x"49",x"d4"),
   362 => (x"08",x"92",x"27",x"79"),
   363 => (x"27",x"0f",x"00",x"00"),
   364 => (x"00",x"00",x"17",x"e8"),
   365 => (x"17",x"e4",x"27",x"58"),
   366 => (x"1e",x"bf",x"00",x"00"),
   367 => (x"00",x"06",x"00",x"27"),
   368 => (x"9c",x"27",x"1e",x"00"),
   369 => (x"0f",x"00",x"00",x"00"),
   370 => (x"48",x"6c",x"86",x"c8"),
   371 => (x"a6",x"c4",x"98",x"73"),
   372 => (x"c0",x"02",x"6e",x"58"),
   373 => (x"48",x"6c",x"87",x"cc"),
   374 => (x"a6",x"c4",x"98",x"73"),
   375 => (x"ff",x"05",x"6e",x"58"),
   376 => (x"7c",x"c0",x"87",x"f4"),
   377 => (x"c3",x"49",x"d4",x"ff"),
   378 => (x"48",x"c1",x"79",x"ff"),
   379 => (x"26",x"4d",x"26",x"26"),
   380 => (x"26",x"4b",x"26",x"4c"),
   381 => (x"49",x"4f",x"26",x"4a"),
   382 => (x"00",x"52",x"52",x"45"),
   383 => (x"00",x"49",x"50",x"53"),
   384 => (x"63",x"20",x"44",x"53"),
   385 => (x"20",x"64",x"72",x"61"),
   386 => (x"65",x"7a",x"69",x"73"),
   387 => (x"20",x"73",x"69",x"20"),
   388 => (x"00",x"0a",x"64",x"25"),
   389 => (x"5b",x"5a",x"5e",x"0e"),
   390 => (x"1e",x"0e",x"5d",x"5c"),
   391 => (x"ff",x"4d",x"ff",x"c3"),
   392 => (x"7c",x"75",x"4c",x"d4"),
   393 => (x"48",x"bf",x"d0",x"ff"),
   394 => (x"98",x"c0",x"c0",x"c8"),
   395 => (x"6e",x"58",x"a6",x"c4"),
   396 => (x"87",x"d2",x"c0",x"02"),
   397 => (x"4a",x"c0",x"c0",x"c8"),
   398 => (x"48",x"bf",x"d0",x"ff"),
   399 => (x"a6",x"c4",x"98",x"72"),
   400 => (x"ff",x"05",x"6e",x"58"),
   401 => (x"d0",x"ff",x"87",x"f2"),
   402 => (x"79",x"c1",x"c4",x"49"),
   403 => (x"66",x"d8",x"7c",x"75"),
   404 => (x"f0",x"ff",x"c0",x"1e"),
   405 => (x"27",x"1e",x"d8",x"c1"),
   406 => (x"00",x"00",x"02",x"4b"),
   407 => (x"70",x"86",x"c8",x"0f"),
   408 => (x"02",x"9a",x"72",x"4a"),
   409 => (x"27",x"87",x"d3",x"c0"),
   410 => (x"00",x"00",x"07",x"1c"),
   411 => (x"00",x"68",x"27",x"1e"),
   412 => (x"c4",x"0f",x"00",x"00"),
   413 => (x"c2",x"48",x"c1",x"86"),
   414 => (x"7c",x"75",x"87",x"d7"),
   415 => (x"76",x"7c",x"fe",x"c3"),
   416 => (x"dc",x"79",x"c0",x"49"),
   417 => (x"72",x"4a",x"bf",x"66"),
   418 => (x"2b",x"b7",x"d8",x"4b"),
   419 => (x"98",x"75",x"48",x"73"),
   420 => (x"4b",x"72",x"7c",x"70"),
   421 => (x"73",x"2b",x"b7",x"d0"),
   422 => (x"70",x"98",x"75",x"48"),
   423 => (x"c8",x"4b",x"72",x"7c"),
   424 => (x"48",x"73",x"2b",x"b7"),
   425 => (x"7c",x"70",x"98",x"75"),
   426 => (x"98",x"75",x"48",x"72"),
   427 => (x"66",x"dc",x"7c",x"70"),
   428 => (x"c0",x"80",x"c4",x"48"),
   429 => (x"6e",x"58",x"a6",x"e0"),
   430 => (x"c4",x"80",x"c1",x"48"),
   431 => (x"49",x"6e",x"58",x"a6"),
   432 => (x"a9",x"b7",x"c0",x"c2"),
   433 => (x"87",x"fb",x"fe",x"04"),
   434 => (x"7c",x"75",x"7c",x"75"),
   435 => (x"da",x"d8",x"7c",x"75"),
   436 => (x"7c",x"75",x"4b",x"e0"),
   437 => (x"9a",x"75",x"4a",x"6c"),
   438 => (x"c0",x"05",x"9a",x"72"),
   439 => (x"8b",x"c1",x"87",x"c8"),
   440 => (x"ff",x"05",x"9b",x"73"),
   441 => (x"7c",x"75",x"87",x"ec"),
   442 => (x"48",x"bf",x"d0",x"ff"),
   443 => (x"98",x"c0",x"c0",x"c8"),
   444 => (x"6e",x"58",x"a6",x"c4"),
   445 => (x"87",x"d2",x"c0",x"02"),
   446 => (x"4a",x"c0",x"c0",x"c8"),
   447 => (x"48",x"bf",x"d0",x"ff"),
   448 => (x"a6",x"c4",x"98",x"72"),
   449 => (x"ff",x"05",x"6e",x"58"),
   450 => (x"d0",x"ff",x"87",x"f2"),
   451 => (x"c0",x"79",x"c0",x"49"),
   452 => (x"4d",x"26",x"26",x"48"),
   453 => (x"4b",x"26",x"4c",x"26"),
   454 => (x"4f",x"26",x"4a",x"26"),
   455 => (x"74",x"69",x"72",x"57"),
   456 => (x"61",x"66",x"20",x"65"),
   457 => (x"64",x"65",x"6c",x"69"),
   458 => (x"5e",x"0e",x"00",x"0a"),
   459 => (x"5d",x"5c",x"5b",x"5a"),
   460 => (x"66",x"d8",x"1e",x"0e"),
   461 => (x"4b",x"66",x"dc",x"4c"),
   462 => (x"79",x"c0",x"49",x"76"),
   463 => (x"df",x"cd",x"ee",x"c5"),
   464 => (x"49",x"d4",x"ff",x"4d"),
   465 => (x"ff",x"79",x"ff",x"c3"),
   466 => (x"c3",x"4a",x"bf",x"d4"),
   467 => (x"fe",x"c3",x"9a",x"ff"),
   468 => (x"c1",x"05",x"aa",x"b7"),
   469 => (x"e0",x"27",x"87",x"e5"),
   470 => (x"49",x"00",x"00",x"17"),
   471 => (x"b7",x"c4",x"79",x"c0"),
   472 => (x"e4",x"c0",x"04",x"ab"),
   473 => (x"02",x"05",x"27",x"87"),
   474 => (x"70",x"0f",x"00",x"00"),
   475 => (x"c4",x"7c",x"72",x"4a"),
   476 => (x"17",x"e0",x"27",x"84"),
   477 => (x"48",x"bf",x"00",x"00"),
   478 => (x"e4",x"27",x"80",x"72"),
   479 => (x"58",x"00",x"00",x"17"),
   480 => (x"b7",x"c4",x"8b",x"c4"),
   481 => (x"dc",x"ff",x"03",x"ab"),
   482 => (x"ab",x"b7",x"c0",x"87"),
   483 => (x"87",x"e5",x"c0",x"06"),
   484 => (x"c3",x"4d",x"d4",x"ff"),
   485 => (x"4a",x"6d",x"7d",x"ff"),
   486 => (x"c1",x"7c",x"97",x"72"),
   487 => (x"17",x"e0",x"27",x"84"),
   488 => (x"48",x"bf",x"00",x"00"),
   489 => (x"e4",x"27",x"80",x"72"),
   490 => (x"58",x"00",x"00",x"17"),
   491 => (x"b7",x"c0",x"8b",x"c1"),
   492 => (x"de",x"ff",x"01",x"ab"),
   493 => (x"76",x"4d",x"c1",x"87"),
   494 => (x"c1",x"79",x"c1",x"49"),
   495 => (x"05",x"9d",x"75",x"8d"),
   496 => (x"ff",x"87",x"fe",x"fd"),
   497 => (x"ff",x"c3",x"49",x"d4"),
   498 => (x"26",x"48",x"6e",x"79"),
   499 => (x"4c",x"26",x"4d",x"26"),
   500 => (x"4a",x"26",x"4b",x"26"),
   501 => (x"5e",x"0e",x"4f",x"26"),
   502 => (x"5d",x"5c",x"5b",x"5a"),
   503 => (x"d0",x"ff",x"1e",x"0e"),
   504 => (x"c0",x"c0",x"c8",x"4b"),
   505 => (x"ff",x"4c",x"c0",x"4a"),
   506 => (x"ff",x"c3",x"49",x"d4"),
   507 => (x"72",x"48",x"6b",x"79"),
   508 => (x"58",x"a6",x"c4",x"98"),
   509 => (x"cc",x"c0",x"02",x"6e"),
   510 => (x"72",x"48",x"6b",x"87"),
   511 => (x"58",x"a6",x"c4",x"98"),
   512 => (x"f4",x"ff",x"05",x"6e"),
   513 => (x"7b",x"c1",x"c4",x"87"),
   514 => (x"c3",x"49",x"d4",x"ff"),
   515 => (x"66",x"d8",x"79",x"ff"),
   516 => (x"f0",x"ff",x"c0",x"1e"),
   517 => (x"27",x"1e",x"d1",x"c1"),
   518 => (x"00",x"00",x"02",x"4b"),
   519 => (x"70",x"86",x"c8",x"0f"),
   520 => (x"02",x"9d",x"75",x"4d"),
   521 => (x"75",x"87",x"d6",x"c0"),
   522 => (x"1e",x"66",x"dc",x"1e"),
   523 => (x"00",x"08",x"72",x"27"),
   524 => (x"9c",x"27",x"1e",x"00"),
   525 => (x"0f",x"00",x"00",x"00"),
   526 => (x"e8",x"c0",x"86",x"cc"),
   527 => (x"1e",x"c0",x"c8",x"87"),
   528 => (x"1e",x"66",x"e0",x"c0"),
   529 => (x"c8",x"87",x"e3",x"fb"),
   530 => (x"6b",x"4c",x"70",x"86"),
   531 => (x"c4",x"98",x"72",x"48"),
   532 => (x"02",x"6e",x"58",x"a6"),
   533 => (x"6b",x"87",x"cc",x"c0"),
   534 => (x"c4",x"98",x"72",x"48"),
   535 => (x"05",x"6e",x"58",x"a6"),
   536 => (x"c0",x"87",x"f4",x"ff"),
   537 => (x"26",x"48",x"74",x"7b"),
   538 => (x"4c",x"26",x"4d",x"26"),
   539 => (x"4a",x"26",x"4b",x"26"),
   540 => (x"65",x"52",x"4f",x"26"),
   541 => (x"63",x"20",x"64",x"61"),
   542 => (x"61",x"6d",x"6d",x"6f"),
   543 => (x"66",x"20",x"64",x"6e"),
   544 => (x"65",x"6c",x"69",x"61"),
   545 => (x"74",x"61",x"20",x"64"),
   546 => (x"20",x"64",x"25",x"20"),
   547 => (x"29",x"64",x"25",x"28"),
   548 => (x"5e",x"0e",x"00",x"0a"),
   549 => (x"5d",x"5c",x"5b",x"5a"),
   550 => (x"1e",x"c0",x"1e",x"0e"),
   551 => (x"c1",x"f0",x"ff",x"c0"),
   552 => (x"4b",x"27",x"1e",x"c9"),
   553 => (x"0f",x"00",x"00",x"02"),
   554 => (x"1e",x"d2",x"86",x"c8"),
   555 => (x"00",x"17",x"f0",x"27"),
   556 => (x"f5",x"f9",x"1e",x"00"),
   557 => (x"c0",x"86",x"c8",x"87"),
   558 => (x"d2",x"85",x"c1",x"4d"),
   559 => (x"ff",x"04",x"ad",x"b7"),
   560 => (x"f0",x"27",x"87",x"f7"),
   561 => (x"97",x"00",x"00",x"17"),
   562 => (x"c0",x"c3",x"4a",x"bf"),
   563 => (x"b7",x"c0",x"c1",x"9a"),
   564 => (x"f2",x"c0",x"05",x"aa"),
   565 => (x"17",x"f7",x"27",x"87"),
   566 => (x"bf",x"97",x"00",x"00"),
   567 => (x"27",x"32",x"d0",x"4a"),
   568 => (x"00",x"00",x"17",x"f8"),
   569 => (x"c8",x"4b",x"bf",x"97"),
   570 => (x"73",x"4a",x"72",x"33"),
   571 => (x"17",x"f9",x"27",x"b2"),
   572 => (x"bf",x"97",x"00",x"00"),
   573 => (x"73",x"4a",x"72",x"4b"),
   574 => (x"ff",x"ff",x"cf",x"b2"),
   575 => (x"4d",x"72",x"9a",x"ff"),
   576 => (x"35",x"ca",x"85",x"c1"),
   577 => (x"27",x"87",x"cb",x"c3"),
   578 => (x"00",x"00",x"17",x"f9"),
   579 => (x"c1",x"4a",x"bf",x"97"),
   580 => (x"27",x"9a",x"c6",x"32"),
   581 => (x"00",x"00",x"17",x"fa"),
   582 => (x"c7",x"4b",x"bf",x"97"),
   583 => (x"4a",x"72",x"2b",x"b7"),
   584 => (x"f5",x"27",x"b2",x"73"),
   585 => (x"97",x"00",x"00",x"17"),
   586 => (x"48",x"73",x"4b",x"bf"),
   587 => (x"a6",x"c4",x"98",x"cf"),
   588 => (x"17",x"f6",x"27",x"58"),
   589 => (x"bf",x"97",x"00",x"00"),
   590 => (x"ca",x"9b",x"c3",x"4b"),
   591 => (x"17",x"f7",x"27",x"33"),
   592 => (x"bf",x"97",x"00",x"00"),
   593 => (x"73",x"34",x"c2",x"4c"),
   594 => (x"27",x"b3",x"74",x"4b"),
   595 => (x"00",x"00",x"17",x"f8"),
   596 => (x"c3",x"4c",x"bf",x"97"),
   597 => (x"b7",x"c6",x"9c",x"c0"),
   598 => (x"74",x"4b",x"73",x"2c"),
   599 => (x"c4",x"1e",x"73",x"b3"),
   600 => (x"1e",x"72",x"1e",x"66"),
   601 => (x"00",x"09",x"df",x"27"),
   602 => (x"9c",x"27",x"1e",x"00"),
   603 => (x"0f",x"00",x"00",x"00"),
   604 => (x"82",x"c2",x"86",x"d0"),
   605 => (x"30",x"72",x"48",x"c1"),
   606 => (x"1e",x"72",x"4a",x"70"),
   607 => (x"00",x"0a",x"0c",x"27"),
   608 => (x"9c",x"27",x"1e",x"00"),
   609 => (x"0f",x"00",x"00",x"00"),
   610 => (x"48",x"c1",x"86",x"c8"),
   611 => (x"a6",x"c4",x"30",x"6e"),
   612 => (x"73",x"83",x"c1",x"58"),
   613 => (x"6e",x"95",x"72",x"4d"),
   614 => (x"27",x"1e",x"75",x"1e"),
   615 => (x"00",x"00",x"0a",x"15"),
   616 => (x"00",x"9c",x"27",x"1e"),
   617 => (x"cc",x"0f",x"00",x"00"),
   618 => (x"c8",x"49",x"6e",x"86"),
   619 => (x"06",x"a9",x"b7",x"c0"),
   620 => (x"6e",x"87",x"cf",x"c0"),
   621 => (x"c1",x"35",x"c1",x"4a"),
   622 => (x"c0",x"c8",x"2a",x"b7"),
   623 => (x"ff",x"01",x"aa",x"b7"),
   624 => (x"1e",x"75",x"87",x"f3"),
   625 => (x"00",x"0a",x"2b",x"27"),
   626 => (x"9c",x"27",x"1e",x"00"),
   627 => (x"0f",x"00",x"00",x"00"),
   628 => (x"48",x"75",x"86",x"c8"),
   629 => (x"26",x"4d",x"26",x"26"),
   630 => (x"26",x"4b",x"26",x"4c"),
   631 => (x"63",x"4f",x"26",x"4a"),
   632 => (x"7a",x"69",x"73",x"5f"),
   633 => (x"75",x"6d",x"5f",x"65"),
   634 => (x"20",x"3a",x"74",x"6c"),
   635 => (x"20",x"2c",x"64",x"25"),
   636 => (x"64",x"61",x"65",x"72"),
   637 => (x"5f",x"6c",x"62",x"5f"),
   638 => (x"3a",x"6e",x"65",x"6c"),
   639 => (x"2c",x"64",x"25",x"20"),
   640 => (x"69",x"73",x"63",x"20"),
   641 => (x"20",x"3a",x"65",x"7a"),
   642 => (x"00",x"0a",x"64",x"25"),
   643 => (x"74",x"6c",x"75",x"4d"),
   644 => (x"0a",x"64",x"25",x"20"),
   645 => (x"20",x"64",x"25",x"00"),
   646 => (x"63",x"6f",x"6c",x"62"),
   647 => (x"6f",x"20",x"73",x"6b"),
   648 => (x"69",x"73",x"20",x"66"),
   649 => (x"25",x"20",x"65",x"7a"),
   650 => (x"25",x"00",x"0a",x"64"),
   651 => (x"6c",x"62",x"20",x"64"),
   652 => (x"73",x"6b",x"63",x"6f"),
   653 => (x"20",x"66",x"6f",x"20"),
   654 => (x"20",x"32",x"31",x"35"),
   655 => (x"65",x"74",x"79",x"62"),
   656 => (x"0e",x"00",x"0a",x"73"),
   657 => (x"c0",x"0e",x"5b",x"5e"),
   658 => (x"48",x"66",x"d0",x"4b"),
   659 => (x"06",x"a8",x"b7",x"c0"),
   660 => (x"c8",x"87",x"f8",x"c0"),
   661 => (x"4a",x"bf",x"97",x"66"),
   662 => (x"ba",x"82",x"c0",x"fe"),
   663 => (x"c1",x"48",x"66",x"c8"),
   664 => (x"58",x"a6",x"cc",x"80"),
   665 => (x"bf",x"97",x"66",x"cc"),
   666 => (x"81",x"c0",x"fe",x"49"),
   667 => (x"48",x"66",x"cc",x"b9"),
   668 => (x"a6",x"d0",x"80",x"c1"),
   669 => (x"aa",x"b7",x"71",x"58"),
   670 => (x"87",x"c5",x"c0",x"02"),
   671 => (x"cc",x"c0",x"48",x"c1"),
   672 => (x"d0",x"83",x"c1",x"87"),
   673 => (x"04",x"ab",x"b7",x"66"),
   674 => (x"c0",x"87",x"c8",x"ff"),
   675 => (x"c4",x"c0",x"c0",x"48"),
   676 => (x"26",x"4d",x"26",x"87"),
   677 => (x"26",x"4b",x"26",x"4c"),
   678 => (x"5b",x"5e",x"0e",x"4f"),
   679 => (x"27",x"0e",x"5d",x"5c"),
   680 => (x"00",x"00",x"18",x"10"),
   681 => (x"27",x"78",x"c0",x"48"),
   682 => (x"00",x"00",x"17",x"24"),
   683 => (x"00",x"68",x"27",x"1e"),
   684 => (x"c4",x"0f",x"00",x"00"),
   685 => (x"18",x"50",x"27",x"86"),
   686 => (x"c0",x"1e",x"00",x"00"),
   687 => (x"07",x"d6",x"27",x"1e"),
   688 => (x"c8",x"0f",x"00",x"00"),
   689 => (x"05",x"98",x"70",x"86"),
   690 => (x"27",x"87",x"d3",x"c0"),
   691 => (x"00",x"00",x"16",x"50"),
   692 => (x"00",x"68",x"27",x"1e"),
   693 => (x"c4",x"0f",x"00",x"00"),
   694 => (x"ce",x"48",x"c0",x"86"),
   695 => (x"31",x"27",x"87",x"d9"),
   696 => (x"1e",x"00",x"00",x"17"),
   697 => (x"00",x"00",x"68",x"27"),
   698 => (x"86",x"c4",x"0f",x"00"),
   699 => (x"3c",x"27",x"4b",x"c0"),
   700 => (x"48",x"00",x"00",x"18"),
   701 => (x"1e",x"c8",x"78",x"c1"),
   702 => (x"00",x"17",x"48",x"27"),
   703 => (x"86",x"27",x"1e",x"00"),
   704 => (x"1e",x"00",x"00",x"18"),
   705 => (x"00",x"0a",x"43",x"27"),
   706 => (x"86",x"cc",x"0f",x"00"),
   707 => (x"c0",x"05",x"98",x"70"),
   708 => (x"3c",x"27",x"87",x"c8"),
   709 => (x"48",x"00",x"00",x"18"),
   710 => (x"1e",x"c8",x"78",x"c0"),
   711 => (x"00",x"17",x"51",x"27"),
   712 => (x"a2",x"27",x"1e",x"00"),
   713 => (x"1e",x"00",x"00",x"18"),
   714 => (x"00",x"0a",x"43",x"27"),
   715 => (x"86",x"cc",x"0f",x"00"),
   716 => (x"c0",x"05",x"98",x"70"),
   717 => (x"3c",x"27",x"87",x"c8"),
   718 => (x"48",x"00",x"00",x"18"),
   719 => (x"3c",x"27",x"78",x"c0"),
   720 => (x"bf",x"00",x"00",x"18"),
   721 => (x"17",x"5a",x"27",x"1e"),
   722 => (x"27",x"1e",x"00",x"00"),
   723 => (x"00",x"00",x"00",x"9c"),
   724 => (x"27",x"86",x"c8",x"0f"),
   725 => (x"00",x"00",x"18",x"3c"),
   726 => (x"fc",x"c2",x"02",x"bf"),
   727 => (x"18",x"50",x"27",x"87"),
   728 => (x"27",x"4d",x"00",x"00"),
   729 => (x"00",x"00",x"1a",x"0e"),
   730 => (x"1a",x"4e",x"27",x"4c"),
   731 => (x"bf",x"9f",x"00",x"00"),
   732 => (x"27",x"1e",x"71",x"49"),
   733 => (x"00",x"00",x"1a",x"4e"),
   734 => (x"18",x"50",x"27",x"49"),
   735 => (x"71",x"89",x"00",x"00"),
   736 => (x"c8",x"1e",x"d0",x"1e"),
   737 => (x"82",x"27",x"1e",x"c0"),
   738 => (x"1e",x"00",x"00",x"16"),
   739 => (x"00",x"00",x"9c",x"27"),
   740 => (x"86",x"d4",x"0f",x"00"),
   741 => (x"81",x"c8",x"49",x"74"),
   742 => (x"4e",x"27",x"4b",x"69"),
   743 => (x"9f",x"00",x"00",x"1a"),
   744 => (x"d6",x"c5",x"49",x"bf"),
   745 => (x"c0",x"05",x"a9",x"ea"),
   746 => (x"49",x"74",x"87",x"d3"),
   747 => (x"1e",x"69",x"81",x"c8"),
   748 => (x"00",x"11",x"8f",x"27"),
   749 => (x"86",x"c4",x"0f",x"00"),
   750 => (x"e3",x"c0",x"4b",x"70"),
   751 => (x"c7",x"49",x"75",x"87"),
   752 => (x"69",x"9f",x"81",x"fe"),
   753 => (x"d5",x"e9",x"ca",x"49"),
   754 => (x"d3",x"c0",x"02",x"a9"),
   755 => (x"16",x"64",x"27",x"87"),
   756 => (x"27",x"1e",x"00",x"00"),
   757 => (x"00",x"00",x"00",x"68"),
   758 => (x"c0",x"86",x"c4",x"0f"),
   759 => (x"87",x"d7",x"ca",x"48"),
   760 => (x"bf",x"27",x"1e",x"73"),
   761 => (x"1e",x"00",x"00",x"16"),
   762 => (x"00",x"00",x"9c",x"27"),
   763 => (x"86",x"c8",x"0f",x"00"),
   764 => (x"00",x"18",x"50",x"27"),
   765 => (x"1e",x"73",x"1e",x"00"),
   766 => (x"00",x"07",x"d6",x"27"),
   767 => (x"86",x"c8",x"0f",x"00"),
   768 => (x"c0",x"05",x"98",x"70"),
   769 => (x"48",x"c0",x"87",x"c5"),
   770 => (x"27",x"87",x"ec",x"c9"),
   771 => (x"00",x"00",x"16",x"d7"),
   772 => (x"00",x"68",x"27",x"1e"),
   773 => (x"c4",x"0f",x"00",x"00"),
   774 => (x"17",x"6d",x"27",x"86"),
   775 => (x"27",x"1e",x"00",x"00"),
   776 => (x"00",x"00",x"00",x"9c"),
   777 => (x"c8",x"86",x"c4",x"0f"),
   778 => (x"17",x"85",x"27",x"1e"),
   779 => (x"27",x"1e",x"00",x"00"),
   780 => (x"00",x"00",x"18",x"a2"),
   781 => (x"0a",x"43",x"27",x"1e"),
   782 => (x"cc",x"0f",x"00",x"00"),
   783 => (x"05",x"98",x"70",x"86"),
   784 => (x"27",x"87",x"cb",x"c0"),
   785 => (x"00",x"00",x"18",x"10"),
   786 => (x"c0",x"78",x"c1",x"48"),
   787 => (x"1e",x"c8",x"87",x"ef"),
   788 => (x"00",x"17",x"8e",x"27"),
   789 => (x"86",x"27",x"1e",x"00"),
   790 => (x"1e",x"00",x"00",x"18"),
   791 => (x"00",x"0a",x"43",x"27"),
   792 => (x"86",x"cc",x"0f",x"00"),
   793 => (x"c0",x"02",x"98",x"70"),
   794 => (x"fe",x"27",x"87",x"d3"),
   795 => (x"1e",x"00",x"00",x"16"),
   796 => (x"00",x"00",x"9c",x"27"),
   797 => (x"86",x"c4",x"0f",x"00"),
   798 => (x"fa",x"c7",x"48",x"c0"),
   799 => (x"1a",x"4e",x"27",x"87"),
   800 => (x"bf",x"97",x"00",x"00"),
   801 => (x"a9",x"d5",x"c1",x"49"),
   802 => (x"87",x"cf",x"c0",x"05"),
   803 => (x"00",x"1a",x"4f",x"27"),
   804 => (x"49",x"bf",x"97",x"00"),
   805 => (x"02",x"a9",x"ea",x"c2"),
   806 => (x"c0",x"87",x"c5",x"c0"),
   807 => (x"87",x"d7",x"c7",x"48"),
   808 => (x"00",x"18",x"50",x"27"),
   809 => (x"49",x"bf",x"97",x"00"),
   810 => (x"02",x"a9",x"e9",x"c3"),
   811 => (x"27",x"87",x"d4",x"c0"),
   812 => (x"00",x"00",x"18",x"50"),
   813 => (x"c3",x"49",x"bf",x"97"),
   814 => (x"c0",x"02",x"a9",x"eb"),
   815 => (x"48",x"c0",x"87",x"c5"),
   816 => (x"27",x"87",x"f4",x"c6"),
   817 => (x"00",x"00",x"18",x"5b"),
   818 => (x"71",x"49",x"bf",x"97"),
   819 => (x"ce",x"c0",x"05",x"99"),
   820 => (x"18",x"5c",x"27",x"87"),
   821 => (x"bf",x"97",x"00",x"00"),
   822 => (x"02",x"a9",x"c2",x"49"),
   823 => (x"c0",x"87",x"c5",x"c0"),
   824 => (x"87",x"d3",x"c6",x"48"),
   825 => (x"00",x"18",x"5d",x"27"),
   826 => (x"48",x"bf",x"97",x"00"),
   827 => (x"00",x"18",x"0c",x"27"),
   828 => (x"08",x"27",x"58",x"00"),
   829 => (x"bf",x"00",x"00",x"18"),
   830 => (x"c1",x"4a",x"71",x"49"),
   831 => (x"18",x"10",x"27",x"8a"),
   832 => (x"72",x"5a",x"00",x"00"),
   833 => (x"27",x"1e",x"71",x"1e"),
   834 => (x"00",x"00",x"17",x"97"),
   835 => (x"00",x"9c",x"27",x"1e"),
   836 => (x"cc",x"0f",x"00",x"00"),
   837 => (x"18",x"5e",x"27",x"86"),
   838 => (x"bf",x"97",x"00",x"00"),
   839 => (x"27",x"81",x"73",x"49"),
   840 => (x"00",x"00",x"18",x"5f"),
   841 => (x"c8",x"4a",x"bf",x"97"),
   842 => (x"71",x"48",x"72",x"32"),
   843 => (x"18",x"20",x"27",x"80"),
   844 => (x"27",x"58",x"00",x"00"),
   845 => (x"00",x"00",x"18",x"60"),
   846 => (x"27",x"48",x"bf",x"97"),
   847 => (x"00",x"00",x"18",x"34"),
   848 => (x"18",x"10",x"27",x"58"),
   849 => (x"02",x"bf",x"00",x"00"),
   850 => (x"c8",x"87",x"c3",x"c3"),
   851 => (x"17",x"1b",x"27",x"1e"),
   852 => (x"27",x"1e",x"00",x"00"),
   853 => (x"00",x"00",x"18",x"a2"),
   854 => (x"0a",x"43",x"27",x"1e"),
   855 => (x"cc",x"0f",x"00",x"00"),
   856 => (x"02",x"98",x"70",x"86"),
   857 => (x"c0",x"87",x"c5",x"c0"),
   858 => (x"87",x"cb",x"c4",x"48"),
   859 => (x"00",x"18",x"08",x"27"),
   860 => (x"72",x"4a",x"bf",x"00"),
   861 => (x"27",x"30",x"c4",x"48"),
   862 => (x"00",x"00",x"18",x"38"),
   863 => (x"18",x"30",x"27",x"58"),
   864 => (x"27",x"5a",x"00",x"00"),
   865 => (x"00",x"00",x"18",x"75"),
   866 => (x"c8",x"49",x"bf",x"97"),
   867 => (x"18",x"74",x"27",x"31"),
   868 => (x"bf",x"97",x"00",x"00"),
   869 => (x"27",x"81",x"73",x"4b"),
   870 => (x"00",x"00",x"18",x"76"),
   871 => (x"d0",x"4b",x"bf",x"97"),
   872 => (x"27",x"81",x"73",x"33"),
   873 => (x"00",x"00",x"18",x"77"),
   874 => (x"d8",x"4b",x"bf",x"97"),
   875 => (x"27",x"81",x"73",x"33"),
   876 => (x"00",x"00",x"18",x"3c"),
   877 => (x"18",x"30",x"27",x"59"),
   878 => (x"91",x"bf",x"00",x"00"),
   879 => (x"00",x"18",x"1c",x"27"),
   880 => (x"27",x"81",x"bf",x"00"),
   881 => (x"00",x"00",x"18",x"24"),
   882 => (x"18",x"7d",x"27",x"59"),
   883 => (x"bf",x"97",x"00",x"00"),
   884 => (x"27",x"33",x"c8",x"4b"),
   885 => (x"00",x"00",x"18",x"7c"),
   886 => (x"74",x"4c",x"bf",x"97"),
   887 => (x"18",x"7e",x"27",x"83"),
   888 => (x"bf",x"97",x"00",x"00"),
   889 => (x"74",x"34",x"d0",x"4c"),
   890 => (x"18",x"7f",x"27",x"83"),
   891 => (x"bf",x"97",x"00",x"00"),
   892 => (x"d8",x"9c",x"cf",x"4c"),
   893 => (x"27",x"83",x"74",x"34"),
   894 => (x"00",x"00",x"18",x"28"),
   895 => (x"73",x"8b",x"c2",x"5b"),
   896 => (x"71",x"48",x"72",x"92"),
   897 => (x"18",x"2c",x"27",x"80"),
   898 => (x"c1",x"58",x"00",x"00"),
   899 => (x"62",x"27",x"87",x"e7"),
   900 => (x"97",x"00",x"00",x"18"),
   901 => (x"31",x"c8",x"49",x"bf"),
   902 => (x"00",x"18",x"61",x"27"),
   903 => (x"4a",x"bf",x"97",x"00"),
   904 => (x"38",x"27",x"81",x"72"),
   905 => (x"59",x"00",x"00",x"18"),
   906 => (x"ff",x"c7",x"31",x"c5"),
   907 => (x"27",x"29",x"c9",x"81"),
   908 => (x"00",x"00",x"18",x"30"),
   909 => (x"18",x"67",x"27",x"59"),
   910 => (x"bf",x"97",x"00",x"00"),
   911 => (x"27",x"32",x"c8",x"4a"),
   912 => (x"00",x"00",x"18",x"66"),
   913 => (x"73",x"4b",x"bf",x"97"),
   914 => (x"18",x"3c",x"27",x"82"),
   915 => (x"27",x"5a",x"00",x"00"),
   916 => (x"00",x"00",x"18",x"30"),
   917 => (x"1c",x"27",x"92",x"bf"),
   918 => (x"bf",x"00",x"00",x"18"),
   919 => (x"18",x"2c",x"27",x"82"),
   920 => (x"27",x"5a",x"00",x"00"),
   921 => (x"00",x"00",x"18",x"24"),
   922 => (x"72",x"78",x"c0",x"48"),
   923 => (x"27",x"80",x"71",x"48"),
   924 => (x"00",x"00",x"18",x"24"),
   925 => (x"ff",x"48",x"c1",x"58"),
   926 => (x"0e",x"87",x"d6",x"f0"),
   927 => (x"0e",x"5c",x"5b",x"5e"),
   928 => (x"00",x"18",x"10",x"27"),
   929 => (x"c0",x"02",x"bf",x"00"),
   930 => (x"66",x"cc",x"87",x"cf"),
   931 => (x"2a",x"b7",x"c7",x"4a"),
   932 => (x"c1",x"4b",x"66",x"cc"),
   933 => (x"cc",x"c0",x"9b",x"ff"),
   934 => (x"4a",x"66",x"cc",x"87"),
   935 => (x"cc",x"2a",x"b7",x"c8"),
   936 => (x"ff",x"c3",x"4b",x"66"),
   937 => (x"18",x"50",x"27",x"9b"),
   938 => (x"27",x"1e",x"00",x"00"),
   939 => (x"00",x"00",x"18",x"1c"),
   940 => (x"81",x"72",x"49",x"bf"),
   941 => (x"d6",x"27",x"1e",x"71"),
   942 => (x"0f",x"00",x"00",x"07"),
   943 => (x"98",x"70",x"86",x"c8"),
   944 => (x"87",x"c5",x"c0",x"05"),
   945 => (x"f0",x"c0",x"48",x"c0"),
   946 => (x"18",x"10",x"27",x"87"),
   947 => (x"02",x"bf",x"00",x"00"),
   948 => (x"73",x"87",x"d6",x"c0"),
   949 => (x"91",x"b7",x"c4",x"49"),
   950 => (x"00",x"18",x"50",x"27"),
   951 => (x"4c",x"69",x"81",x"00"),
   952 => (x"ff",x"ff",x"ff",x"cf"),
   953 => (x"ce",x"c0",x"9c",x"ff"),
   954 => (x"c2",x"49",x"73",x"87"),
   955 => (x"50",x"27",x"91",x"b7"),
   956 => (x"81",x"00",x"00",x"18"),
   957 => (x"74",x"4c",x"69",x"9f"),
   958 => (x"d6",x"ee",x"ff",x"48"),
   959 => (x"5b",x"5e",x"0e",x"87"),
   960 => (x"f4",x"0e",x"5d",x"5c"),
   961 => (x"76",x"4b",x"c0",x"86"),
   962 => (x"18",x"24",x"27",x"48"),
   963 => (x"78",x"bf",x"00",x"00"),
   964 => (x"28",x"27",x"80",x"c4"),
   965 => (x"bf",x"00",x"00",x"18"),
   966 => (x"18",x"10",x"27",x"78"),
   967 => (x"02",x"bf",x"00",x"00"),
   968 => (x"27",x"87",x"cc",x"c0"),
   969 => (x"00",x"00",x"18",x"08"),
   970 => (x"31",x"c4",x"49",x"bf"),
   971 => (x"27",x"87",x"c9",x"c0"),
   972 => (x"00",x"00",x"18",x"2c"),
   973 => (x"31",x"c4",x"49",x"bf"),
   974 => (x"c0",x"59",x"a6",x"cc"),
   975 => (x"48",x"66",x"c8",x"4d"),
   976 => (x"c3",x"06",x"a8",x"c0"),
   977 => (x"49",x"75",x"87",x"c3"),
   978 => (x"99",x"71",x"99",x"cf"),
   979 => (x"87",x"e2",x"c0",x"05"),
   980 => (x"00",x"18",x"50",x"27"),
   981 => (x"66",x"c8",x"1e",x"00"),
   982 => (x"80",x"c1",x"48",x"49"),
   983 => (x"71",x"58",x"a6",x"cc"),
   984 => (x"07",x"d6",x"27",x"1e"),
   985 => (x"c8",x"0f",x"00",x"00"),
   986 => (x"18",x"50",x"27",x"86"),
   987 => (x"c0",x"4b",x"00",x"00"),
   988 => (x"e0",x"c0",x"87",x"c3"),
   989 => (x"49",x"6b",x"97",x"83"),
   990 => (x"c2",x"02",x"99",x"71"),
   991 => (x"6b",x"97",x"87",x"c2"),
   992 => (x"a9",x"e5",x"c3",x"49"),
   993 => (x"87",x"f8",x"c1",x"02"),
   994 => (x"81",x"cb",x"49",x"73"),
   995 => (x"d8",x"49",x"69",x"97"),
   996 => (x"05",x"99",x"71",x"99"),
   997 => (x"73",x"87",x"e9",x"c1"),
   998 => (x"00",x"68",x"27",x"1e"),
   999 => (x"c4",x"0f",x"00",x"00"),
  1000 => (x"c0",x"1e",x"cb",x"86"),
  1001 => (x"73",x"1e",x"66",x"e4"),
  1002 => (x"0a",x"43",x"27",x"1e"),
  1003 => (x"cc",x"0f",x"00",x"00"),
  1004 => (x"05",x"98",x"70",x"86"),
  1005 => (x"73",x"87",x"c9",x"c1"),
  1006 => (x"dc",x"82",x"dc",x"4a"),
  1007 => (x"81",x"c4",x"49",x"66"),
  1008 => (x"4a",x"73",x"79",x"6a"),
  1009 => (x"66",x"dc",x"82",x"da"),
  1010 => (x"9f",x"81",x"c8",x"49"),
  1011 => (x"79",x"70",x"48",x"6a"),
  1012 => (x"10",x"27",x"4c",x"71"),
  1013 => (x"bf",x"00",x"00",x"18"),
  1014 => (x"87",x"d2",x"c0",x"02"),
  1015 => (x"81",x"d4",x"49",x"73"),
  1016 => (x"c0",x"49",x"69",x"9f"),
  1017 => (x"71",x"99",x"ff",x"ff"),
  1018 => (x"c0",x"32",x"d0",x"4a"),
  1019 => (x"4a",x"c0",x"87",x"c2"),
  1020 => (x"80",x"6c",x"48",x"72"),
  1021 => (x"66",x"dc",x"7c",x"70"),
  1022 => (x"c1",x"78",x"c0",x"48"),
  1023 => (x"87",x"c9",x"c1",x"48"),
  1024 => (x"66",x"c8",x"85",x"c1"),
  1025 => (x"fd",x"fc",x"04",x"ad"),
  1026 => (x"18",x"10",x"27",x"87"),
  1027 => (x"02",x"bf",x"00",x"00"),
  1028 => (x"6e",x"87",x"f4",x"c0"),
  1029 => (x"0e",x"7b",x"27",x"1e"),
  1030 => (x"c4",x"0f",x"00",x"00"),
  1031 => (x"58",x"a6",x"c4",x"86"),
  1032 => (x"ff",x"cf",x"49",x"6e"),
  1033 => (x"99",x"f8",x"ff",x"ff"),
  1034 => (x"da",x"c0",x"02",x"a9"),
  1035 => (x"c2",x"49",x"6e",x"87"),
  1036 => (x"18",x"08",x"27",x"89"),
  1037 => (x"91",x"bf",x"00",x"00"),
  1038 => (x"00",x"18",x"20",x"27"),
  1039 => (x"71",x"48",x"bf",x"00"),
  1040 => (x"58",x"a6",x"c8",x"80"),
  1041 => (x"c0",x"87",x"f4",x"fb"),
  1042 => (x"ff",x"8e",x"f4",x"48"),
  1043 => (x"0e",x"87",x"c2",x"e9"),
  1044 => (x"c8",x"0e",x"5b",x"5e"),
  1045 => (x"c1",x"49",x"bf",x"66"),
  1046 => (x"09",x"66",x"c8",x"81"),
  1047 => (x"0c",x"27",x"09",x"79"),
  1048 => (x"bf",x"00",x"00",x"18"),
  1049 => (x"05",x"99",x"71",x"99"),
  1050 => (x"c8",x"87",x"d3",x"c0"),
  1051 => (x"83",x"c8",x"4b",x"66"),
  1052 => (x"7b",x"27",x"1e",x"6b"),
  1053 => (x"0f",x"00",x"00",x"0e"),
  1054 => (x"49",x"70",x"86",x"c4"),
  1055 => (x"48",x"c1",x"7b",x"71"),
  1056 => (x"87",x"d1",x"e8",x"ff"),
  1057 => (x"27",x"0e",x"5e",x"0e"),
  1058 => (x"00",x"00",x"18",x"20"),
  1059 => (x"66",x"c4",x"49",x"bf"),
  1060 => (x"6a",x"82",x"c8",x"4a"),
  1061 => (x"27",x"8a",x"c2",x"4a"),
  1062 => (x"00",x"00",x"18",x"08"),
  1063 => (x"81",x"72",x"92",x"bf"),
  1064 => (x"00",x"18",x"0c",x"27"),
  1065 => (x"c4",x"4a",x"bf",x"00"),
  1066 => (x"72",x"9a",x"bf",x"66"),
  1067 => (x"1e",x"66",x"c8",x"81"),
  1068 => (x"d6",x"27",x"1e",x"71"),
  1069 => (x"0f",x"00",x"00",x"07"),
  1070 => (x"98",x"70",x"86",x"c8"),
  1071 => (x"87",x"c5",x"c0",x"05"),
  1072 => (x"c2",x"c0",x"48",x"c0"),
  1073 => (x"ff",x"48",x"c1",x"87"),
  1074 => (x"0e",x"87",x"cc",x"e7"),
  1075 => (x"0e",x"5c",x"5b",x"5e"),
  1076 => (x"27",x"1e",x"66",x"cc"),
  1077 => (x"00",x"00",x"18",x"40"),
  1078 => (x"0e",x"fd",x"27",x"1e"),
  1079 => (x"c8",x"0f",x"00",x"00"),
  1080 => (x"02",x"98",x"70",x"86"),
  1081 => (x"27",x"87",x"e4",x"c1"),
  1082 => (x"00",x"00",x"18",x"44"),
  1083 => (x"ff",x"c7",x"49",x"bf"),
  1084 => (x"71",x"29",x"c9",x"81"),
  1085 => (x"27",x"4b",x"c0",x"4c"),
  1086 => (x"00",x"00",x"11",x"67"),
  1087 => (x"00",x"68",x"27",x"1e"),
  1088 => (x"c4",x"0f",x"00",x"00"),
  1089 => (x"ac",x"b7",x"c0",x"86"),
  1090 => (x"87",x"d5",x"c1",x"06"),
  1091 => (x"27",x"1e",x"66",x"d0"),
  1092 => (x"00",x"00",x"18",x"40"),
  1093 => (x"10",x"84",x"27",x"1e"),
  1094 => (x"c8",x"0f",x"00",x"00"),
  1095 => (x"05",x"98",x"70",x"86"),
  1096 => (x"c0",x"87",x"c5",x"c0"),
  1097 => (x"87",x"fb",x"c0",x"48"),
  1098 => (x"00",x"18",x"40",x"27"),
  1099 => (x"4f",x"27",x"1e",x"00"),
  1100 => (x"0f",x"00",x"00",x"10"),
  1101 => (x"66",x"d0",x"86",x"c4"),
  1102 => (x"80",x"c0",x"c8",x"48"),
  1103 => (x"c1",x"58",x"a6",x"d4"),
  1104 => (x"ab",x"b7",x"74",x"83"),
  1105 => (x"87",x"c4",x"ff",x"04"),
  1106 => (x"cc",x"87",x"d6",x"c0"),
  1107 => (x"80",x"27",x"1e",x"66"),
  1108 => (x"1e",x"00",x"00",x"11"),
  1109 => (x"00",x"00",x"9c",x"27"),
  1110 => (x"86",x"c8",x"0f",x"00"),
  1111 => (x"c2",x"c0",x"48",x"c0"),
  1112 => (x"ff",x"48",x"c1",x"87"),
  1113 => (x"4f",x"87",x"ec",x"e4"),
  1114 => (x"65",x"6e",x"65",x"70"),
  1115 => (x"69",x"66",x"20",x"64"),
  1116 => (x"20",x"2c",x"65",x"6c"),
  1117 => (x"64",x"61",x"6f",x"6c"),
  1118 => (x"2e",x"67",x"6e",x"69"),
  1119 => (x"00",x"0a",x"2e",x"2e"),
  1120 => (x"27",x"6e",x"61",x"43"),
  1121 => (x"70",x"6f",x"20",x"74"),
  1122 => (x"25",x"20",x"6e",x"65"),
  1123 => (x"0e",x"00",x"0a",x"73"),
  1124 => (x"66",x"c4",x"0e",x"5e"),
  1125 => (x"c3",x"29",x"d8",x"49"),
  1126 => (x"66",x"c4",x"99",x"ff"),
  1127 => (x"cf",x"2a",x"c8",x"4a"),
  1128 => (x"72",x"9a",x"c0",x"fc"),
  1129 => (x"4a",x"66",x"c4",x"b1"),
  1130 => (x"ff",x"c0",x"32",x"c8"),
  1131 => (x"9a",x"c0",x"c0",x"f0"),
  1132 => (x"66",x"c4",x"b1",x"72"),
  1133 => (x"ff",x"32",x"d8",x"4a"),
  1134 => (x"c0",x"c0",x"c0",x"c0"),
  1135 => (x"71",x"b1",x"72",x"9a"),
  1136 => (x"c6",x"c0",x"c0",x"48"),
  1137 => (x"26",x"4d",x"26",x"87"),
  1138 => (x"26",x"4b",x"26",x"4c"),
  1139 => (x"0e",x"5e",x"0e",x"4f"),
  1140 => (x"c8",x"4a",x"66",x"c4"),
  1141 => (x"9a",x"ff",x"c3",x"2a"),
  1142 => (x"9a",x"ff",x"ff",x"cf"),
  1143 => (x"c8",x"49",x"66",x"c4"),
  1144 => (x"c0",x"fc",x"cf",x"31"),
  1145 => (x"cf",x"b1",x"72",x"99"),
  1146 => (x"71",x"99",x"ff",x"ff"),
  1147 => (x"da",x"ff",x"ff",x"48"),
  1148 => (x"0e",x"5e",x"0e",x"87"),
  1149 => (x"d0",x"49",x"66",x"c4"),
  1150 => (x"ff",x"ff",x"cf",x"29"),
  1151 => (x"4a",x"66",x"c4",x"99"),
  1152 => (x"c0",x"f0",x"32",x"d0"),
  1153 => (x"b1",x"72",x"9a",x"c0"),
  1154 => (x"fe",x"ff",x"48",x"71"),
  1155 => (x"73",x"1e",x"87",x"fd"),
  1156 => (x"c0",x"c0",x"d0",x"1e"),
  1157 => (x"73",x"4b",x"c0",x"c0"),
  1158 => (x"87",x"fd",x"ff",x"0f"),
  1159 => (x"87",x"c4",x"c0",x"c0"),
  1160 => (x"4c",x"26",x"4d",x"26"),
  1161 => (x"4f",x"26",x"4b",x"26"),
  1162 => (x"49",x"66",x"c8",x"1e"),
  1163 => (x"c0",x"99",x"df",x"c3"),
  1164 => (x"b7",x"c0",x"89",x"f7"),
  1165 => (x"c3",x"c0",x"03",x"a9"),
  1166 => (x"81",x"e7",x"c0",x"87"),
  1167 => (x"c4",x"48",x"66",x"c4"),
  1168 => (x"58",x"a6",x"c8",x"30"),
  1169 => (x"71",x"48",x"66",x"c4"),
  1170 => (x"58",x"a6",x"c8",x"b0"),
  1171 => (x"ff",x"48",x"66",x"c4"),
  1172 => (x"0e",x"87",x"d3",x"ff"),
  1173 => (x"0e",x"5c",x"5b",x"5e"),
  1174 => (x"c0",x"c0",x"c0",x"d0"),
  1175 => (x"50",x"27",x"4c",x"c0"),
  1176 => (x"bf",x"00",x"00",x"1a"),
  1177 => (x"27",x"80",x"c1",x"48"),
  1178 => (x"00",x"00",x"1a",x"54"),
  1179 => (x"66",x"cc",x"97",x"58"),
  1180 => (x"81",x"c0",x"fe",x"49"),
  1181 => (x"a9",x"d3",x"c1",x"b9"),
  1182 => (x"87",x"e9",x"c0",x"05"),
  1183 => (x"00",x"1a",x"50",x"27"),
  1184 => (x"78",x"c0",x"48",x"00"),
  1185 => (x"00",x"1a",x"54",x"27"),
  1186 => (x"78",x"c0",x"48",x"00"),
  1187 => (x"00",x"1a",x"5c",x"27"),
  1188 => (x"78",x"c0",x"48",x"00"),
  1189 => (x"00",x"1a",x"60",x"27"),
  1190 => (x"78",x"c0",x"48",x"00"),
  1191 => (x"c1",x"48",x"c0",x"ff"),
  1192 => (x"e3",x"c9",x"78",x"d3"),
  1193 => (x"1a",x"50",x"27",x"87"),
  1194 => (x"48",x"bf",x"00",x"00"),
  1195 => (x"c1",x"05",x"a8",x"c1"),
  1196 => (x"c0",x"ff",x"87",x"d4"),
  1197 => (x"78",x"f4",x"c1",x"48"),
  1198 => (x"49",x"66",x"cc",x"97"),
  1199 => (x"b9",x"81",x"c0",x"fe"),
  1200 => (x"60",x"27",x"1e",x"71"),
  1201 => (x"bf",x"00",x"00",x"1a"),
  1202 => (x"12",x"28",x"27",x"1e"),
  1203 => (x"c8",x"0f",x"00",x"00"),
  1204 => (x"1a",x"64",x"27",x"86"),
  1205 => (x"27",x"58",x"00",x"00"),
  1206 => (x"00",x"00",x"1a",x"60"),
  1207 => (x"b7",x"c3",x"4a",x"bf"),
  1208 => (x"c6",x"c0",x"06",x"aa"),
  1209 => (x"72",x"48",x"ca",x"87"),
  1210 => (x"72",x"4a",x"70",x"88"),
  1211 => (x"71",x"81",x"c1",x"49"),
  1212 => (x"27",x"30",x"c1",x"48"),
  1213 => (x"00",x"00",x"1a",x"5c"),
  1214 => (x"c0",x"48",x"72",x"58"),
  1215 => (x"c0",x"ff",x"80",x"f0"),
  1216 => (x"c8",x"08",x"78",x"08"),
  1217 => (x"60",x"27",x"87",x"c2"),
  1218 => (x"bf",x"00",x"00",x"1a"),
  1219 => (x"a8",x"b7",x"c9",x"48"),
  1220 => (x"87",x"f4",x"c7",x"01"),
  1221 => (x"00",x"1a",x"60",x"27"),
  1222 => (x"c0",x"48",x"bf",x"00"),
  1223 => (x"c7",x"06",x"a8",x"b7"),
  1224 => (x"60",x"27",x"87",x"e6"),
  1225 => (x"bf",x"00",x"00",x"1a"),
  1226 => (x"80",x"f0",x"c0",x"48"),
  1227 => (x"78",x"08",x"c0",x"ff"),
  1228 => (x"1a",x"50",x"27",x"08"),
  1229 => (x"48",x"bf",x"00",x"00"),
  1230 => (x"01",x"a8",x"b7",x"c3"),
  1231 => (x"97",x"87",x"e2",x"c0"),
  1232 => (x"fe",x"49",x"66",x"cc"),
  1233 => (x"71",x"b9",x"81",x"c0"),
  1234 => (x"1a",x"5c",x"27",x"1e"),
  1235 => (x"1e",x"bf",x"00",x"00"),
  1236 => (x"00",x"12",x"28",x"27"),
  1237 => (x"86",x"c8",x"0f",x"00"),
  1238 => (x"00",x"1a",x"60",x"27"),
  1239 => (x"e7",x"c6",x"58",x"00"),
  1240 => (x"1a",x"58",x"27",x"87"),
  1241 => (x"49",x"bf",x"00",x"00"),
  1242 => (x"50",x"27",x"81",x"c3"),
  1243 => (x"bf",x"00",x"00",x"1a"),
  1244 => (x"c0",x"04",x"a9",x"b7"),
  1245 => (x"cc",x"97",x"87",x"ea"),
  1246 => (x"c0",x"fe",x"49",x"66"),
  1247 => (x"1e",x"71",x"b9",x"81"),
  1248 => (x"00",x"1a",x"54",x"27"),
  1249 => (x"27",x"1e",x"bf",x"00"),
  1250 => (x"00",x"00",x"12",x"28"),
  1251 => (x"27",x"86",x"c8",x"0f"),
  1252 => (x"00",x"00",x"1a",x"58"),
  1253 => (x"1a",x"64",x"27",x"58"),
  1254 => (x"c1",x"48",x"00",x"00"),
  1255 => (x"87",x"e8",x"c5",x"78"),
  1256 => (x"00",x"1a",x"60",x"27"),
  1257 => (x"c0",x"48",x"bf",x"00"),
  1258 => (x"c3",x"06",x"a8",x"b7"),
  1259 => (x"60",x"27",x"87",x"c4"),
  1260 => (x"bf",x"00",x"00",x"1a"),
  1261 => (x"a8",x"b7",x"c3",x"48"),
  1262 => (x"87",x"f6",x"c2",x"01"),
  1263 => (x"00",x"1a",x"5c",x"27"),
  1264 => (x"c1",x"49",x"bf",x"00"),
  1265 => (x"50",x"27",x"81",x"31"),
  1266 => (x"bf",x"00",x"00",x"1a"),
  1267 => (x"c1",x"04",x"a9",x"b7"),
  1268 => (x"cc",x"97",x"87",x"fa"),
  1269 => (x"c0",x"fe",x"49",x"66"),
  1270 => (x"1e",x"71",x"b9",x"81"),
  1271 => (x"00",x"1a",x"68",x"27"),
  1272 => (x"27",x"1e",x"bf",x"00"),
  1273 => (x"00",x"00",x"12",x"28"),
  1274 => (x"27",x"86",x"c8",x"0f"),
  1275 => (x"00",x"00",x"1a",x"6c"),
  1276 => (x"1a",x"64",x"27",x"58"),
  1277 => (x"49",x"bf",x"00",x"00"),
  1278 => (x"68",x"27",x"89",x"c1"),
  1279 => (x"59",x"00",x"00",x"1a"),
  1280 => (x"03",x"a9",x"b7",x"c0"),
  1281 => (x"27",x"87",x"c1",x"c4"),
  1282 => (x"00",x"00",x"1a",x"54"),
  1283 => (x"68",x"27",x"49",x"bf"),
  1284 => (x"97",x"00",x"00",x"1a"),
  1285 => (x"ff",x"c3",x"51",x"bf"),
  1286 => (x"1a",x"54",x"27",x"98"),
  1287 => (x"49",x"bf",x"00",x"00"),
  1288 => (x"58",x"27",x"81",x"c1"),
  1289 => (x"59",x"00",x"00",x"1a"),
  1290 => (x"00",x"1a",x"6c",x"27"),
  1291 => (x"a9",x"b7",x"bf",x"00"),
  1292 => (x"87",x"cd",x"c0",x"06"),
  1293 => (x"00",x"1a",x"6c",x"27"),
  1294 => (x"54",x"27",x"48",x"00"),
  1295 => (x"bf",x"00",x"00",x"1a"),
  1296 => (x"1a",x"64",x"27",x"78"),
  1297 => (x"c1",x"48",x"00",x"00"),
  1298 => (x"87",x"fc",x"c2",x"78"),
  1299 => (x"00",x"1a",x"64",x"27"),
  1300 => (x"c2",x"05",x"bf",x"00"),
  1301 => (x"68",x"27",x"87",x"f2"),
  1302 => (x"bf",x"00",x"00",x"1a"),
  1303 => (x"27",x"31",x"c4",x"49"),
  1304 => (x"00",x"00",x"1a",x"6c"),
  1305 => (x"1a",x"54",x"27",x"59"),
  1306 => (x"09",x"bf",x"00",x"00"),
  1307 => (x"c2",x"09",x"79",x"97"),
  1308 => (x"60",x"27",x"87",x"d6"),
  1309 => (x"bf",x"00",x"00",x"1a"),
  1310 => (x"a8",x"b7",x"c7",x"48"),
  1311 => (x"87",x"f9",x"c1",x"04"),
  1312 => (x"f4",x"fe",x"4b",x"c0"),
  1313 => (x"27",x"78",x"c1",x"48"),
  1314 => (x"00",x"00",x"1a",x"6c"),
  1315 => (x"1e",x"74",x"1e",x"bf"),
  1316 => (x"00",x"17",x"bb",x"27"),
  1317 => (x"9c",x"27",x"1e",x"00"),
  1318 => (x"0f",x"00",x"00",x"00"),
  1319 => (x"58",x"27",x"86",x"cc"),
  1320 => (x"5c",x"00",x"00",x"1a"),
  1321 => (x"00",x"1a",x"54",x"27"),
  1322 => (x"27",x"48",x"bf",x"00"),
  1323 => (x"00",x"00",x"1a",x"6c"),
  1324 => (x"03",x"a8",x"b7",x"bf"),
  1325 => (x"27",x"87",x"e3",x"c0"),
  1326 => (x"00",x"00",x"1a",x"54"),
  1327 => (x"27",x"83",x"bf",x"bf"),
  1328 => (x"00",x"00",x"1a",x"54"),
  1329 => (x"81",x"c4",x"49",x"bf"),
  1330 => (x"00",x"1a",x"58",x"27"),
  1331 => (x"6c",x"27",x"59",x"00"),
  1332 => (x"bf",x"00",x"00",x"1a"),
  1333 => (x"ff",x"04",x"a9",x"b7"),
  1334 => (x"1e",x"73",x"87",x"dd"),
  1335 => (x"00",x"17",x"da",x"27"),
  1336 => (x"9c",x"27",x"1e",x"00"),
  1337 => (x"0f",x"00",x"00",x"00"),
  1338 => (x"c0",x"ff",x"86",x"c8"),
  1339 => (x"78",x"c2",x"c1",x"48"),
  1340 => (x"00",x"12",x"0e",x"27"),
  1341 => (x"cf",x"c0",x"0f",x"00"),
  1342 => (x"1a",x"60",x"27",x"87"),
  1343 => (x"48",x"bf",x"00",x"00"),
  1344 => (x"ff",x"80",x"f0",x"c0"),
  1345 => (x"08",x"78",x"08",x"c0"),
  1346 => (x"87",x"d6",x"f4",x"ff"),
  1347 => (x"5c",x"5b",x"5e",x"0e"),
  1348 => (x"0e",x"27",x"0e",x"5d"),
  1349 => (x"1e",x"00",x"00",x"16"),
  1350 => (x"00",x"00",x"68",x"27"),
  1351 => (x"86",x"c4",x"0f",x"00"),
  1352 => (x"00",x"04",x"df",x"27"),
  1353 => (x"98",x"70",x"0f",x"00"),
  1354 => (x"87",x"d1",x"c0",x"02"),
  1355 => (x"00",x"0a",x"99",x"27"),
  1356 => (x"98",x"70",x"0f",x"00"),
  1357 => (x"87",x"c5",x"c0",x"02"),
  1358 => (x"c2",x"c0",x"49",x"c1"),
  1359 => (x"71",x"49",x"c0",x"87"),
  1360 => (x"16",x"24",x"27",x"4d"),
  1361 => (x"27",x"1e",x"00",x"00"),
  1362 => (x"00",x"00",x"00",x"68"),
  1363 => (x"27",x"86",x"c4",x"0f"),
  1364 => (x"00",x"00",x"1a",x"6c"),
  1365 => (x"c0",x"78",x"c0",x"48"),
  1366 => (x"45",x"27",x"1e",x"ee"),
  1367 => (x"0f",x"00",x"00",x"00"),
  1368 => (x"f4",x"c3",x"86",x"c4"),
  1369 => (x"ff",x"4a",x"ff",x"c8"),
  1370 => (x"74",x"4c",x"bf",x"c0"),
  1371 => (x"99",x"c0",x"c8",x"49"),
  1372 => (x"c1",x"02",x"99",x"71"),
  1373 => (x"4b",x"74",x"87",x"df"),
  1374 => (x"db",x"9b",x"ff",x"c3"),
  1375 => (x"c5",x"c1",x"05",x"ab"),
  1376 => (x"02",x"9d",x"75",x"87"),
  1377 => (x"d0",x"87",x"f1",x"c0"),
  1378 => (x"c0",x"c0",x"c0",x"c0"),
  1379 => (x"15",x"f2",x"27",x"1e"),
  1380 => (x"27",x"1e",x"00",x"00"),
  1381 => (x"00",x"00",x"10",x"cb"),
  1382 => (x"70",x"86",x"c8",x"0f"),
  1383 => (x"d7",x"c0",x"02",x"98"),
  1384 => (x"15",x"e6",x"27",x"87"),
  1385 => (x"27",x"1e",x"00",x"00"),
  1386 => (x"00",x"00",x"00",x"68"),
  1387 => (x"27",x"86",x"c4",x"0f"),
  1388 => (x"00",x"00",x"12",x"0e"),
  1389 => (x"87",x"ce",x"c0",x"0f"),
  1390 => (x"00",x"15",x"fe",x"27"),
  1391 => (x"68",x"27",x"1e",x"00"),
  1392 => (x"0f",x"00",x"00",x"00"),
  1393 => (x"1e",x"73",x"86",x"c4"),
  1394 => (x"00",x"12",x"53",x"27"),
  1395 => (x"86",x"c4",x"0f",x"00"),
  1396 => (x"c0",x"c9",x"f4",x"c3"),
  1397 => (x"c1",x"49",x"72",x"4a"),
  1398 => (x"05",x"99",x"71",x"8a"),
  1399 => (x"fd",x"87",x"c8",x"fe"),
  1400 => (x"f0",x"ff",x"87",x"f5"),
  1401 => (x"6f",x"42",x"87",x"fa"),
  1402 => (x"6e",x"69",x"74",x"6f"),
  1403 => (x"2e",x"2e",x"2e",x"67"),
  1404 => (x"4f",x"42",x"00",x"0a"),
  1405 => (x"33",x"38",x"54",x"4f"),
  1406 => (x"49",x"42",x"20",x"32"),
  1407 => (x"44",x"53",x"00",x"4e"),
  1408 => (x"6f",x"6f",x"62",x"20"),
  1409 => (x"61",x"66",x"20",x"74"),
  1410 => (x"64",x"65",x"6c",x"69"),
  1411 => (x"6e",x"49",x"00",x"0a"),
  1412 => (x"61",x"69",x"74",x"69"),
  1413 => (x"69",x"7a",x"69",x"6c"),
  1414 => (x"53",x"20",x"67",x"6e"),
  1415 => (x"61",x"63",x"20",x"44"),
  1416 => (x"00",x"0a",x"64",x"72"),
  1417 => (x"33",x"32",x"53",x"52"),
  1418 => (x"6f",x"62",x"20",x"32"),
  1419 => (x"2d",x"20",x"74",x"6f"),
  1420 => (x"65",x"72",x"70",x"20"),
  1421 => (x"45",x"20",x"73",x"73"),
  1422 => (x"74",x"20",x"43",x"53"),
  1423 => (x"6f",x"62",x"20",x"6f"),
  1424 => (x"66",x"20",x"74",x"6f"),
  1425 => (x"20",x"6d",x"6f",x"72"),
  1426 => (x"00",x"2e",x"44",x"53"),
  1427 => (x"00",x"44",x"4d",x"43"),
  1428 => (x"64",x"61",x"65",x"52"),
  1429 => (x"20",x"66",x"6f",x"20"),
  1430 => (x"20",x"52",x"42",x"4d"),
  1431 => (x"6c",x"69",x"61",x"66"),
  1432 => (x"00",x"0a",x"64",x"65"),
  1433 => (x"70",x"20",x"6f",x"4e"),
  1434 => (x"69",x"74",x"72",x"61"),
  1435 => (x"6e",x"6f",x"69",x"74"),
  1436 => (x"67",x"69",x"73",x"20"),
  1437 => (x"75",x"74",x"61",x"6e"),
  1438 => (x"66",x"20",x"65",x"72"),
  1439 => (x"64",x"6e",x"75",x"6f"),
  1440 => (x"42",x"4d",x"00",x"0a"),
  1441 => (x"7a",x"69",x"73",x"52"),
  1442 => (x"25",x"20",x"3a",x"65"),
  1443 => (x"70",x"20",x"2c",x"64"),
  1444 => (x"69",x"74",x"72",x"61"),
  1445 => (x"6e",x"6f",x"69",x"74"),
  1446 => (x"65",x"7a",x"69",x"73"),
  1447 => (x"64",x"25",x"20",x"3a"),
  1448 => (x"66",x"6f",x"20",x"2c"),
  1449 => (x"74",x"65",x"73",x"66"),
  1450 => (x"20",x"66",x"6f",x"20"),
  1451 => (x"3a",x"67",x"69",x"73"),
  1452 => (x"2c",x"64",x"25",x"20"),
  1453 => (x"67",x"69",x"73",x"20"),
  1454 => (x"25",x"78",x"30",x"20"),
  1455 => (x"52",x"00",x"0a",x"78"),
  1456 => (x"69",x"64",x"61",x"65"),
  1457 => (x"62",x"20",x"67",x"6e"),
  1458 => (x"20",x"74",x"6f",x"6f"),
  1459 => (x"74",x"63",x"65",x"73"),
  1460 => (x"25",x"20",x"72",x"6f"),
  1461 => (x"52",x"00",x"0a",x"64"),
  1462 => (x"20",x"64",x"61",x"65"),
  1463 => (x"74",x"6f",x"6f",x"62"),
  1464 => (x"63",x"65",x"73",x"20"),
  1465 => (x"20",x"72",x"6f",x"74"),
  1466 => (x"6d",x"6f",x"72",x"66"),
  1467 => (x"72",x"69",x"66",x"20"),
  1468 => (x"70",x"20",x"74",x"73"),
  1469 => (x"69",x"74",x"72",x"61"),
  1470 => (x"6e",x"6f",x"69",x"74"),
  1471 => (x"6e",x"55",x"00",x"0a"),
  1472 => (x"70",x"70",x"75",x"73"),
  1473 => (x"65",x"74",x"72",x"6f"),
  1474 => (x"61",x"70",x"20",x"64"),
  1475 => (x"74",x"69",x"74",x"72"),
  1476 => (x"20",x"6e",x"6f",x"69"),
  1477 => (x"65",x"70",x"79",x"74"),
  1478 => (x"46",x"00",x"0d",x"21"),
  1479 => (x"32",x"33",x"54",x"41"),
  1480 => (x"00",x"20",x"20",x"20"),
  1481 => (x"64",x"61",x"65",x"52"),
  1482 => (x"20",x"67",x"6e",x"69"),
  1483 => (x"0a",x"52",x"42",x"4d"),
  1484 => (x"52",x"42",x"4d",x"00"),
  1485 => (x"63",x"75",x"73",x"20"),
  1486 => (x"73",x"73",x"65",x"63"),
  1487 => (x"6c",x"6c",x"75",x"66"),
  1488 => (x"65",x"72",x"20",x"79"),
  1489 => (x"00",x"0a",x"64",x"61"),
  1490 => (x"31",x"54",x"41",x"46"),
  1491 => (x"20",x"20",x"20",x"36"),
  1492 => (x"54",x"41",x"46",x"00"),
  1493 => (x"20",x"20",x"32",x"33"),
  1494 => (x"61",x"50",x"00",x"20"),
  1495 => (x"74",x"69",x"74",x"72"),
  1496 => (x"63",x"6e",x"6f",x"69"),
  1497 => (x"74",x"6e",x"75",x"6f"),
  1498 => (x"0a",x"64",x"25",x"20"),
  1499 => (x"6e",x"75",x"48",x"00"),
  1500 => (x"67",x"6e",x"69",x"74"),
  1501 => (x"72",x"6f",x"66",x"20"),
  1502 => (x"6c",x"69",x"66",x"20"),
  1503 => (x"73",x"79",x"73",x"65"),
  1504 => (x"0a",x"6d",x"65",x"74"),
  1505 => (x"54",x"41",x"46",x"00"),
  1506 => (x"20",x"20",x"32",x"33"),
  1507 => (x"41",x"46",x"00",x"20"),
  1508 => (x"20",x"36",x"31",x"54"),
  1509 => (x"43",x"00",x"20",x"20"),
  1510 => (x"74",x"73",x"75",x"6c"),
  1511 => (x"73",x"20",x"72",x"65"),
  1512 => (x"3a",x"65",x"7a",x"69"),
  1513 => (x"2c",x"64",x"25",x"20"),
  1514 => (x"75",x"6c",x"43",x"20"),
  1515 => (x"72",x"65",x"74",x"73"),
  1516 => (x"73",x"61",x"6d",x"20"),
  1517 => (x"25",x"20",x"2c",x"6b"),
  1518 => (x"43",x"00",x"0a",x"64"),
  1519 => (x"6b",x"63",x"65",x"68"),
  1520 => (x"6d",x"6d",x"75",x"73"),
  1521 => (x"20",x"67",x"6e",x"69"),
  1522 => (x"6d",x"6f",x"72",x"66"),
  1523 => (x"20",x"64",x"25",x"20"),
  1524 => (x"25",x"20",x"6f",x"74"),
  1525 => (x"2e",x"2e",x"2e",x"64"),
  1526 => (x"64",x"25",x"00",x"20"),
  1527 => (x"64",x"25",x"00",x"0a"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
