
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"2c",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"29"),
    10 => (x"87",x"fd",x"00",x"4f"),
    11 => (x"c4",x"f2",x"c3",x"4f"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"c4",x"f2",x"c3"),
    14 => (x"48",x"cc",x"cf",x"c1"),
    15 => (x"03",x"89",x"d0",x"89"),
    16 => (x"40",x"40",x"40",x"c0"),
    17 => (x"d0",x"87",x"f6",x"40"),
    18 => (x"50",x"c0",x"05",x"81"),
    19 => (x"f9",x"05",x"89",x"c1"),
    20 => (x"c9",x"cf",x"c1",x"87"),
    21 => (x"c9",x"cf",x"c1",x"4d"),
    22 => (x"02",x"ad",x"74",x"4c"),
    23 => (x"0f",x"24",x"87",x"c4"),
    24 => (x"ed",x"cd",x"87",x"f7"),
    25 => (x"c9",x"cf",x"c1",x"87"),
    26 => (x"c9",x"cf",x"c1",x"4d"),
    27 => (x"02",x"ad",x"74",x"4c"),
    28 => (x"8c",x"c4",x"87",x"c6"),
    29 => (x"87",x"f5",x"0f",x"6c"),
    30 => (x"0e",x"87",x"fd",x"00"),
    31 => (x"5d",x"5c",x"5b",x"5e"),
    32 => (x"71",x"86",x"fc",x"0e"),
    33 => (x"66",x"e0",x"c0",x"4a"),
    34 => (x"cc",x"cf",x"c1",x"4c"),
    35 => (x"72",x"7e",x"c0",x"4b"),
    36 => (x"87",x"ce",x"05",x"9a"),
    37 => (x"4b",x"cd",x"cf",x"c1"),
    38 => (x"48",x"cc",x"cf",x"c1"),
    39 => (x"c1",x"50",x"f0",x"c0"),
    40 => (x"9a",x"72",x"87",x"d1"),
    41 => (x"87",x"e8",x"c0",x"02"),
    42 => (x"72",x"4d",x"66",x"d4"),
    43 => (x"75",x"49",x"72",x"1e"),
    44 => (x"87",x"f9",x"ca",x"4a"),
    45 => (x"e4",x"c4",x"4a",x"26"),
    46 => (x"71",x"53",x"11",x"81"),
    47 => (x"75",x"49",x"72",x"1e"),
    48 => (x"87",x"e9",x"ca",x"4a"),
    49 => (x"49",x"26",x"4a",x"70"),
    50 => (x"9a",x"72",x"8c",x"c1"),
    51 => (x"87",x"db",x"ff",x"05"),
    52 => (x"06",x"ac",x"b7",x"c0"),
    53 => (x"e4",x"c0",x"87",x"dd"),
    54 => (x"87",x"c5",x"02",x"66"),
    55 => (x"c3",x"4a",x"f0",x"c0"),
    56 => (x"4a",x"e0",x"c0",x"87"),
    57 => (x"7a",x"97",x"0a",x"73"),
    58 => (x"8c",x"83",x"c1",x"0a"),
    59 => (x"01",x"ac",x"b7",x"c0"),
    60 => (x"c1",x"87",x"e3",x"ff"),
    61 => (x"02",x"ab",x"cc",x"cf"),
    62 => (x"66",x"d8",x"87",x"de"),
    63 => (x"1e",x"66",x"dc",x"4c"),
    64 => (x"6b",x"97",x"8b",x"c1"),
    65 => (x"c4",x"0f",x"74",x"49"),
    66 => (x"c1",x"48",x"6e",x"86"),
    67 => (x"58",x"a6",x"c4",x"80"),
    68 => (x"ab",x"cc",x"cf",x"c1"),
    69 => (x"87",x"e5",x"ff",x"05"),
    70 => (x"8e",x"fc",x"48",x"6e"),
    71 => (x"4c",x"26",x"4d",x"26"),
    72 => (x"4f",x"26",x"4b",x"26"),
    73 => (x"33",x"32",x"31",x"30"),
    74 => (x"37",x"36",x"35",x"34"),
    75 => (x"42",x"41",x"39",x"38"),
    76 => (x"46",x"45",x"44",x"43"),
    77 => (x"5b",x"5e",x"0e",x"00"),
    78 => (x"71",x"0e",x"5d",x"5c"),
    79 => (x"13",x"4d",x"ff",x"4b"),
    80 => (x"02",x"9c",x"74",x"4c"),
    81 => (x"85",x"c1",x"87",x"d8"),
    82 => (x"74",x"1e",x"66",x"d4"),
    83 => (x"0f",x"66",x"d4",x"49"),
    84 => (x"a8",x"74",x"86",x"c4"),
    85 => (x"13",x"87",x"c7",x"05"),
    86 => (x"05",x"9c",x"74",x"4c"),
    87 => (x"48",x"75",x"87",x"e8"),
    88 => (x"4c",x"26",x"4d",x"26"),
    89 => (x"4f",x"26",x"4b",x"26"),
    90 => (x"5c",x"5b",x"5e",x"0e"),
    91 => (x"86",x"e8",x"0e",x"5d"),
    92 => (x"c0",x"59",x"a6",x"c4"),
    93 => (x"c0",x"4d",x"66",x"e8"),
    94 => (x"48",x"a6",x"c8",x"4c"),
    95 => (x"97",x"6e",x"78",x"c0"),
    96 => (x"48",x"6e",x"4b",x"bf"),
    97 => (x"a6",x"c4",x"80",x"c1"),
    98 => (x"02",x"9b",x"73",x"58"),
    99 => (x"c8",x"87",x"d3",x"c6"),
   100 => (x"db",x"c5",x"02",x"66"),
   101 => (x"48",x"a6",x"cc",x"87"),
   102 => (x"80",x"fc",x"78",x"c0"),
   103 => (x"4a",x"73",x"78",x"c0"),
   104 => (x"02",x"8a",x"e0",x"c0"),
   105 => (x"c3",x"87",x"c6",x"c3"),
   106 => (x"c0",x"c3",x"02",x"8a"),
   107 => (x"02",x"8a",x"c2",x"87"),
   108 => (x"c2",x"87",x"e8",x"c2"),
   109 => (x"f4",x"c2",x"02",x"8a"),
   110 => (x"02",x"8a",x"c4",x"87"),
   111 => (x"c2",x"87",x"ee",x"c2"),
   112 => (x"e8",x"c2",x"02",x"8a"),
   113 => (x"02",x"8a",x"c3",x"87"),
   114 => (x"d4",x"87",x"ea",x"c2"),
   115 => (x"f6",x"c0",x"02",x"8a"),
   116 => (x"02",x"8a",x"d4",x"87"),
   117 => (x"ca",x"87",x"c0",x"c1"),
   118 => (x"f2",x"c0",x"02",x"8a"),
   119 => (x"02",x"8a",x"c1",x"87"),
   120 => (x"c1",x"87",x"e1",x"c1"),
   121 => (x"87",x"df",x"02",x"8a"),
   122 => (x"c1",x"02",x"8a",x"c8"),
   123 => (x"8a",x"c4",x"87",x"ce"),
   124 => (x"87",x"e3",x"c0",x"02"),
   125 => (x"c0",x"02",x"8a",x"c3"),
   126 => (x"8a",x"c2",x"87",x"e5"),
   127 => (x"c3",x"87",x"c8",x"02"),
   128 => (x"87",x"d3",x"02",x"8a"),
   129 => (x"cc",x"87",x"fa",x"c1"),
   130 => (x"78",x"ca",x"48",x"a6"),
   131 => (x"cc",x"87",x"d2",x"c2"),
   132 => (x"78",x"c2",x"48",x"a6"),
   133 => (x"cc",x"87",x"ca",x"c2"),
   134 => (x"78",x"d0",x"48",x"a6"),
   135 => (x"c0",x"87",x"c2",x"c2"),
   136 => (x"c0",x"1e",x"66",x"f0"),
   137 => (x"c4",x"1e",x"66",x"f0"),
   138 => (x"c4",x"4a",x"75",x"85"),
   139 => (x"fc",x"49",x"6a",x"8a"),
   140 => (x"86",x"c8",x"87",x"c3"),
   141 => (x"a4",x"71",x"49",x"70"),
   142 => (x"87",x"e5",x"c1",x"4c"),
   143 => (x"c1",x"48",x"a6",x"c8"),
   144 => (x"87",x"dd",x"c1",x"78"),
   145 => (x"1e",x"66",x"f0",x"c0"),
   146 => (x"4a",x"75",x"85",x"c4"),
   147 => (x"49",x"6a",x"8a",x"c4"),
   148 => (x"0f",x"66",x"f0",x"c0"),
   149 => (x"84",x"c1",x"86",x"c4"),
   150 => (x"c0",x"87",x"c6",x"c1"),
   151 => (x"c0",x"1e",x"66",x"f0"),
   152 => (x"f0",x"c0",x"49",x"e5"),
   153 => (x"86",x"c4",x"0f",x"66"),
   154 => (x"f4",x"c0",x"84",x"c1"),
   155 => (x"48",x"a6",x"c8",x"87"),
   156 => (x"ec",x"c0",x"78",x"c1"),
   157 => (x"48",x"a6",x"d0",x"87"),
   158 => (x"80",x"f8",x"78",x"c1"),
   159 => (x"e0",x"c0",x"78",x"c1"),
   160 => (x"ab",x"f0",x"c0",x"87"),
   161 => (x"c0",x"87",x"da",x"06"),
   162 => (x"d4",x"03",x"ab",x"f9"),
   163 => (x"49",x"66",x"d4",x"87"),
   164 => (x"4a",x"73",x"91",x"ca"),
   165 => (x"d4",x"8a",x"f0",x"c0"),
   166 => (x"a1",x"72",x"48",x"a6"),
   167 => (x"c1",x"80",x"f4",x"78"),
   168 => (x"02",x"66",x"cc",x"78"),
   169 => (x"c4",x"87",x"ea",x"c1"),
   170 => (x"c4",x"49",x"75",x"85"),
   171 => (x"69",x"48",x"a6",x"89"),
   172 => (x"ab",x"e4",x"c1",x"78"),
   173 => (x"c4",x"87",x"d8",x"05"),
   174 => (x"b7",x"c0",x"48",x"66"),
   175 => (x"87",x"cf",x"03",x"a8"),
   176 => (x"c1",x"49",x"ed",x"c0"),
   177 => (x"66",x"c4",x"87",x"fb"),
   178 => (x"88",x"08",x"c0",x"48"),
   179 => (x"d0",x"58",x"a6",x"c8"),
   180 => (x"66",x"d8",x"1e",x"66"),
   181 => (x"66",x"f8",x"c0",x"1e"),
   182 => (x"66",x"f8",x"c0",x"1e"),
   183 => (x"1e",x"66",x"dc",x"1e"),
   184 => (x"f6",x"49",x"66",x"d8"),
   185 => (x"86",x"d4",x"87",x"d5"),
   186 => (x"a4",x"71",x"49",x"70"),
   187 => (x"87",x"e1",x"c0",x"4c"),
   188 => (x"05",x"ab",x"e5",x"c0"),
   189 => (x"a6",x"d0",x"87",x"cf"),
   190 => (x"c4",x"78",x"c0",x"48"),
   191 => (x"f4",x"78",x"c0",x"80"),
   192 => (x"cc",x"78",x"c1",x"80"),
   193 => (x"66",x"f0",x"c0",x"87"),
   194 => (x"c0",x"49",x"73",x"1e"),
   195 => (x"c4",x"0f",x"66",x"f0"),
   196 => (x"bf",x"97",x"6e",x"86"),
   197 => (x"c1",x"48",x"6e",x"4b"),
   198 => (x"58",x"a6",x"c4",x"80"),
   199 => (x"f9",x"05",x"9b",x"73"),
   200 => (x"48",x"74",x"87",x"ed"),
   201 => (x"4d",x"26",x"8e",x"e8"),
   202 => (x"4b",x"26",x"4c",x"26"),
   203 => (x"c0",x"1e",x"4f",x"26"),
   204 => (x"1e",x"c1",x"cd",x"1e"),
   205 => (x"d0",x"1e",x"a6",x"d0"),
   206 => (x"eb",x"f8",x"49",x"66"),
   207 => (x"26",x"8e",x"f4",x"87"),
   208 => (x"86",x"fc",x"1e",x"4f"),
   209 => (x"c0",x"ff",x"4a",x"71"),
   210 => (x"c4",x"48",x"69",x"49"),
   211 => (x"a6",x"c4",x"98",x"c0"),
   212 => (x"f4",x"02",x"6e",x"58"),
   213 => (x"48",x"79",x"72",x"87"),
   214 => (x"4f",x"26",x"8e",x"fc"),
   215 => (x"12",x"1e",x"72",x"1e"),
   216 => (x"c4",x"02",x"11",x"48"),
   217 => (x"f6",x"02",x"88",x"87"),
   218 => (x"26",x"4a",x"26",x"87"),
   219 => (x"1e",x"73",x"1e",x"4f"),
   220 => (x"c0",x"02",x"9a",x"72"),
   221 => (x"48",x"c0",x"87",x"e7"),
   222 => (x"a9",x"72",x"4b",x"c1"),
   223 => (x"72",x"87",x"d1",x"06"),
   224 => (x"87",x"c9",x"06",x"82"),
   225 => (x"a9",x"72",x"83",x"73"),
   226 => (x"c3",x"87",x"f4",x"01"),
   227 => (x"3a",x"b2",x"c1",x"87"),
   228 => (x"89",x"03",x"a9",x"72"),
   229 => (x"c1",x"07",x"80",x"73"),
   230 => (x"f3",x"05",x"2b",x"2a"),
   231 => (x"26",x"4b",x"26",x"87"),
   232 => (x"1e",x"75",x"1e",x"4f"),
   233 => (x"b7",x"71",x"4d",x"c4"),
   234 => (x"b9",x"ff",x"04",x"a1"),
   235 => (x"bd",x"c3",x"81",x"c1"),
   236 => (x"a2",x"b7",x"72",x"07"),
   237 => (x"c1",x"ba",x"ff",x"04"),
   238 => (x"07",x"bd",x"c1",x"82"),
   239 => (x"c1",x"87",x"ee",x"fe"),
   240 => (x"b8",x"ff",x"04",x"2d"),
   241 => (x"2d",x"07",x"80",x"c1"),
   242 => (x"c1",x"b9",x"ff",x"04"),
   243 => (x"4d",x"26",x"07",x"81"),
   244 => (x"5e",x"0e",x"4f",x"26"),
   245 => (x"0e",x"5d",x"5c",x"5b"),
   246 => (x"c1",x"86",x"dc",x"ff"),
   247 => (x"c3",x"48",x"e0",x"cf"),
   248 => (x"c1",x"78",x"e4",x"ef"),
   249 => (x"c3",x"48",x"dc",x"cf"),
   250 => (x"48",x"78",x"d4",x"f0"),
   251 => (x"78",x"e4",x"ef",x"c3"),
   252 => (x"48",x"d8",x"f0",x"c3"),
   253 => (x"80",x"c4",x"78",x"c0"),
   254 => (x"80",x"c4",x"78",x"c2"),
   255 => (x"71",x"78",x"e8",x"c0"),
   256 => (x"c8",x"ee",x"c0",x"1e"),
   257 => (x"e4",x"f0",x"c3",x"48"),
   258 => (x"20",x"41",x"20",x"49"),
   259 => (x"20",x"41",x"20",x"41"),
   260 => (x"20",x"41",x"20",x"41"),
   261 => (x"10",x"41",x"20",x"41"),
   262 => (x"10",x"51",x"10",x"51"),
   263 => (x"1e",x"49",x"26",x"51"),
   264 => (x"48",x"e8",x"ee",x"c0"),
   265 => (x"49",x"c4",x"f1",x"c3"),
   266 => (x"41",x"20",x"41",x"20"),
   267 => (x"41",x"20",x"41",x"20"),
   268 => (x"41",x"20",x"41",x"20"),
   269 => (x"51",x"10",x"41",x"20"),
   270 => (x"51",x"10",x"51",x"10"),
   271 => (x"ec",x"c1",x"49",x"26"),
   272 => (x"78",x"ca",x"48",x"d8"),
   273 => (x"1e",x"c8",x"ef",x"c0"),
   274 => (x"c0",x"87",x"e3",x"fb"),
   275 => (x"fb",x"1e",x"cc",x"ef"),
   276 => (x"ef",x"c0",x"87",x"dc"),
   277 => (x"d5",x"fb",x"1e",x"fc"),
   278 => (x"c0",x"86",x"cc",x"87"),
   279 => (x"02",x"bf",x"ec",x"e7"),
   280 => (x"e7",x"c0",x"87",x"d2"),
   281 => (x"c5",x"fb",x"1e",x"f4"),
   282 => (x"e0",x"e8",x"c0",x"87"),
   283 => (x"87",x"fe",x"fa",x"1e"),
   284 => (x"87",x"d0",x"86",x"c8"),
   285 => (x"1e",x"e4",x"e8",x"c0"),
   286 => (x"c0",x"87",x"f3",x"fa"),
   287 => (x"fa",x"1e",x"d4",x"e9"),
   288 => (x"86",x"c8",x"87",x"ec"),
   289 => (x"bf",x"f0",x"e7",x"c0"),
   290 => (x"c0",x"f0",x"c0",x"1e"),
   291 => (x"87",x"de",x"fa",x"1e"),
   292 => (x"ef",x"c3",x"86",x"c8"),
   293 => (x"c8",x"ff",x"48",x"cc"),
   294 => (x"a6",x"c4",x"78",x"bf"),
   295 => (x"c0",x"78",x"c1",x"48"),
   296 => (x"48",x"bf",x"f0",x"e7"),
   297 => (x"06",x"a8",x"b7",x"c0"),
   298 => (x"c8",x"87",x"eb",x"c8"),
   299 => (x"a6",x"d0",x"48",x"a6"),
   300 => (x"48",x"a6",x"d0",x"58"),
   301 => (x"d8",x"58",x"a6",x"d8"),
   302 => (x"a6",x"c4",x"48",x"a6"),
   303 => (x"ec",x"cf",x"c1",x"58"),
   304 => (x"50",x"c1",x"c1",x"48"),
   305 => (x"48",x"e8",x"cf",x"c1"),
   306 => (x"cf",x"c1",x"78",x"c0"),
   307 => (x"49",x"bf",x"97",x"ec"),
   308 => (x"02",x"a9",x"c1",x"c1"),
   309 => (x"dc",x"87",x"c8",x"c0"),
   310 => (x"78",x"c0",x"48",x"a6"),
   311 => (x"dc",x"87",x"c5",x"c0"),
   312 => (x"78",x"c1",x"48",x"a6"),
   313 => (x"bf",x"e8",x"cf",x"c1"),
   314 => (x"b0",x"66",x"dc",x"48"),
   315 => (x"58",x"ec",x"cf",x"c1"),
   316 => (x"48",x"f0",x"cf",x"c1"),
   317 => (x"d8",x"50",x"c2",x"c1"),
   318 => (x"78",x"c2",x"48",x"a6"),
   319 => (x"78",x"c3",x"80",x"c8"),
   320 => (x"48",x"f8",x"e9",x"c0"),
   321 => (x"49",x"e4",x"f1",x"c3"),
   322 => (x"41",x"20",x"41",x"20"),
   323 => (x"41",x"20",x"41",x"20"),
   324 => (x"41",x"20",x"41",x"20"),
   325 => (x"51",x"10",x"41",x"20"),
   326 => (x"51",x"10",x"51",x"10"),
   327 => (x"c1",x"48",x"a6",x"d0"),
   328 => (x"e4",x"f1",x"c3",x"78"),
   329 => (x"c4",x"f1",x"c3",x"1e"),
   330 => (x"e6",x"f8",x"c0",x"49"),
   331 => (x"70",x"86",x"c4",x"87"),
   332 => (x"c8",x"c0",x"05",x"98"),
   333 => (x"48",x"a6",x"dc",x"87"),
   334 => (x"c5",x"c0",x"78",x"c1"),
   335 => (x"48",x"a6",x"dc",x"87"),
   336 => (x"cf",x"c1",x"78",x"c0"),
   337 => (x"66",x"dc",x"48",x"e8"),
   338 => (x"48",x"66",x"d8",x"78"),
   339 => (x"03",x"a8",x"b7",x"c3"),
   340 => (x"d8",x"87",x"ea",x"c0"),
   341 => (x"91",x"c5",x"49",x"66"),
   342 => (x"88",x"c3",x"48",x"71"),
   343 => (x"cc",x"58",x"a6",x"cc"),
   344 => (x"1e",x"c3",x"1e",x"66"),
   345 => (x"49",x"66",x"e0",x"c0"),
   346 => (x"87",x"f0",x"f4",x"c0"),
   347 => (x"66",x"d8",x"86",x"c8"),
   348 => (x"dc",x"80",x"c1",x"48"),
   349 => (x"b7",x"c3",x"58",x"a6"),
   350 => (x"d6",x"ff",x"04",x"a8"),
   351 => (x"1e",x"66",x"c8",x"87"),
   352 => (x"c1",x"1e",x"66",x"dc"),
   353 => (x"c1",x"1e",x"fc",x"d2"),
   354 => (x"c0",x"49",x"f4",x"cf"),
   355 => (x"cc",x"87",x"df",x"f4"),
   356 => (x"dc",x"cf",x"c1",x"86"),
   357 => (x"cf",x"c1",x"4c",x"bf"),
   358 => (x"4b",x"bf",x"bf",x"dc"),
   359 => (x"cf",x"c1",x"1e",x"72"),
   360 => (x"73",x"48",x"bf",x"dc"),
   361 => (x"a1",x"f0",x"c0",x"49"),
   362 => (x"71",x"41",x"20",x"4a"),
   363 => (x"f8",x"ff",x"05",x"aa"),
   364 => (x"cc",x"4a",x"26",x"87"),
   365 => (x"79",x"c5",x"49",x"a4"),
   366 => (x"69",x"4d",x"a3",x"cc"),
   367 => (x"73",x"7b",x"6c",x"7d"),
   368 => (x"87",x"c0",x"d0",x"49"),
   369 => (x"69",x"49",x"a3",x"c4"),
   370 => (x"87",x"e5",x"c0",x"05"),
   371 => (x"c6",x"49",x"a3",x"c8"),
   372 => (x"c8",x"1e",x"71",x"7d"),
   373 => (x"49",x"6a",x"4a",x"a4"),
   374 => (x"87",x"e3",x"f1",x"c0"),
   375 => (x"bf",x"dc",x"cf",x"c1"),
   376 => (x"1e",x"75",x"7b",x"bf"),
   377 => (x"49",x"6d",x"1e",x"ca"),
   378 => (x"87",x"f0",x"f2",x"c0"),
   379 => (x"d9",x"c0",x"86",x"cc"),
   380 => (x"1e",x"49",x"6c",x"87"),
   381 => (x"48",x"71",x"1e",x"72"),
   382 => (x"f0",x"c0",x"49",x"74"),
   383 => (x"41",x"20",x"4a",x"a1"),
   384 => (x"ff",x"05",x"aa",x"71"),
   385 => (x"4a",x"26",x"87",x"f8"),
   386 => (x"a6",x"dc",x"49",x"26"),
   387 => (x"50",x"c1",x"c1",x"48"),
   388 => (x"97",x"f0",x"cf",x"c1"),
   389 => (x"c1",x"c1",x"49",x"bf"),
   390 => (x"c1",x"04",x"a9",x"b7"),
   391 => (x"97",x"dc",x"87",x"db"),
   392 => (x"c3",x"c1",x"4b",x"66"),
   393 => (x"c0",x"49",x"73",x"1e"),
   394 => (x"c4",x"87",x"c6",x"f4"),
   395 => (x"a8",x"66",x"d0",x"86"),
   396 => (x"87",x"f5",x"c0",x"05"),
   397 => (x"c0",x"1e",x"66",x"d4"),
   398 => (x"c2",x"f0",x"c0",x"49"),
   399 => (x"c0",x"86",x"c4",x"87"),
   400 => (x"c3",x"48",x"d8",x"e9"),
   401 => (x"20",x"49",x"e4",x"f1"),
   402 => (x"20",x"41",x"20",x"41"),
   403 => (x"20",x"41",x"20",x"41"),
   404 => (x"20",x"41",x"20",x"41"),
   405 => (x"10",x"51",x"10",x"41"),
   406 => (x"c0",x"51",x"10",x"51"),
   407 => (x"c4",x"48",x"a6",x"e0"),
   408 => (x"cf",x"c1",x"78",x"66"),
   409 => (x"66",x"c4",x"48",x"e4"),
   410 => (x"73",x"83",x"c1",x"78"),
   411 => (x"f0",x"cf",x"c1",x"4a"),
   412 => (x"b7",x"49",x"bf",x"97"),
   413 => (x"e9",x"fe",x"06",x"aa"),
   414 => (x"66",x"e0",x"c0",x"87"),
   415 => (x"90",x"66",x"d8",x"48"),
   416 => (x"58",x"a6",x"e4",x"c0"),
   417 => (x"49",x"70",x"1e",x"72"),
   418 => (x"f4",x"4a",x"66",x"cc"),
   419 => (x"4a",x"26",x"87",x"d3"),
   420 => (x"c0",x"58",x"a6",x"dc"),
   421 => (x"c8",x"49",x"66",x"e0"),
   422 => (x"91",x"c7",x"89",x"66"),
   423 => (x"66",x"d8",x"48",x"71"),
   424 => (x"a6",x"e4",x"c0",x"88"),
   425 => (x"4a",x"bf",x"6e",x"58"),
   426 => (x"cf",x"c1",x"82",x"ca"),
   427 => (x"49",x"bf",x"97",x"ec"),
   428 => (x"05",x"a9",x"c1",x"c1"),
   429 => (x"c1",x"87",x"cd",x"c0"),
   430 => (x"c1",x"48",x"72",x"8a"),
   431 => (x"88",x"bf",x"e4",x"cf"),
   432 => (x"08",x"78",x"08",x"6e"),
   433 => (x"c1",x"48",x"66",x"c4"),
   434 => (x"58",x"a6",x"c8",x"80"),
   435 => (x"bf",x"f0",x"e7",x"c0"),
   436 => (x"f7",x"06",x"a8",x"b7"),
   437 => (x"ef",x"c3",x"87",x"e7"),
   438 => (x"c8",x"ff",x"48",x"d0"),
   439 => (x"f0",x"c0",x"78",x"bf"),
   440 => (x"c9",x"f1",x"1e",x"f0"),
   441 => (x"c0",x"f1",x"c0",x"87"),
   442 => (x"87",x"c2",x"f1",x"1e"),
   443 => (x"1e",x"c4",x"f1",x"c0"),
   444 => (x"c0",x"87",x"fb",x"f0"),
   445 => (x"f0",x"1e",x"fc",x"f1"),
   446 => (x"cf",x"c1",x"87",x"f4"),
   447 => (x"c0",x"1e",x"bf",x"e4"),
   448 => (x"f0",x"1e",x"c0",x"f2"),
   449 => (x"1e",x"c5",x"87",x"e8"),
   450 => (x"1e",x"dc",x"f2",x"c0"),
   451 => (x"c1",x"87",x"df",x"f0"),
   452 => (x"1e",x"bf",x"e8",x"cf"),
   453 => (x"1e",x"f8",x"f2",x"c0"),
   454 => (x"c1",x"87",x"d3",x"f0"),
   455 => (x"d4",x"f3",x"c0",x"1e"),
   456 => (x"87",x"ca",x"f0",x"1e"),
   457 => (x"97",x"ec",x"cf",x"c1"),
   458 => (x"c0",x"1e",x"49",x"bf"),
   459 => (x"ef",x"1e",x"f0",x"f3"),
   460 => (x"c1",x"c1",x"87",x"fc"),
   461 => (x"cc",x"f4",x"c0",x"1e"),
   462 => (x"87",x"f2",x"ef",x"1e"),
   463 => (x"97",x"f0",x"cf",x"c1"),
   464 => (x"c0",x"1e",x"49",x"bf"),
   465 => (x"ef",x"1e",x"e8",x"f4"),
   466 => (x"c2",x"c1",x"87",x"e4"),
   467 => (x"c4",x"f5",x"c0",x"1e"),
   468 => (x"87",x"da",x"ef",x"1e"),
   469 => (x"bf",x"d4",x"d0",x"c1"),
   470 => (x"e0",x"f5",x"c0",x"1e"),
   471 => (x"87",x"ce",x"ef",x"1e"),
   472 => (x"f5",x"c0",x"1e",x"c7"),
   473 => (x"c5",x"ef",x"1e",x"fc"),
   474 => (x"d8",x"ec",x"c1",x"87"),
   475 => (x"f6",x"c0",x"1e",x"bf"),
   476 => (x"f9",x"ee",x"1e",x"d8"),
   477 => (x"f4",x"f6",x"c0",x"87"),
   478 => (x"87",x"f2",x"ee",x"1e"),
   479 => (x"1e",x"e0",x"f7",x"c0"),
   480 => (x"c1",x"87",x"eb",x"ee"),
   481 => (x"bf",x"bf",x"dc",x"cf"),
   482 => (x"ec",x"f7",x"c0",x"1e"),
   483 => (x"87",x"de",x"ee",x"1e"),
   484 => (x"1e",x"c8",x"f8",x"c0"),
   485 => (x"c1",x"87",x"d7",x"ee"),
   486 => (x"49",x"bf",x"dc",x"cf"),
   487 => (x"1e",x"69",x"81",x"c4"),
   488 => (x"1e",x"fc",x"f8",x"c0"),
   489 => (x"c0",x"87",x"c7",x"ee"),
   490 => (x"d8",x"f9",x"c0",x"1e"),
   491 => (x"87",x"fe",x"ed",x"1e"),
   492 => (x"bf",x"dc",x"cf",x"c1"),
   493 => (x"69",x"81",x"c8",x"49"),
   494 => (x"f4",x"f9",x"c0",x"1e"),
   495 => (x"87",x"ee",x"ed",x"1e"),
   496 => (x"fa",x"c0",x"1e",x"c2"),
   497 => (x"e5",x"ed",x"1e",x"d0"),
   498 => (x"dc",x"cf",x"c1",x"87"),
   499 => (x"81",x"cc",x"49",x"bf"),
   500 => (x"fa",x"c0",x"1e",x"69"),
   501 => (x"d5",x"ed",x"1e",x"ec"),
   502 => (x"c0",x"1e",x"d1",x"87"),
   503 => (x"ed",x"1e",x"c8",x"fb"),
   504 => (x"cf",x"c1",x"87",x"cc"),
   505 => (x"d0",x"49",x"bf",x"dc"),
   506 => (x"c0",x"1e",x"71",x"81"),
   507 => (x"ec",x"1e",x"e4",x"fb"),
   508 => (x"fc",x"c0",x"87",x"fc"),
   509 => (x"f5",x"ec",x"1e",x"c0"),
   510 => (x"f8",x"fc",x"c0",x"87"),
   511 => (x"87",x"ee",x"ec",x"1e"),
   512 => (x"bf",x"e0",x"cf",x"c1"),
   513 => (x"fd",x"c0",x"1e",x"bf"),
   514 => (x"e1",x"ec",x"1e",x"cc"),
   515 => (x"e8",x"fd",x"c0",x"87"),
   516 => (x"87",x"da",x"ec",x"1e"),
   517 => (x"bf",x"e0",x"cf",x"c1"),
   518 => (x"69",x"81",x"c4",x"49"),
   519 => (x"e8",x"fe",x"c0",x"1e"),
   520 => (x"87",x"ca",x"ec",x"1e"),
   521 => (x"ff",x"c0",x"1e",x"c0"),
   522 => (x"c1",x"ec",x"1e",x"c4"),
   523 => (x"e0",x"cf",x"c1",x"87"),
   524 => (x"81",x"c8",x"49",x"bf"),
   525 => (x"ff",x"c0",x"1e",x"69"),
   526 => (x"f1",x"eb",x"1e",x"e0"),
   527 => (x"c0",x"1e",x"c1",x"87"),
   528 => (x"eb",x"1e",x"fc",x"ff"),
   529 => (x"cf",x"c1",x"87",x"e8"),
   530 => (x"cc",x"49",x"bf",x"e0"),
   531 => (x"c1",x"1e",x"69",x"81"),
   532 => (x"eb",x"1e",x"d8",x"c0"),
   533 => (x"1e",x"d2",x"87",x"d8"),
   534 => (x"1e",x"f4",x"c0",x"c1"),
   535 => (x"c1",x"87",x"cf",x"eb"),
   536 => (x"49",x"bf",x"e0",x"cf"),
   537 => (x"1e",x"71",x"81",x"d0"),
   538 => (x"1e",x"d0",x"c1",x"c1"),
   539 => (x"c1",x"87",x"ff",x"ea"),
   540 => (x"ea",x"1e",x"ec",x"c1"),
   541 => (x"dc",x"c4",x"87",x"f8"),
   542 => (x"c2",x"c1",x"1e",x"66"),
   543 => (x"ed",x"ea",x"1e",x"e4"),
   544 => (x"c1",x"1e",x"c5",x"87"),
   545 => (x"ea",x"1e",x"c0",x"c3"),
   546 => (x"f4",x"c4",x"87",x"e4"),
   547 => (x"c3",x"c1",x"1e",x"66"),
   548 => (x"d9",x"ea",x"1e",x"dc"),
   549 => (x"c1",x"1e",x"cd",x"87"),
   550 => (x"ea",x"1e",x"f8",x"c3"),
   551 => (x"ec",x"c4",x"87",x"d0"),
   552 => (x"c4",x"c1",x"1e",x"66"),
   553 => (x"c5",x"ea",x"1e",x"d4"),
   554 => (x"c1",x"1e",x"c7",x"87"),
   555 => (x"e9",x"1e",x"f0",x"c4"),
   556 => (x"c4",x"c5",x"87",x"fc"),
   557 => (x"c5",x"c1",x"1e",x"66"),
   558 => (x"f1",x"e9",x"1e",x"cc"),
   559 => (x"c1",x"1e",x"c1",x"87"),
   560 => (x"e9",x"1e",x"e8",x"c5"),
   561 => (x"f1",x"c3",x"87",x"e8"),
   562 => (x"c6",x"c1",x"1e",x"c4"),
   563 => (x"dd",x"e9",x"1e",x"c4"),
   564 => (x"e0",x"c6",x"c1",x"87"),
   565 => (x"87",x"d6",x"e9",x"1e"),
   566 => (x"1e",x"e4",x"f1",x"c3"),
   567 => (x"1e",x"d8",x"c7",x"c1"),
   568 => (x"c1",x"87",x"cb",x"e9"),
   569 => (x"e9",x"1e",x"f4",x"c7"),
   570 => (x"c8",x"c1",x"87",x"c4"),
   571 => (x"fd",x"e8",x"1e",x"ec"),
   572 => (x"d0",x"ef",x"c3",x"87"),
   573 => (x"ef",x"c3",x"49",x"bf"),
   574 => (x"c3",x"89",x"bf",x"cc"),
   575 => (x"71",x"59",x"d8",x"ef"),
   576 => (x"f0",x"c8",x"c1",x"1e"),
   577 => (x"87",x"e6",x"e8",x"1e"),
   578 => (x"c3",x"86",x"e8",x"c5"),
   579 => (x"48",x"bf",x"d4",x"ef"),
   580 => (x"a8",x"b7",x"f8",x"c1"),
   581 => (x"87",x"d7",x"c0",x"03"),
   582 => (x"1e",x"d8",x"ea",x"c0"),
   583 => (x"c0",x"87",x"cf",x"e8"),
   584 => (x"e8",x"1e",x"d0",x"eb"),
   585 => (x"eb",x"c0",x"87",x"c8"),
   586 => (x"c1",x"e8",x"1e",x"f0"),
   587 => (x"c3",x"86",x"cc",x"87"),
   588 => (x"49",x"bf",x"d4",x"ef"),
   589 => (x"92",x"e8",x"cf",x"4a"),
   590 => (x"1e",x"72",x"1e",x"71"),
   591 => (x"e7",x"c0",x"49",x"72"),
   592 => (x"e9",x"4a",x"bf",x"f0"),
   593 => (x"4a",x"26",x"87",x"db"),
   594 => (x"ef",x"c3",x"49",x"26"),
   595 => (x"e7",x"c0",x"58",x"dc"),
   596 => (x"4b",x"4a",x"bf",x"f0"),
   597 => (x"71",x"93",x"e8",x"cf"),
   598 => (x"73",x"1e",x"72",x"1e"),
   599 => (x"c0",x"e9",x"4a",x"09"),
   600 => (x"26",x"4a",x"26",x"87"),
   601 => (x"e0",x"ef",x"c3",x"49"),
   602 => (x"92",x"f9",x"c8",x"58"),
   603 => (x"1e",x"72",x"1e",x"71"),
   604 => (x"e8",x"4a",x"09",x"72"),
   605 => (x"4a",x"26",x"87",x"eb"),
   606 => (x"ef",x"c3",x"49",x"26"),
   607 => (x"eb",x"c0",x"58",x"e4"),
   608 => (x"e9",x"e6",x"1e",x"f4"),
   609 => (x"d8",x"ef",x"c3",x"87"),
   610 => (x"ec",x"c0",x"1e",x"bf"),
   611 => (x"dd",x"e6",x"1e",x"e4"),
   612 => (x"ec",x"ec",x"c0",x"87"),
   613 => (x"87",x"d6",x"e6",x"1e"),
   614 => (x"bf",x"dc",x"ef",x"c3"),
   615 => (x"dc",x"ed",x"c0",x"1e"),
   616 => (x"87",x"ca",x"e6",x"1e"),
   617 => (x"bf",x"e0",x"ef",x"c3"),
   618 => (x"e4",x"ed",x"c0",x"1e"),
   619 => (x"87",x"fe",x"e5",x"1e"),
   620 => (x"1e",x"c4",x"ee",x"c0"),
   621 => (x"c0",x"87",x"f7",x"e5"),
   622 => (x"8e",x"f8",x"fe",x"48"),
   623 => (x"4c",x"26",x"4d",x"26"),
   624 => (x"4f",x"26",x"4b",x"26"),
   625 => (x"c1",x"4a",x"71",x"1e"),
   626 => (x"02",x"bf",x"dc",x"cf"),
   627 => (x"cf",x"c1",x"87",x"c6"),
   628 => (x"7a",x"bf",x"bf",x"dc"),
   629 => (x"bf",x"dc",x"cf",x"c1"),
   630 => (x"71",x"81",x"cc",x"49"),
   631 => (x"e4",x"cf",x"c1",x"1e"),
   632 => (x"49",x"ca",x"1e",x"bf"),
   633 => (x"87",x"f4",x"e2",x"c0"),
   634 => (x"4f",x"26",x"8e",x"f8"),
   635 => (x"00",x"00",x"00",x"00"),
   636 => (x"00",x"00",x"61",x"a8"),
   637 => (x"67",x"6f",x"72",x"50"),
   638 => (x"20",x"6d",x"61",x"72"),
   639 => (x"70",x"6d",x"6f",x"63"),
   640 => (x"64",x"65",x"6c",x"69"),
   641 => (x"74",x"69",x"77",x"20"),
   642 => (x"72",x"27",x"20",x"68"),
   643 => (x"73",x"69",x"67",x"65"),
   644 => (x"27",x"72",x"65",x"74"),
   645 => (x"74",x"74",x"61",x"20"),
   646 => (x"75",x"62",x"69",x"72"),
   647 => (x"00",x"0a",x"65",x"74"),
   648 => (x"00",x"00",x"00",x"0a"),
   649 => (x"67",x"6f",x"72",x"50"),
   650 => (x"20",x"6d",x"61",x"72"),
   651 => (x"70",x"6d",x"6f",x"63"),
   652 => (x"64",x"65",x"6c",x"69"),
   653 => (x"74",x"69",x"77",x"20"),
   654 => (x"74",x"75",x"6f",x"68"),
   655 => (x"65",x"72",x"27",x"20"),
   656 => (x"74",x"73",x"69",x"67"),
   657 => (x"20",x"27",x"72",x"65"),
   658 => (x"72",x"74",x"74",x"61"),
   659 => (x"74",x"75",x"62",x"69"),
   660 => (x"00",x"00",x"0a",x"65"),
   661 => (x"00",x"00",x"00",x"0a"),
   662 => (x"59",x"52",x"48",x"44"),
   663 => (x"4e",x"4f",x"54",x"53"),
   664 => (x"52",x"50",x"20",x"45"),
   665 => (x"41",x"52",x"47",x"4f"),
   666 => (x"33",x"20",x"2c",x"4d"),
   667 => (x"20",x"44",x"52",x"27"),
   668 => (x"49",x"52",x"54",x"53"),
   669 => (x"00",x"00",x"47",x"4e"),
   670 => (x"59",x"52",x"48",x"44"),
   671 => (x"4e",x"4f",x"54",x"53"),
   672 => (x"52",x"50",x"20",x"45"),
   673 => (x"41",x"52",x"47",x"4f"),
   674 => (x"32",x"20",x"2c",x"4d"),
   675 => (x"20",x"44",x"4e",x"27"),
   676 => (x"49",x"52",x"54",x"53"),
   677 => (x"00",x"00",x"47",x"4e"),
   678 => (x"73",x"61",x"65",x"4d"),
   679 => (x"64",x"65",x"72",x"75"),
   680 => (x"6d",x"69",x"74",x"20"),
   681 => (x"6f",x"74",x"20",x"65"),
   682 => (x"6d",x"73",x"20",x"6f"),
   683 => (x"20",x"6c",x"6c",x"61"),
   684 => (x"6f",x"20",x"6f",x"74"),
   685 => (x"69",x"61",x"74",x"62"),
   686 => (x"65",x"6d",x"20",x"6e"),
   687 => (x"6e",x"69",x"6e",x"61"),
   688 => (x"6c",x"75",x"66",x"67"),
   689 => (x"73",x"65",x"72",x"20"),
   690 => (x"73",x"74",x"6c",x"75"),
   691 => (x"00",x"00",x"00",x"0a"),
   692 => (x"61",x"65",x"6c",x"50"),
   693 => (x"69",x"20",x"65",x"73"),
   694 => (x"65",x"72",x"63",x"6e"),
   695 => (x"20",x"65",x"73",x"61"),
   696 => (x"62",x"6d",x"75",x"6e"),
   697 => (x"6f",x"20",x"72",x"65"),
   698 => (x"75",x"72",x"20",x"66"),
   699 => (x"00",x"0a",x"73",x"6e"),
   700 => (x"00",x"00",x"00",x"0a"),
   701 => (x"72",x"63",x"69",x"4d"),
   702 => (x"63",x"65",x"73",x"6f"),
   703 => (x"73",x"64",x"6e",x"6f"),
   704 => (x"72",x"6f",x"66",x"20"),
   705 => (x"65",x"6e",x"6f",x"20"),
   706 => (x"6e",x"75",x"72",x"20"),
   707 => (x"72",x"68",x"74",x"20"),
   708 => (x"68",x"67",x"75",x"6f"),
   709 => (x"72",x"68",x"44",x"20"),
   710 => (x"6f",x"74",x"73",x"79"),
   711 => (x"20",x"3a",x"65",x"6e"),
   712 => (x"00",x"00",x"00",x"00"),
   713 => (x"0a",x"20",x"64",x"25"),
   714 => (x"00",x"00",x"00",x"00"),
   715 => (x"79",x"72",x"68",x"44"),
   716 => (x"6e",x"6f",x"74",x"73"),
   717 => (x"70",x"20",x"73",x"65"),
   718 => (x"53",x"20",x"72",x"65"),
   719 => (x"6e",x"6f",x"63",x"65"),
   720 => (x"20",x"20",x"3a",x"64"),
   721 => (x"20",x"20",x"20",x"20"),
   722 => (x"20",x"20",x"20",x"20"),
   723 => (x"20",x"20",x"20",x"20"),
   724 => (x"20",x"20",x"20",x"20"),
   725 => (x"20",x"20",x"20",x"20"),
   726 => (x"00",x"00",x"00",x"00"),
   727 => (x"0a",x"20",x"64",x"25"),
   728 => (x"00",x"00",x"00",x"00"),
   729 => (x"20",x"58",x"41",x"56"),
   730 => (x"53",x"50",x"49",x"4d"),
   731 => (x"74",x"61",x"72",x"20"),
   732 => (x"20",x"67",x"6e",x"69"),
   733 => (x"30",x"31",x"20",x"2a"),
   734 => (x"3d",x"20",x"30",x"30"),
   735 => (x"20",x"64",x"25",x"20"),
   736 => (x"00",x"00",x"00",x"0a"),
   737 => (x"00",x"00",x"00",x"0a"),
   738 => (x"59",x"52",x"48",x"44"),
   739 => (x"4e",x"4f",x"54",x"53"),
   740 => (x"52",x"50",x"20",x"45"),
   741 => (x"41",x"52",x"47",x"4f"),
   742 => (x"53",x"20",x"2c",x"4d"),
   743 => (x"20",x"45",x"4d",x"4f"),
   744 => (x"49",x"52",x"54",x"53"),
   745 => (x"00",x"00",x"47",x"4e"),
   746 => (x"59",x"52",x"48",x"44"),
   747 => (x"4e",x"4f",x"54",x"53"),
   748 => (x"52",x"50",x"20",x"45"),
   749 => (x"41",x"52",x"47",x"4f"),
   750 => (x"31",x"20",x"2c",x"4d"),
   751 => (x"20",x"54",x"53",x"27"),
   752 => (x"49",x"52",x"54",x"53"),
   753 => (x"00",x"00",x"47",x"4e"),
   754 => (x"00",x"00",x"00",x"0a"),
   755 => (x"79",x"72",x"68",x"44"),
   756 => (x"6e",x"6f",x"74",x"73"),
   757 => (x"65",x"42",x"20",x"65"),
   758 => (x"6d",x"68",x"63",x"6e"),
   759 => (x"2c",x"6b",x"72",x"61"),
   760 => (x"72",x"65",x"56",x"20"),
   761 => (x"6e",x"6f",x"69",x"73"),
   762 => (x"31",x"2e",x"32",x"20"),
   763 => (x"61",x"4c",x"28",x"20"),
   764 => (x"61",x"75",x"67",x"6e"),
   765 => (x"20",x"3a",x"65",x"67"),
   766 => (x"00",x"0a",x"29",x"43"),
   767 => (x"00",x"00",x"00",x"0a"),
   768 => (x"63",x"65",x"78",x"45"),
   769 => (x"6f",x"69",x"74",x"75"),
   770 => (x"74",x"73",x"20",x"6e"),
   771 => (x"73",x"74",x"72",x"61"),
   772 => (x"64",x"25",x"20",x"2c"),
   773 => (x"6e",x"75",x"72",x"20"),
   774 => (x"68",x"74",x"20",x"73"),
   775 => (x"67",x"75",x"6f",x"72"),
   776 => (x"68",x"44",x"20",x"68"),
   777 => (x"74",x"73",x"79",x"72"),
   778 => (x"0a",x"65",x"6e",x"6f"),
   779 => (x"00",x"00",x"00",x"00"),
   780 => (x"63",x"65",x"78",x"45"),
   781 => (x"6f",x"69",x"74",x"75"),
   782 => (x"6e",x"65",x"20",x"6e"),
   783 => (x"00",x"0a",x"73",x"64"),
   784 => (x"00",x"00",x"00",x"0a"),
   785 => (x"61",x"6e",x"69",x"46"),
   786 => (x"61",x"76",x"20",x"6c"),
   787 => (x"73",x"65",x"75",x"6c"),
   788 => (x"20",x"66",x"6f",x"20"),
   789 => (x"20",x"65",x"68",x"74"),
   790 => (x"69",x"72",x"61",x"76"),
   791 => (x"65",x"6c",x"62",x"61"),
   792 => (x"73",x"75",x"20",x"73"),
   793 => (x"69",x"20",x"64",x"65"),
   794 => (x"68",x"74",x"20",x"6e"),
   795 => (x"65",x"62",x"20",x"65"),
   796 => (x"6d",x"68",x"63",x"6e"),
   797 => (x"3a",x"6b",x"72",x"61"),
   798 => (x"00",x"00",x"00",x"0a"),
   799 => (x"00",x"00",x"00",x"0a"),
   800 => (x"5f",x"74",x"6e",x"49"),
   801 => (x"62",x"6f",x"6c",x"47"),
   802 => (x"20",x"20",x"20",x"3a"),
   803 => (x"20",x"20",x"20",x"20"),
   804 => (x"20",x"20",x"20",x"20"),
   805 => (x"0a",x"64",x"25",x"20"),
   806 => (x"00",x"00",x"00",x"00"),
   807 => (x"20",x"20",x"20",x"20"),
   808 => (x"20",x"20",x"20",x"20"),
   809 => (x"75",x"6f",x"68",x"73"),
   810 => (x"62",x"20",x"64",x"6c"),
   811 => (x"20",x"20",x"3a",x"65"),
   812 => (x"0a",x"64",x"25",x"20"),
   813 => (x"00",x"00",x"00",x"00"),
   814 => (x"6c",x"6f",x"6f",x"42"),
   815 => (x"6f",x"6c",x"47",x"5f"),
   816 => (x"20",x"20",x"3a",x"62"),
   817 => (x"20",x"20",x"20",x"20"),
   818 => (x"20",x"20",x"20",x"20"),
   819 => (x"0a",x"64",x"25",x"20"),
   820 => (x"00",x"00",x"00",x"00"),
   821 => (x"20",x"20",x"20",x"20"),
   822 => (x"20",x"20",x"20",x"20"),
   823 => (x"75",x"6f",x"68",x"73"),
   824 => (x"62",x"20",x"64",x"6c"),
   825 => (x"20",x"20",x"3a",x"65"),
   826 => (x"0a",x"64",x"25",x"20"),
   827 => (x"00",x"00",x"00",x"00"),
   828 => (x"31",x"5f",x"68",x"43"),
   829 => (x"6f",x"6c",x"47",x"5f"),
   830 => (x"20",x"20",x"3a",x"62"),
   831 => (x"20",x"20",x"20",x"20"),
   832 => (x"20",x"20",x"20",x"20"),
   833 => (x"0a",x"63",x"25",x"20"),
   834 => (x"00",x"00",x"00",x"00"),
   835 => (x"20",x"20",x"20",x"20"),
   836 => (x"20",x"20",x"20",x"20"),
   837 => (x"75",x"6f",x"68",x"73"),
   838 => (x"62",x"20",x"64",x"6c"),
   839 => (x"20",x"20",x"3a",x"65"),
   840 => (x"0a",x"63",x"25",x"20"),
   841 => (x"00",x"00",x"00",x"00"),
   842 => (x"32",x"5f",x"68",x"43"),
   843 => (x"6f",x"6c",x"47",x"5f"),
   844 => (x"20",x"20",x"3a",x"62"),
   845 => (x"20",x"20",x"20",x"20"),
   846 => (x"20",x"20",x"20",x"20"),
   847 => (x"0a",x"63",x"25",x"20"),
   848 => (x"00",x"00",x"00",x"00"),
   849 => (x"20",x"20",x"20",x"20"),
   850 => (x"20",x"20",x"20",x"20"),
   851 => (x"75",x"6f",x"68",x"73"),
   852 => (x"62",x"20",x"64",x"6c"),
   853 => (x"20",x"20",x"3a",x"65"),
   854 => (x"0a",x"63",x"25",x"20"),
   855 => (x"00",x"00",x"00",x"00"),
   856 => (x"5f",x"72",x"72",x"41"),
   857 => (x"6c",x"47",x"5f",x"31"),
   858 => (x"38",x"5b",x"62",x"6f"),
   859 => (x"20",x"20",x"3a",x"5d"),
   860 => (x"20",x"20",x"20",x"20"),
   861 => (x"0a",x"64",x"25",x"20"),
   862 => (x"00",x"00",x"00",x"00"),
   863 => (x"20",x"20",x"20",x"20"),
   864 => (x"20",x"20",x"20",x"20"),
   865 => (x"75",x"6f",x"68",x"73"),
   866 => (x"62",x"20",x"64",x"6c"),
   867 => (x"20",x"20",x"3a",x"65"),
   868 => (x"0a",x"64",x"25",x"20"),
   869 => (x"00",x"00",x"00",x"00"),
   870 => (x"5f",x"72",x"72",x"41"),
   871 => (x"6c",x"47",x"5f",x"32"),
   872 => (x"38",x"5b",x"62",x"6f"),
   873 => (x"5d",x"37",x"5b",x"5d"),
   874 => (x"20",x"20",x"20",x"3a"),
   875 => (x"0a",x"64",x"25",x"20"),
   876 => (x"00",x"00",x"00",x"00"),
   877 => (x"20",x"20",x"20",x"20"),
   878 => (x"20",x"20",x"20",x"20"),
   879 => (x"75",x"6f",x"68",x"73"),
   880 => (x"62",x"20",x"64",x"6c"),
   881 => (x"20",x"20",x"3a",x"65"),
   882 => (x"6d",x"75",x"4e",x"20"),
   883 => (x"5f",x"72",x"65",x"62"),
   884 => (x"52",x"5f",x"66",x"4f"),
   885 => (x"20",x"73",x"6e",x"75"),
   886 => (x"30",x"31",x"20",x"2b"),
   887 => (x"00",x"00",x"00",x"0a"),
   888 => (x"5f",x"72",x"74",x"50"),
   889 => (x"62",x"6f",x"6c",x"47"),
   890 => (x"00",x"0a",x"3e",x"2d"),
   891 => (x"74",x"50",x"20",x"20"),
   892 => (x"6f",x"43",x"5f",x"72"),
   893 => (x"20",x"3a",x"70",x"6d"),
   894 => (x"20",x"20",x"20",x"20"),
   895 => (x"20",x"20",x"20",x"20"),
   896 => (x"0a",x"64",x"25",x"20"),
   897 => (x"00",x"00",x"00",x"00"),
   898 => (x"20",x"20",x"20",x"20"),
   899 => (x"20",x"20",x"20",x"20"),
   900 => (x"75",x"6f",x"68",x"73"),
   901 => (x"62",x"20",x"64",x"6c"),
   902 => (x"20",x"20",x"3a",x"65"),
   903 => (x"6d",x"69",x"28",x"20"),
   904 => (x"6d",x"65",x"6c",x"70"),
   905 => (x"61",x"74",x"6e",x"65"),
   906 => (x"6e",x"6f",x"69",x"74"),
   907 => (x"70",x"65",x"64",x"2d"),
   908 => (x"65",x"64",x"6e",x"65"),
   909 => (x"0a",x"29",x"74",x"6e"),
   910 => (x"00",x"00",x"00",x"00"),
   911 => (x"69",x"44",x"20",x"20"),
   912 => (x"3a",x"72",x"63",x"73"),
   913 => (x"20",x"20",x"20",x"20"),
   914 => (x"20",x"20",x"20",x"20"),
   915 => (x"20",x"20",x"20",x"20"),
   916 => (x"0a",x"64",x"25",x"20"),
   917 => (x"00",x"00",x"00",x"00"),
   918 => (x"20",x"20",x"20",x"20"),
   919 => (x"20",x"20",x"20",x"20"),
   920 => (x"75",x"6f",x"68",x"73"),
   921 => (x"62",x"20",x"64",x"6c"),
   922 => (x"20",x"20",x"3a",x"65"),
   923 => (x"0a",x"64",x"25",x"20"),
   924 => (x"00",x"00",x"00",x"00"),
   925 => (x"6e",x"45",x"20",x"20"),
   926 => (x"43",x"5f",x"6d",x"75"),
   927 => (x"3a",x"70",x"6d",x"6f"),
   928 => (x"20",x"20",x"20",x"20"),
   929 => (x"20",x"20",x"20",x"20"),
   930 => (x"0a",x"64",x"25",x"20"),
   931 => (x"00",x"00",x"00",x"00"),
   932 => (x"20",x"20",x"20",x"20"),
   933 => (x"20",x"20",x"20",x"20"),
   934 => (x"75",x"6f",x"68",x"73"),
   935 => (x"62",x"20",x"64",x"6c"),
   936 => (x"20",x"20",x"3a",x"65"),
   937 => (x"0a",x"64",x"25",x"20"),
   938 => (x"00",x"00",x"00",x"00"),
   939 => (x"6e",x"49",x"20",x"20"),
   940 => (x"6f",x"43",x"5f",x"74"),
   941 => (x"20",x"3a",x"70",x"6d"),
   942 => (x"20",x"20",x"20",x"20"),
   943 => (x"20",x"20",x"20",x"20"),
   944 => (x"0a",x"64",x"25",x"20"),
   945 => (x"00",x"00",x"00",x"00"),
   946 => (x"20",x"20",x"20",x"20"),
   947 => (x"20",x"20",x"20",x"20"),
   948 => (x"75",x"6f",x"68",x"73"),
   949 => (x"62",x"20",x"64",x"6c"),
   950 => (x"20",x"20",x"3a",x"65"),
   951 => (x"0a",x"64",x"25",x"20"),
   952 => (x"00",x"00",x"00",x"00"),
   953 => (x"74",x"53",x"20",x"20"),
   954 => (x"6f",x"43",x"5f",x"72"),
   955 => (x"20",x"3a",x"70",x"6d"),
   956 => (x"20",x"20",x"20",x"20"),
   957 => (x"20",x"20",x"20",x"20"),
   958 => (x"0a",x"73",x"25",x"20"),
   959 => (x"00",x"00",x"00",x"00"),
   960 => (x"20",x"20",x"20",x"20"),
   961 => (x"20",x"20",x"20",x"20"),
   962 => (x"75",x"6f",x"68",x"73"),
   963 => (x"62",x"20",x"64",x"6c"),
   964 => (x"20",x"20",x"3a",x"65"),
   965 => (x"52",x"48",x"44",x"20"),
   966 => (x"4f",x"54",x"53",x"59"),
   967 => (x"50",x"20",x"45",x"4e"),
   968 => (x"52",x"47",x"4f",x"52"),
   969 => (x"20",x"2c",x"4d",x"41"),
   970 => (x"45",x"4d",x"4f",x"53"),
   971 => (x"52",x"54",x"53",x"20"),
   972 => (x"0a",x"47",x"4e",x"49"),
   973 => (x"00",x"00",x"00",x"00"),
   974 => (x"74",x"78",x"65",x"4e"),
   975 => (x"72",x"74",x"50",x"5f"),
   976 => (x"6f",x"6c",x"47",x"5f"),
   977 => (x"0a",x"3e",x"2d",x"62"),
   978 => (x"00",x"00",x"00",x"00"),
   979 => (x"74",x"50",x"20",x"20"),
   980 => (x"6f",x"43",x"5f",x"72"),
   981 => (x"20",x"3a",x"70",x"6d"),
   982 => (x"20",x"20",x"20",x"20"),
   983 => (x"20",x"20",x"20",x"20"),
   984 => (x"0a",x"64",x"25",x"20"),
   985 => (x"00",x"00",x"00",x"00"),
   986 => (x"20",x"20",x"20",x"20"),
   987 => (x"20",x"20",x"20",x"20"),
   988 => (x"75",x"6f",x"68",x"73"),
   989 => (x"62",x"20",x"64",x"6c"),
   990 => (x"20",x"20",x"3a",x"65"),
   991 => (x"6d",x"69",x"28",x"20"),
   992 => (x"6d",x"65",x"6c",x"70"),
   993 => (x"61",x"74",x"6e",x"65"),
   994 => (x"6e",x"6f",x"69",x"74"),
   995 => (x"70",x"65",x"64",x"2d"),
   996 => (x"65",x"64",x"6e",x"65"),
   997 => (x"2c",x"29",x"74",x"6e"),
   998 => (x"6d",x"61",x"73",x"20"),
   999 => (x"73",x"61",x"20",x"65"),
  1000 => (x"6f",x"62",x"61",x"20"),
  1001 => (x"00",x"0a",x"65",x"76"),
  1002 => (x"69",x"44",x"20",x"20"),
  1003 => (x"3a",x"72",x"63",x"73"),
  1004 => (x"20",x"20",x"20",x"20"),
  1005 => (x"20",x"20",x"20",x"20"),
  1006 => (x"20",x"20",x"20",x"20"),
  1007 => (x"0a",x"64",x"25",x"20"),
  1008 => (x"00",x"00",x"00",x"00"),
  1009 => (x"20",x"20",x"20",x"20"),
  1010 => (x"20",x"20",x"20",x"20"),
  1011 => (x"75",x"6f",x"68",x"73"),
  1012 => (x"62",x"20",x"64",x"6c"),
  1013 => (x"20",x"20",x"3a",x"65"),
  1014 => (x"0a",x"64",x"25",x"20"),
  1015 => (x"00",x"00",x"00",x"00"),
  1016 => (x"6e",x"45",x"20",x"20"),
  1017 => (x"43",x"5f",x"6d",x"75"),
  1018 => (x"3a",x"70",x"6d",x"6f"),
  1019 => (x"20",x"20",x"20",x"20"),
  1020 => (x"20",x"20",x"20",x"20"),
  1021 => (x"0a",x"64",x"25",x"20"),
  1022 => (x"00",x"00",x"00",x"00"),
  1023 => (x"20",x"20",x"20",x"20"),
  1024 => (x"20",x"20",x"20",x"20"),
  1025 => (x"75",x"6f",x"68",x"73"),
  1026 => (x"62",x"20",x"64",x"6c"),
  1027 => (x"20",x"20",x"3a",x"65"),
  1028 => (x"0a",x"64",x"25",x"20"),
  1029 => (x"00",x"00",x"00",x"00"),
  1030 => (x"6e",x"49",x"20",x"20"),
  1031 => (x"6f",x"43",x"5f",x"74"),
  1032 => (x"20",x"3a",x"70",x"6d"),
  1033 => (x"20",x"20",x"20",x"20"),
  1034 => (x"20",x"20",x"20",x"20"),
  1035 => (x"0a",x"64",x"25",x"20"),
  1036 => (x"00",x"00",x"00",x"00"),
  1037 => (x"20",x"20",x"20",x"20"),
  1038 => (x"20",x"20",x"20",x"20"),
  1039 => (x"75",x"6f",x"68",x"73"),
  1040 => (x"62",x"20",x"64",x"6c"),
  1041 => (x"20",x"20",x"3a",x"65"),
  1042 => (x"0a",x"64",x"25",x"20"),
  1043 => (x"00",x"00",x"00",x"00"),
  1044 => (x"74",x"53",x"20",x"20"),
  1045 => (x"6f",x"43",x"5f",x"72"),
  1046 => (x"20",x"3a",x"70",x"6d"),
  1047 => (x"20",x"20",x"20",x"20"),
  1048 => (x"20",x"20",x"20",x"20"),
  1049 => (x"0a",x"73",x"25",x"20"),
  1050 => (x"00",x"00",x"00",x"00"),
  1051 => (x"20",x"20",x"20",x"20"),
  1052 => (x"20",x"20",x"20",x"20"),
  1053 => (x"75",x"6f",x"68",x"73"),
  1054 => (x"62",x"20",x"64",x"6c"),
  1055 => (x"20",x"20",x"3a",x"65"),
  1056 => (x"52",x"48",x"44",x"20"),
  1057 => (x"4f",x"54",x"53",x"59"),
  1058 => (x"50",x"20",x"45",x"4e"),
  1059 => (x"52",x"47",x"4f",x"52"),
  1060 => (x"20",x"2c",x"4d",x"41"),
  1061 => (x"45",x"4d",x"4f",x"53"),
  1062 => (x"52",x"54",x"53",x"20"),
  1063 => (x"0a",x"47",x"4e",x"49"),
  1064 => (x"00",x"00",x"00",x"00"),
  1065 => (x"5f",x"74",x"6e",x"49"),
  1066 => (x"6f",x"4c",x"5f",x"31"),
  1067 => (x"20",x"20",x"3a",x"63"),
  1068 => (x"20",x"20",x"20",x"20"),
  1069 => (x"20",x"20",x"20",x"20"),
  1070 => (x"0a",x"64",x"25",x"20"),
  1071 => (x"00",x"00",x"00",x"00"),
  1072 => (x"20",x"20",x"20",x"20"),
  1073 => (x"20",x"20",x"20",x"20"),
  1074 => (x"75",x"6f",x"68",x"73"),
  1075 => (x"62",x"20",x"64",x"6c"),
  1076 => (x"20",x"20",x"3a",x"65"),
  1077 => (x"0a",x"64",x"25",x"20"),
  1078 => (x"00",x"00",x"00",x"00"),
  1079 => (x"5f",x"74",x"6e",x"49"),
  1080 => (x"6f",x"4c",x"5f",x"32"),
  1081 => (x"20",x"20",x"3a",x"63"),
  1082 => (x"20",x"20",x"20",x"20"),
  1083 => (x"20",x"20",x"20",x"20"),
  1084 => (x"0a",x"64",x"25",x"20"),
  1085 => (x"00",x"00",x"00",x"00"),
  1086 => (x"20",x"20",x"20",x"20"),
  1087 => (x"20",x"20",x"20",x"20"),
  1088 => (x"75",x"6f",x"68",x"73"),
  1089 => (x"62",x"20",x"64",x"6c"),
  1090 => (x"20",x"20",x"3a",x"65"),
  1091 => (x"0a",x"64",x"25",x"20"),
  1092 => (x"00",x"00",x"00",x"00"),
  1093 => (x"5f",x"74",x"6e",x"49"),
  1094 => (x"6f",x"4c",x"5f",x"33"),
  1095 => (x"20",x"20",x"3a",x"63"),
  1096 => (x"20",x"20",x"20",x"20"),
  1097 => (x"20",x"20",x"20",x"20"),
  1098 => (x"0a",x"64",x"25",x"20"),
  1099 => (x"00",x"00",x"00",x"00"),
  1100 => (x"20",x"20",x"20",x"20"),
  1101 => (x"20",x"20",x"20",x"20"),
  1102 => (x"75",x"6f",x"68",x"73"),
  1103 => (x"62",x"20",x"64",x"6c"),
  1104 => (x"20",x"20",x"3a",x"65"),
  1105 => (x"0a",x"64",x"25",x"20"),
  1106 => (x"00",x"00",x"00",x"00"),
  1107 => (x"6d",x"75",x"6e",x"45"),
  1108 => (x"63",x"6f",x"4c",x"5f"),
  1109 => (x"20",x"20",x"20",x"3a"),
  1110 => (x"20",x"20",x"20",x"20"),
  1111 => (x"20",x"20",x"20",x"20"),
  1112 => (x"0a",x"64",x"25",x"20"),
  1113 => (x"00",x"00",x"00",x"00"),
  1114 => (x"20",x"20",x"20",x"20"),
  1115 => (x"20",x"20",x"20",x"20"),
  1116 => (x"75",x"6f",x"68",x"73"),
  1117 => (x"62",x"20",x"64",x"6c"),
  1118 => (x"20",x"20",x"3a",x"65"),
  1119 => (x"0a",x"64",x"25",x"20"),
  1120 => (x"00",x"00",x"00",x"00"),
  1121 => (x"5f",x"72",x"74",x"53"),
  1122 => (x"6f",x"4c",x"5f",x"31"),
  1123 => (x"20",x"20",x"3a",x"63"),
  1124 => (x"20",x"20",x"20",x"20"),
  1125 => (x"20",x"20",x"20",x"20"),
  1126 => (x"0a",x"73",x"25",x"20"),
  1127 => (x"00",x"00",x"00",x"00"),
  1128 => (x"20",x"20",x"20",x"20"),
  1129 => (x"20",x"20",x"20",x"20"),
  1130 => (x"75",x"6f",x"68",x"73"),
  1131 => (x"62",x"20",x"64",x"6c"),
  1132 => (x"20",x"20",x"3a",x"65"),
  1133 => (x"52",x"48",x"44",x"20"),
  1134 => (x"4f",x"54",x"53",x"59"),
  1135 => (x"50",x"20",x"45",x"4e"),
  1136 => (x"52",x"47",x"4f",x"52"),
  1137 => (x"20",x"2c",x"4d",x"41"),
  1138 => (x"54",x"53",x"27",x"31"),
  1139 => (x"52",x"54",x"53",x"20"),
  1140 => (x"0a",x"47",x"4e",x"49"),
  1141 => (x"00",x"00",x"00",x"00"),
  1142 => (x"5f",x"72",x"74",x"53"),
  1143 => (x"6f",x"4c",x"5f",x"32"),
  1144 => (x"20",x"20",x"3a",x"63"),
  1145 => (x"20",x"20",x"20",x"20"),
  1146 => (x"20",x"20",x"20",x"20"),
  1147 => (x"0a",x"73",x"25",x"20"),
  1148 => (x"00",x"00",x"00",x"00"),
  1149 => (x"20",x"20",x"20",x"20"),
  1150 => (x"20",x"20",x"20",x"20"),
  1151 => (x"75",x"6f",x"68",x"73"),
  1152 => (x"62",x"20",x"64",x"6c"),
  1153 => (x"20",x"20",x"3a",x"65"),
  1154 => (x"52",x"48",x"44",x"20"),
  1155 => (x"4f",x"54",x"53",x"59"),
  1156 => (x"50",x"20",x"45",x"4e"),
  1157 => (x"52",x"47",x"4f",x"52"),
  1158 => (x"20",x"2c",x"4d",x"41"),
  1159 => (x"44",x"4e",x"27",x"32"),
  1160 => (x"52",x"54",x"53",x"20"),
  1161 => (x"0a",x"47",x"4e",x"49"),
  1162 => (x"00",x"00",x"00",x"00"),
  1163 => (x"00",x"00",x"00",x"0a"),
  1164 => (x"72",x"65",x"73",x"55"),
  1165 => (x"6d",x"69",x"74",x"20"),
  1166 => (x"25",x"20",x"3a",x"65"),
  1167 => (x"1e",x"00",x"0a",x"64"),
  1168 => (x"1e",x"74",x"1e",x"73"),
  1169 => (x"66",x"cc",x"4b",x"71"),
  1170 => (x"c2",x"7a",x"73",x"4a"),
  1171 => (x"87",x"c4",x"05",x"ab"),
  1172 => (x"87",x"c2",x"4c",x"c1"),
  1173 => (x"9c",x"74",x"4c",x"c0"),
  1174 => (x"c3",x"87",x"c2",x"05"),
  1175 => (x"02",x"9b",x"73",x"7a"),
  1176 => (x"c1",x"49",x"87",x"d6"),
  1177 => (x"87",x"d4",x"02",x"89"),
  1178 => (x"e3",x"c0",x"02",x"89"),
  1179 => (x"c0",x"02",x"89",x"87"),
  1180 => (x"02",x"89",x"87",x"e4"),
  1181 => (x"87",x"de",x"87",x"de"),
  1182 => (x"87",x"da",x"7a",x"c0"),
  1183 => (x"bf",x"e4",x"cf",x"c1"),
  1184 => (x"b7",x"e4",x"c1",x"48"),
  1185 => (x"87",x"c4",x"06",x"a8"),
  1186 => (x"87",x"ca",x"7a",x"c0"),
  1187 => (x"87",x"c6",x"7a",x"c3"),
  1188 => (x"87",x"c2",x"7a",x"c1"),
  1189 => (x"4c",x"26",x"7a",x"c2"),
  1190 => (x"4f",x"26",x"4b",x"26"),
  1191 => (x"49",x"4a",x"71",x"1e"),
  1192 => (x"66",x"c4",x"81",x"c2"),
  1193 => (x"c8",x"80",x"71",x"48"),
  1194 => (x"08",x"78",x"08",x"66"),
  1195 => (x"5e",x"0e",x"4f",x"26"),
  1196 => (x"0e",x"5d",x"5c",x"5b"),
  1197 => (x"a6",x"c4",x"86",x"f4"),
  1198 => (x"66",x"e0",x"c0",x"59"),
  1199 => (x"74",x"84",x"c5",x"4c"),
  1200 => (x"c8",x"90",x"c4",x"48"),
  1201 => (x"4d",x"6e",x"58",x"a6"),
  1202 => (x"e4",x"c0",x"85",x"70"),
  1203 => (x"a5",x"c4",x"7d",x"66"),
  1204 => (x"66",x"e4",x"c0",x"49"),
  1205 => (x"a5",x"f8",x"c1",x"79"),
  1206 => (x"c8",x"79",x"74",x"49"),
  1207 => (x"a4",x"c1",x"48",x"a6"),
  1208 => (x"01",x"ac",x"b7",x"78"),
  1209 => (x"49",x"74",x"87",x"dd"),
  1210 => (x"dc",x"91",x"c8",x"c3"),
  1211 => (x"82",x"71",x"4a",x"66"),
  1212 => (x"c8",x"82",x"66",x"c4"),
  1213 => (x"8b",x"74",x"4b",x"66"),
  1214 => (x"7a",x"74",x"83",x"c1"),
  1215 => (x"8b",x"c1",x"82",x"c4"),
  1216 => (x"74",x"87",x"f7",x"01"),
  1217 => (x"91",x"c8",x"c3",x"49"),
  1218 => (x"71",x"81",x"66",x"dc"),
  1219 => (x"82",x"66",x"c4",x"4a"),
  1220 => (x"48",x"6a",x"8a",x"c4"),
  1221 => (x"7a",x"70",x"80",x"c1"),
  1222 => (x"81",x"e0",x"fe",x"c0"),
  1223 => (x"6d",x"81",x"66",x"c4"),
  1224 => (x"e4",x"cf",x"c1",x"79"),
  1225 => (x"f4",x"78",x"c5",x"48"),
  1226 => (x"26",x"4d",x"26",x"8e"),
  1227 => (x"26",x"4b",x"26",x"4c"),
  1228 => (x"1e",x"73",x"1e",x"4f"),
  1229 => (x"4b",x"71",x"1e",x"74"),
  1230 => (x"66",x"cc",x"4a",x"4c"),
  1231 => (x"02",x"aa",x"b7",x"49"),
  1232 => (x"48",x"c0",x"87",x"c4"),
  1233 => (x"cf",x"c1",x"87",x"c7"),
  1234 => (x"c1",x"5c",x"97",x"f0"),
  1235 => (x"26",x"4c",x"26",x"48"),
  1236 => (x"0e",x"4f",x"26",x"4b"),
  1237 => (x"5d",x"5c",x"5b",x"5e"),
  1238 => (x"c4",x"86",x"f4",x"0e"),
  1239 => (x"4d",x"c2",x"59",x"a6"),
  1240 => (x"c1",x"49",x"66",x"dc"),
  1241 => (x"c2",x"4c",x"6e",x"81"),
  1242 => (x"6b",x"4b",x"a1",x"84"),
  1243 => (x"99",x"ff",x"c3",x"49"),
  1244 => (x"6c",x"48",x"a6",x"c4"),
  1245 => (x"66",x"97",x"c4",x"50"),
  1246 => (x"aa",x"b7",x"71",x"4a"),
  1247 => (x"c8",x"87",x"c7",x"02"),
  1248 => (x"78",x"c0",x"48",x"a6"),
  1249 => (x"cf",x"c1",x"87",x"cd"),
  1250 => (x"97",x"c4",x"48",x"ec"),
  1251 => (x"a6",x"c8",x"50",x"66"),
  1252 => (x"c8",x"78",x"c1",x"48"),
  1253 => (x"87",x"c4",x"05",x"66"),
  1254 => (x"84",x"83",x"85",x"c1"),
  1255 => (x"06",x"ad",x"b7",x"c2"),
  1256 => (x"6e",x"87",x"c8",x"ff"),
  1257 => (x"49",x"66",x"dc",x"4a"),
  1258 => (x"87",x"f0",x"fe",x"fe"),
  1259 => (x"06",x"a8",x"b7",x"c0"),
  1260 => (x"cf",x"c1",x"87",x"cb"),
  1261 => (x"a5",x"c7",x"48",x"e4"),
  1262 => (x"c2",x"48",x"c1",x"78"),
  1263 => (x"f4",x"48",x"c0",x"87"),
  1264 => (x"26",x"4d",x"26",x"8e"),
  1265 => (x"26",x"4b",x"26",x"4c"),
  1266 => (x"26",x"4b",x"26",x"4f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
