
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"c9",x"01"),
     1 => (x"cf",x"03",x"87",x"cc"),
     2 => (x"87",x"fd",x"00",x"87"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"36",x"27",x"4f",x"00"),
     5 => (x"4f",x"00",x"00",x"00"),
     6 => (x"0e",x"1e",x"18",x"0e"),
     7 => (x"00",x"00",x"44",x"27"),
     8 => (x"48",x"26",x"0f",x"00"),
     9 => (x"08",x"26",x"80",x"ff"),
    10 => (x"c0",x"c0",x"c2",x"4f"),
    11 => (x"05",x"3a",x"27",x"4e"),
    12 => (x"00",x"0f",x"00",x"00"),
    13 => (x"f0",x"c1",x"87",x"fd"),
    14 => (x"43",x"27",x"4e",x"c0"),
    15 => (x"0f",x"00",x"00",x"00"),
    16 => (x"4f",x"87",x"fd",x"00"),
    17 => (x"0e",x"1e",x"18",x"0e"),
    18 => (x"80",x"ff",x"48",x"26"),
    19 => (x"1e",x"4f",x"08",x"26"),
    20 => (x"ff",x"1e",x"1e",x"72"),
    21 => (x"48",x"6a",x"4a",x"c0"),
    22 => (x"c4",x"98",x"c0",x"c4"),
    23 => (x"02",x"6e",x"58",x"a6"),
    24 => (x"cc",x"87",x"f3",x"ff"),
    25 => (x"66",x"cc",x"7a",x"66"),
    26 => (x"4a",x"26",x"26",x"48"),
    27 => (x"5e",x"0e",x"4f",x"26"),
    28 => (x"5d",x"5c",x"5b",x"5a"),
    29 => (x"4b",x"66",x"d4",x"0e"),
    30 => (x"4c",x"13",x"4d",x"c0"),
    31 => (x"c0",x"02",x"9c",x"74"),
    32 => (x"4a",x"74",x"87",x"d6"),
    33 => (x"4f",x"27",x"1e",x"72"),
    34 => (x"0f",x"00",x"00",x"00"),
    35 => (x"85",x"c1",x"86",x"c4"),
    36 => (x"9c",x"74",x"4c",x"13"),
    37 => (x"87",x"ea",x"ff",x"05"),
    38 => (x"4d",x"26",x"48",x"75"),
    39 => (x"4b",x"26",x"4c",x"26"),
    40 => (x"4f",x"26",x"4a",x"26"),
    41 => (x"5b",x"5a",x"5e",x"0e"),
    42 => (x"c8",x"0e",x"5d",x"5c"),
    43 => (x"66",x"e0",x"c0",x"8e"),
    44 => (x"4c",x"66",x"dc",x"4d"),
    45 => (x"00",x"16",x"90",x"27"),
    46 => (x"49",x"76",x"4b",x"00"),
    47 => (x"00",x"0e",x"d4",x"27"),
    48 => (x"a6",x"c4",x"79",x"00"),
    49 => (x"c0",x"79",x"c0",x"49"),
    50 => (x"c0",x"03",x"ac",x"b7"),
    51 => (x"ed",x"c0",x"87",x"ce"),
    52 => (x"00",x"4f",x"27",x"1e"),
    53 => (x"c4",x"0f",x"00",x"00"),
    54 => (x"8c",x"0c",x"c0",x"86"),
    55 => (x"c0",x"05",x"9c",x"74"),
    56 => (x"f0",x"c0",x"87",x"c6"),
    57 => (x"87",x"f6",x"c0",x"53"),
    58 => (x"c0",x"02",x"9c",x"74"),
    59 => (x"49",x"74",x"87",x"f0"),
    60 => (x"e8",x"c0",x"1e",x"72"),
    61 => (x"db",x"27",x"4a",x"66"),
    62 => (x"0f",x"00",x"00",x"04"),
    63 => (x"4a",x"71",x"4a",x"26"),
    64 => (x"82",x"6e",x"4a",x"72"),
    65 => (x"49",x"74",x"53",x"12"),
    66 => (x"e8",x"c0",x"1e",x"72"),
    67 => (x"db",x"27",x"4a",x"66"),
    68 => (x"0f",x"00",x"00",x"04"),
    69 => (x"4c",x"70",x"4a",x"26"),
    70 => (x"ff",x"05",x"9c",x"74"),
    71 => (x"90",x"27",x"87",x"d0"),
    72 => (x"b7",x"00",x"00",x"16"),
    73 => (x"d8",x"c0",x"02",x"ab"),
    74 => (x"97",x"8b",x"c1",x"87"),
    75 => (x"66",x"c4",x"55",x"6b"),
    76 => (x"c8",x"80",x"c1",x"48"),
    77 => (x"90",x"27",x"58",x"a6"),
    78 => (x"b7",x"00",x"00",x"16"),
    79 => (x"e8",x"ff",x"05",x"ab"),
    80 => (x"c4",x"55",x"c0",x"87"),
    81 => (x"86",x"c8",x"48",x"66"),
    82 => (x"4c",x"26",x"4d",x"26"),
    83 => (x"4a",x"26",x"4b",x"26"),
    84 => (x"5e",x"0e",x"4f",x"26"),
    85 => (x"5d",x"5c",x"5b",x"5a"),
    86 => (x"4c",x"c0",x"1e",x"0e"),
    87 => (x"79",x"c0",x"49",x"76"),
    88 => (x"d8",x"4b",x"a6",x"dc"),
    89 => (x"66",x"d8",x"4a",x"66"),
    90 => (x"dc",x"80",x"c1",x"48"),
    91 => (x"4d",x"12",x"58",x"a6"),
    92 => (x"c0",x"c0",x"c0",x"c1"),
    93 => (x"c0",x"c4",x"95",x"c0"),
    94 => (x"75",x"4d",x"95",x"b7"),
    95 => (x"d2",x"c4",x"02",x"9d"),
    96 => (x"c3",x"02",x"6e",x"87"),
    97 => (x"49",x"76",x"87",x"d7"),
    98 => (x"4a",x"75",x"79",x"c0"),
    99 => (x"02",x"ad",x"e3",x"c1"),
   100 => (x"c1",x"87",x"dd",x"c2"),
   101 => (x"c0",x"02",x"aa",x"e4"),
   102 => (x"ec",x"c1",x"87",x"d8"),
   103 => (x"c8",x"c2",x"02",x"aa"),
   104 => (x"aa",x"f3",x"c1",x"87"),
   105 => (x"87",x"e8",x"c1",x"02"),
   106 => (x"02",x"aa",x"f8",x"c1"),
   107 => (x"c2",x"87",x"f2",x"c0"),
   108 => (x"1e",x"ca",x"87",x"d3"),
   109 => (x"00",x"16",x"e0",x"27"),
   110 => (x"83",x"c4",x"1e",x"00"),
   111 => (x"8a",x"c4",x"4a",x"73"),
   112 => (x"a4",x"27",x"1e",x"6a"),
   113 => (x"0f",x"00",x"00",x"00"),
   114 => (x"4a",x"70",x"86",x"cc"),
   115 => (x"84",x"72",x"4c",x"74"),
   116 => (x"00",x"16",x"e0",x"27"),
   117 => (x"6e",x"27",x"1e",x"00"),
   118 => (x"0f",x"00",x"00",x"00"),
   119 => (x"d4",x"c2",x"86",x"c4"),
   120 => (x"27",x"1e",x"d0",x"87"),
   121 => (x"00",x"00",x"16",x"e0"),
   122 => (x"73",x"83",x"c4",x"1e"),
   123 => (x"6a",x"8a",x"c4",x"4a"),
   124 => (x"00",x"a4",x"27",x"1e"),
   125 => (x"cc",x"0f",x"00",x"00"),
   126 => (x"74",x"4a",x"70",x"86"),
   127 => (x"27",x"84",x"72",x"4c"),
   128 => (x"00",x"00",x"16",x"e0"),
   129 => (x"00",x"6e",x"27",x"1e"),
   130 => (x"c4",x"0f",x"00",x"00"),
   131 => (x"87",x"e5",x"c1",x"86"),
   132 => (x"4a",x"73",x"83",x"c4"),
   133 => (x"1e",x"6a",x"8a",x"c4"),
   134 => (x"00",x"00",x"6e",x"27"),
   135 => (x"86",x"c4",x"0f",x"00"),
   136 => (x"4c",x"74",x"4a",x"70"),
   137 => (x"cc",x"c1",x"84",x"72"),
   138 => (x"c1",x"49",x"76",x"87"),
   139 => (x"87",x"c5",x"c1",x"79"),
   140 => (x"4a",x"73",x"83",x"c4"),
   141 => (x"1e",x"6a",x"8a",x"c4"),
   142 => (x"00",x"00",x"4f",x"27"),
   143 => (x"86",x"c4",x"0f",x"00"),
   144 => (x"f0",x"c0",x"84",x"c1"),
   145 => (x"1e",x"e5",x"c0",x"87"),
   146 => (x"00",x"00",x"4f",x"27"),
   147 => (x"86",x"c4",x"0f",x"00"),
   148 => (x"4f",x"27",x"1e",x"75"),
   149 => (x"0f",x"00",x"00",x"00"),
   150 => (x"d8",x"c0",x"86",x"c4"),
   151 => (x"ad",x"e5",x"c0",x"87"),
   152 => (x"87",x"c7",x"c0",x"05"),
   153 => (x"79",x"c1",x"49",x"76"),
   154 => (x"75",x"87",x"ca",x"c0"),
   155 => (x"00",x"4f",x"27",x"1e"),
   156 => (x"c4",x"0f",x"00",x"00"),
   157 => (x"4a",x"66",x"d8",x"86"),
   158 => (x"c1",x"48",x"66",x"d8"),
   159 => (x"58",x"a6",x"dc",x"80"),
   160 => (x"c0",x"c1",x"4d",x"12"),
   161 => (x"95",x"c0",x"c0",x"c0"),
   162 => (x"95",x"b7",x"c0",x"c4"),
   163 => (x"05",x"9d",x"75",x"4d"),
   164 => (x"74",x"87",x"ee",x"fb"),
   165 => (x"4d",x"26",x"26",x"48"),
   166 => (x"4b",x"26",x"4c",x"26"),
   167 => (x"4f",x"26",x"4a",x"26"),
   168 => (x"5b",x"5a",x"5e",x"0e"),
   169 => (x"4b",x"66",x"d0",x"0e"),
   170 => (x"cc",x"7b",x"66",x"cc"),
   171 => (x"c7",x"27",x"1e",x"66"),
   172 => (x"0f",x"00",x"00",x"04"),
   173 => (x"4a",x"70",x"86",x"c4"),
   174 => (x"c0",x"05",x"9a",x"72"),
   175 => (x"7b",x"c3",x"87",x"c2"),
   176 => (x"cc",x"4a",x"66",x"cc"),
   177 => (x"b7",x"c0",x"49",x"66"),
   178 => (x"df",x"c0",x"02",x"a9"),
   179 => (x"aa",x"b7",x"c1",x"87"),
   180 => (x"87",x"dd",x"c0",x"02"),
   181 => (x"02",x"aa",x"b7",x"c2"),
   182 => (x"c3",x"87",x"ef",x"c0"),
   183 => (x"c0",x"02",x"aa",x"b7"),
   184 => (x"b7",x"c4",x"87",x"ef"),
   185 => (x"e6",x"c0",x"02",x"aa"),
   186 => (x"87",x"e5",x"c0",x"87"),
   187 => (x"e0",x"c0",x"7b",x"c0"),
   188 => (x"17",x"08",x"27",x"87"),
   189 => (x"49",x"bf",x"00",x"00"),
   190 => (x"a9",x"b7",x"e4",x"c1"),
   191 => (x"87",x"c5",x"c0",x"06"),
   192 => (x"cc",x"c0",x"7b",x"c0"),
   193 => (x"c0",x"7b",x"c3",x"87"),
   194 => (x"7b",x"c1",x"87",x"c7"),
   195 => (x"c2",x"87",x"c2",x"c0"),
   196 => (x"26",x"4b",x"26",x"7b"),
   197 => (x"1e",x"4f",x"26",x"4a"),
   198 => (x"66",x"c8",x"1e",x"72"),
   199 => (x"cc",x"82",x"c2",x"4a"),
   200 => (x"80",x"72",x"48",x"66"),
   201 => (x"70",x"49",x"66",x"d0"),
   202 => (x"26",x"4a",x"26",x"79"),
   203 => (x"5a",x"5e",x"0e",x"4f"),
   204 => (x"0e",x"5d",x"5c",x"5b"),
   205 => (x"c5",x"4d",x"66",x"dc"),
   206 => (x"c4",x"4a",x"75",x"85"),
   207 => (x"d4",x"4a",x"72",x"92"),
   208 => (x"e0",x"c0",x"82",x"66"),
   209 => (x"4b",x"72",x"7a",x"66"),
   210 => (x"7b",x"6a",x"83",x"c4"),
   211 => (x"75",x"82",x"f8",x"c1"),
   212 => (x"75",x"4c",x"75",x"7a"),
   213 => (x"72",x"82",x"c1",x"4a"),
   214 => (x"c0",x"01",x"ad",x"b7"),
   215 => (x"4b",x"75",x"87",x"e1"),
   216 => (x"73",x"93",x"c8",x"c3"),
   217 => (x"83",x"66",x"d8",x"4b"),
   218 => (x"92",x"c4",x"4a",x"74"),
   219 => (x"82",x"73",x"4a",x"72"),
   220 => (x"84",x"c1",x"7a",x"75"),
   221 => (x"82",x"c1",x"4a",x"75"),
   222 => (x"06",x"ac",x"b7",x"72"),
   223 => (x"75",x"87",x"df",x"ff"),
   224 => (x"94",x"c8",x"c3",x"4c"),
   225 => (x"66",x"d8",x"4c",x"74"),
   226 => (x"c4",x"4a",x"75",x"84"),
   227 => (x"72",x"4b",x"74",x"92"),
   228 => (x"6b",x"8b",x"c4",x"83"),
   229 => (x"70",x"80",x"c1",x"48"),
   230 => (x"4b",x"66",x"d4",x"7b"),
   231 => (x"fe",x"c0",x"83",x"72"),
   232 => (x"4a",x"72",x"84",x"e0"),
   233 => (x"7a",x"6b",x"82",x"74"),
   234 => (x"00",x"17",x"08",x"27"),
   235 => (x"79",x"c5",x"49",x"00"),
   236 => (x"4c",x"26",x"4d",x"26"),
   237 => (x"4a",x"26",x"4b",x"26"),
   238 => (x"5e",x"0e",x"4f",x"26"),
   239 => (x"0e",x"5c",x"5b",x"5a"),
   240 => (x"4c",x"66",x"d0",x"97"),
   241 => (x"c0",x"c1",x"4b",x"74"),
   242 => (x"93",x"c0",x"c0",x"c0"),
   243 => (x"93",x"b7",x"c0",x"c4"),
   244 => (x"66",x"d4",x"97",x"4b"),
   245 => (x"c0",x"c0",x"c1",x"4a"),
   246 => (x"c4",x"92",x"c0",x"c0"),
   247 => (x"4a",x"92",x"b7",x"c0"),
   248 => (x"02",x"ab",x"b7",x"72"),
   249 => (x"c0",x"87",x"c5",x"c0"),
   250 => (x"87",x"ca",x"c0",x"48"),
   251 => (x"00",x"17",x"10",x"27"),
   252 => (x"51",x"74",x"49",x"00"),
   253 => (x"4c",x"26",x"48",x"c1"),
   254 => (x"4a",x"26",x"4b",x"26"),
   255 => (x"5e",x"0e",x"4f",x"26"),
   256 => (x"0e",x"5c",x"5b",x"5a"),
   257 => (x"4c",x"6e",x"97",x"1e"),
   258 => (x"66",x"d8",x"4b",x"c2"),
   259 => (x"73",x"82",x"c1",x"4a"),
   260 => (x"4a",x"6a",x"97",x"82"),
   261 => (x"c0",x"c0",x"c0",x"c1"),
   262 => (x"c0",x"c4",x"92",x"c0"),
   263 => (x"72",x"4a",x"92",x"b7"),
   264 => (x"4a",x"66",x"d8",x"1e"),
   265 => (x"6a",x"97",x"82",x"73"),
   266 => (x"c0",x"c0",x"c1",x"4a"),
   267 => (x"c4",x"92",x"c0",x"c0"),
   268 => (x"4a",x"92",x"b7",x"c0"),
   269 => (x"ba",x"27",x"1e",x"72"),
   270 => (x"0f",x"00",x"00",x"03"),
   271 => (x"4a",x"70",x"86",x"c8"),
   272 => (x"c0",x"05",x"9a",x"72"),
   273 => (x"c1",x"c1",x"87",x"c5"),
   274 => (x"c2",x"83",x"c1",x"4c"),
   275 => (x"fe",x"06",x"ab",x"b7"),
   276 => (x"4a",x"74",x"87",x"f8"),
   277 => (x"c0",x"c0",x"c0",x"c1"),
   278 => (x"c0",x"c4",x"92",x"c0"),
   279 => (x"c1",x"4a",x"92",x"b7"),
   280 => (x"04",x"aa",x"b7",x"d7"),
   281 => (x"74",x"87",x"d7",x"c0"),
   282 => (x"c0",x"c0",x"c1",x"4a"),
   283 => (x"c4",x"92",x"c0",x"c0"),
   284 => (x"4a",x"92",x"b7",x"c0"),
   285 => (x"aa",x"b7",x"da",x"c1"),
   286 => (x"87",x"c2",x"c0",x"03"),
   287 => (x"4a",x"74",x"4b",x"c7"),
   288 => (x"c0",x"c0",x"c0",x"c1"),
   289 => (x"c0",x"c4",x"92",x"c0"),
   290 => (x"c1",x"4a",x"92",x"b7"),
   291 => (x"05",x"aa",x"b7",x"d2"),
   292 => (x"c1",x"87",x"c5",x"c0"),
   293 => (x"87",x"e6",x"c0",x"48"),
   294 => (x"d8",x"4a",x"66",x"d4"),
   295 => (x"25",x"27",x"49",x"66"),
   296 => (x"0f",x"00",x"00",x"05"),
   297 => (x"b7",x"c0",x"4a",x"70"),
   298 => (x"cf",x"c0",x"06",x"aa"),
   299 => (x"c7",x"48",x"73",x"87"),
   300 => (x"17",x"0c",x"27",x"80"),
   301 => (x"c1",x"58",x"00",x"00"),
   302 => (x"87",x"c2",x"c0",x"48"),
   303 => (x"26",x"26",x"48",x"c0"),
   304 => (x"26",x"4b",x"26",x"4c"),
   305 => (x"1e",x"4f",x"26",x"4a"),
   306 => (x"c2",x"49",x"66",x"c4"),
   307 => (x"c0",x"05",x"a9",x"b7"),
   308 => (x"48",x"c1",x"87",x"c5"),
   309 => (x"c0",x"87",x"c2",x"c0"),
   310 => (x"1e",x"4f",x"26",x"48"),
   311 => (x"9a",x"72",x"1e",x"73"),
   312 => (x"c0",x"87",x"d9",x"02"),
   313 => (x"72",x"4b",x"c1",x"48"),
   314 => (x"73",x"82",x"01",x"a9"),
   315 => (x"72",x"87",x"f8",x"83"),
   316 => (x"73",x"89",x"03",x"a9"),
   317 => (x"2a",x"c1",x"07",x"80"),
   318 => (x"87",x"f3",x"05",x"2b"),
   319 => (x"4f",x"26",x"4b",x"26"),
   320 => (x"c0",x"1e",x"75",x"1e"),
   321 => (x"04",x"a1",x"71",x"4d"),
   322 => (x"81",x"c1",x"b9",x"ff"),
   323 => (x"a2",x"72",x"07",x"bd"),
   324 => (x"c1",x"ba",x"ff",x"04"),
   325 => (x"c2",x"07",x"bd",x"82"),
   326 => (x"05",x"9d",x"75",x"87"),
   327 => (x"80",x"c1",x"b8",x"ff"),
   328 => (x"26",x"4d",x"25",x"07"),
   329 => (x"48",x"12",x"1e",x"4f"),
   330 => (x"87",x"c4",x"02",x"11"),
   331 => (x"87",x"f6",x"02",x"88"),
   332 => (x"ff",x"1e",x"4f",x"26"),
   333 => (x"48",x"68",x"48",x"c8"),
   334 => (x"5e",x"0e",x"4f",x"26"),
   335 => (x"5d",x"5c",x"5b",x"5a"),
   336 => (x"c4",x"8e",x"d0",x"0e"),
   337 => (x"04",x"27",x"4c",x"66"),
   338 => (x"49",x"00",x"00",x"17"),
   339 => (x"00",x"3f",x"08",x"27"),
   340 => (x"00",x"27",x"79",x"00"),
   341 => (x"49",x"00",x"00",x"17"),
   342 => (x"00",x"3f",x"38",x"27"),
   343 => (x"38",x"27",x"79",x"00"),
   344 => (x"49",x"00",x"00",x"3f"),
   345 => (x"00",x"3f",x"08",x"27"),
   346 => (x"3c",x"27",x"79",x"00"),
   347 => (x"49",x"00",x"00",x"3f"),
   348 => (x"40",x"27",x"79",x"c0"),
   349 => (x"49",x"00",x"00",x"3f"),
   350 => (x"44",x"27",x"79",x"c2"),
   351 => (x"49",x"00",x"00",x"3f"),
   352 => (x"27",x"79",x"e8",x"c0"),
   353 => (x"00",x"00",x"3f",x"48"),
   354 => (x"10",x"5e",x"27",x"49"),
   355 => (x"72",x"48",x"00",x"00"),
   356 => (x"c4",x"79",x"20",x"1e"),
   357 => (x"c4",x"79",x"20",x"81"),
   358 => (x"c4",x"79",x"20",x"81"),
   359 => (x"c4",x"79",x"20",x"81"),
   360 => (x"c4",x"79",x"20",x"81"),
   361 => (x"c4",x"79",x"20",x"81"),
   362 => (x"c4",x"79",x"20",x"81"),
   363 => (x"10",x"51",x"10",x"81"),
   364 => (x"26",x"51",x"10",x"51"),
   365 => (x"3f",x"68",x"27",x"4a"),
   366 => (x"27",x"49",x"00",x"00"),
   367 => (x"00",x"00",x"10",x"7d"),
   368 => (x"20",x"1e",x"72",x"48"),
   369 => (x"20",x"81",x"c4",x"79"),
   370 => (x"20",x"81",x"c4",x"79"),
   371 => (x"20",x"81",x"c4",x"79"),
   372 => (x"20",x"81",x"c4",x"79"),
   373 => (x"20",x"81",x"c4",x"79"),
   374 => (x"20",x"81",x"c4",x"79"),
   375 => (x"10",x"81",x"c4",x"79"),
   376 => (x"10",x"51",x"10",x"51"),
   377 => (x"27",x"4a",x"26",x"51"),
   378 => (x"00",x"00",x"1e",x"3c"),
   379 => (x"27",x"79",x"ca",x"49"),
   380 => (x"00",x"00",x"10",x"9c"),
   381 => (x"01",x"52",x"27",x"1e"),
   382 => (x"c4",x"0f",x"00",x"00"),
   383 => (x"10",x"9e",x"27",x"86"),
   384 => (x"27",x"1e",x"00",x"00"),
   385 => (x"00",x"00",x"01",x"52"),
   386 => (x"27",x"86",x"c4",x"0f"),
   387 => (x"00",x"00",x"10",x"ce"),
   388 => (x"01",x"52",x"27",x"1e"),
   389 => (x"c4",x"0f",x"00",x"00"),
   390 => (x"16",x"84",x"27",x"86"),
   391 => (x"02",x"bf",x"00",x"00"),
   392 => (x"27",x"87",x"df",x"c0"),
   393 => (x"00",x"00",x"0e",x"e5"),
   394 => (x"01",x"52",x"27",x"1e"),
   395 => (x"c4",x"0f",x"00",x"00"),
   396 => (x"0f",x"11",x"27",x"86"),
   397 => (x"27",x"1e",x"00",x"00"),
   398 => (x"00",x"00",x"01",x"52"),
   399 => (x"c0",x"86",x"c4",x"0f"),
   400 => (x"13",x"27",x"87",x"dc"),
   401 => (x"1e",x"00",x"00",x"0f"),
   402 => (x"00",x"01",x"52",x"27"),
   403 => (x"86",x"c4",x"0f",x"00"),
   404 => (x"00",x"0f",x"42",x"27"),
   405 => (x"52",x"27",x"1e",x"00"),
   406 => (x"0f",x"00",x"00",x"01"),
   407 => (x"88",x"27",x"86",x"c4"),
   408 => (x"bf",x"00",x"00",x"16"),
   409 => (x"10",x"d0",x"27",x"1e"),
   410 => (x"27",x"1e",x"00",x"00"),
   411 => (x"00",x"00",x"01",x"52"),
   412 => (x"27",x"86",x"c8",x"0f"),
   413 => (x"00",x"00",x"05",x"32"),
   414 => (x"3e",x"f4",x"27",x"0f"),
   415 => (x"c1",x"58",x"00",x"00"),
   416 => (x"16",x"88",x"27",x"4d"),
   417 => (x"49",x"bf",x"00",x"00"),
   418 => (x"06",x"a9",x"b7",x"c0"),
   419 => (x"27",x"87",x"d5",x"c7"),
   420 => (x"00",x"00",x"0e",x"bf"),
   421 => (x"0e",x"7e",x"27",x"0f"),
   422 => (x"76",x"0f",x"00",x"00"),
   423 => (x"c3",x"79",x"c2",x"49"),
   424 => (x"3f",x"88",x"27",x"4c"),
   425 => (x"27",x"49",x"00",x"00"),
   426 => (x"00",x"00",x"0f",x"63"),
   427 => (x"20",x"1e",x"72",x"48"),
   428 => (x"20",x"81",x"c4",x"79"),
   429 => (x"20",x"81",x"c4",x"79"),
   430 => (x"20",x"81",x"c4",x"79"),
   431 => (x"20",x"81",x"c4",x"79"),
   432 => (x"20",x"81",x"c4",x"79"),
   433 => (x"20",x"81",x"c4",x"79"),
   434 => (x"10",x"81",x"c4",x"79"),
   435 => (x"10",x"51",x"10",x"51"),
   436 => (x"c8",x"4a",x"26",x"51"),
   437 => (x"79",x"c1",x"49",x"a6"),
   438 => (x"00",x"3f",x"88",x"27"),
   439 => (x"68",x"27",x"1e",x"00"),
   440 => (x"1e",x"00",x"00",x"3f"),
   441 => (x"00",x"03",x"fe",x"27"),
   442 => (x"86",x"c8",x"0f",x"00"),
   443 => (x"9a",x"72",x"4a",x"70"),
   444 => (x"87",x"c5",x"c0",x"05"),
   445 => (x"c2",x"c0",x"4a",x"c1"),
   446 => (x"27",x"4a",x"c0",x"87"),
   447 => (x"00",x"00",x"17",x"0c"),
   448 => (x"6e",x"79",x"72",x"49"),
   449 => (x"a9",x"b7",x"74",x"49"),
   450 => (x"87",x"ed",x"c0",x"03"),
   451 => (x"92",x"c5",x"4a",x"6e"),
   452 => (x"88",x"74",x"48",x"72"),
   453 => (x"cc",x"58",x"a6",x"d0"),
   454 => (x"1e",x"72",x"4a",x"a6"),
   455 => (x"66",x"c8",x"1e",x"74"),
   456 => (x"03",x"17",x"27",x"1e"),
   457 => (x"cc",x"0f",x"00",x"00"),
   458 => (x"c1",x"48",x"6e",x"86"),
   459 => (x"58",x"a6",x"c4",x"80"),
   460 => (x"b7",x"74",x"49",x"6e"),
   461 => (x"d3",x"ff",x"04",x"a9"),
   462 => (x"1e",x"66",x"cc",x"87"),
   463 => (x"27",x"1e",x"66",x"c4"),
   464 => (x"00",x"00",x"17",x"e0"),
   465 => (x"17",x"18",x"27",x"1e"),
   466 => (x"27",x"1e",x"00",x"00"),
   467 => (x"00",x"00",x"03",x"2d"),
   468 => (x"27",x"86",x"d0",x"0f"),
   469 => (x"00",x"00",x"17",x"00"),
   470 => (x"56",x"27",x"1e",x"bf"),
   471 => (x"0f",x"00",x"00",x"0d"),
   472 => (x"a6",x"c4",x"86",x"c4"),
   473 => (x"51",x"c1",x"c1",x"49"),
   474 => (x"00",x"17",x"11",x"27"),
   475 => (x"4a",x"bf",x"97",x"00"),
   476 => (x"c0",x"c0",x"c0",x"c1"),
   477 => (x"c0",x"c4",x"92",x"c0"),
   478 => (x"c1",x"4a",x"92",x"b7"),
   479 => (x"04",x"aa",x"b7",x"c1"),
   480 => (x"c1",x"87",x"e6",x"c2"),
   481 => (x"c8",x"97",x"1e",x"c3"),
   482 => (x"c0",x"c1",x"4a",x"66"),
   483 => (x"92",x"c0",x"c0",x"c0"),
   484 => (x"92",x"b7",x"c0",x"c4"),
   485 => (x"27",x"1e",x"72",x"4a"),
   486 => (x"00",x"00",x"03",x"ba"),
   487 => (x"70",x"86",x"c8",x"0f"),
   488 => (x"49",x"66",x"c8",x"4a"),
   489 => (x"05",x"a9",x"b7",x"72"),
   490 => (x"c8",x"87",x"cb",x"c1"),
   491 => (x"1e",x"72",x"4a",x"a6"),
   492 => (x"a0",x"27",x"1e",x"c0"),
   493 => (x"0f",x"00",x"00",x"02"),
   494 => (x"88",x"27",x"86",x"c8"),
   495 => (x"49",x"00",x"00",x"3f"),
   496 => (x"00",x"0f",x"44",x"27"),
   497 => (x"1e",x"72",x"48",x"00"),
   498 => (x"81",x"c4",x"79",x"20"),
   499 => (x"81",x"c4",x"79",x"20"),
   500 => (x"81",x"c4",x"79",x"20"),
   501 => (x"81",x"c4",x"79",x"20"),
   502 => (x"81",x"c4",x"79",x"20"),
   503 => (x"81",x"c4",x"79",x"20"),
   504 => (x"81",x"c4",x"79",x"20"),
   505 => (x"51",x"10",x"51",x"10"),
   506 => (x"4a",x"26",x"51",x"10"),
   507 => (x"08",x"27",x"4c",x"75"),
   508 => (x"49",x"00",x"00",x"17"),
   509 => (x"c4",x"97",x"79",x"75"),
   510 => (x"80",x"c1",x"48",x"66"),
   511 => (x"50",x"08",x"a6",x"c4"),
   512 => (x"4b",x"66",x"c4",x"97"),
   513 => (x"c0",x"c0",x"c0",x"c1"),
   514 => (x"c0",x"c4",x"93",x"c0"),
   515 => (x"27",x"4b",x"93",x"b7"),
   516 => (x"00",x"00",x"17",x"11"),
   517 => (x"c1",x"4a",x"bf",x"97"),
   518 => (x"c0",x"c0",x"c0",x"c0"),
   519 => (x"b7",x"c0",x"c4",x"92"),
   520 => (x"b7",x"72",x"4a",x"92"),
   521 => (x"da",x"fd",x"06",x"ab"),
   522 => (x"74",x"94",x"6e",x"87"),
   523 => (x"d0",x"1e",x"72",x"49"),
   524 => (x"db",x"27",x"4a",x"66"),
   525 => (x"0f",x"00",x"00",x"04"),
   526 => (x"48",x"70",x"4a",x"26"),
   527 => (x"74",x"58",x"a6",x"c4"),
   528 => (x"8a",x"66",x"cc",x"4a"),
   529 => (x"4c",x"72",x"92",x"c7"),
   530 => (x"4a",x"76",x"8c",x"6e"),
   531 => (x"f9",x"27",x"1e",x"72"),
   532 => (x"0f",x"00",x"00",x"0d"),
   533 => (x"85",x"c1",x"86",x"c4"),
   534 => (x"00",x"16",x"88",x"27"),
   535 => (x"ad",x"b7",x"bf",x"00"),
   536 => (x"87",x"eb",x"f8",x"06"),
   537 => (x"00",x"05",x"32",x"27"),
   538 => (x"f8",x"27",x"0f",x"00"),
   539 => (x"58",x"00",x"00",x"3e"),
   540 => (x"00",x"10",x"fd",x"27"),
   541 => (x"52",x"27",x"1e",x"00"),
   542 => (x"0f",x"00",x"00",x"01"),
   543 => (x"0d",x"27",x"86",x"c4"),
   544 => (x"1e",x"00",x"00",x"11"),
   545 => (x"00",x"01",x"52",x"27"),
   546 => (x"86",x"c4",x"0f",x"00"),
   547 => (x"00",x"11",x"0f",x"27"),
   548 => (x"52",x"27",x"1e",x"00"),
   549 => (x"0f",x"00",x"00",x"01"),
   550 => (x"45",x"27",x"86",x"c4"),
   551 => (x"1e",x"00",x"00",x"11"),
   552 => (x"00",x"01",x"52",x"27"),
   553 => (x"86",x"c4",x"0f",x"00"),
   554 => (x"00",x"17",x"08",x"27"),
   555 => (x"27",x"1e",x"bf",x"00"),
   556 => (x"00",x"00",x"11",x"47"),
   557 => (x"01",x"52",x"27",x"1e"),
   558 => (x"c8",x"0f",x"00",x"00"),
   559 => (x"27",x"1e",x"c5",x"86"),
   560 => (x"00",x"00",x"11",x"60"),
   561 => (x"01",x"52",x"27",x"1e"),
   562 => (x"c8",x"0f",x"00",x"00"),
   563 => (x"17",x"0c",x"27",x"86"),
   564 => (x"1e",x"bf",x"00",x"00"),
   565 => (x"00",x"11",x"79",x"27"),
   566 => (x"52",x"27",x"1e",x"00"),
   567 => (x"0f",x"00",x"00",x"01"),
   568 => (x"1e",x"c1",x"86",x"c8"),
   569 => (x"00",x"11",x"92",x"27"),
   570 => (x"52",x"27",x"1e",x"00"),
   571 => (x"0f",x"00",x"00",x"01"),
   572 => (x"10",x"27",x"86",x"c8"),
   573 => (x"97",x"00",x"00",x"17"),
   574 => (x"c0",x"c1",x"4a",x"bf"),
   575 => (x"92",x"c0",x"c0",x"c0"),
   576 => (x"92",x"b7",x"c0",x"c4"),
   577 => (x"27",x"1e",x"72",x"4a"),
   578 => (x"00",x"00",x"11",x"ab"),
   579 => (x"01",x"52",x"27",x"1e"),
   580 => (x"c8",x"0f",x"00",x"00"),
   581 => (x"1e",x"c1",x"c1",x"86"),
   582 => (x"00",x"11",x"c4",x"27"),
   583 => (x"52",x"27",x"1e",x"00"),
   584 => (x"0f",x"00",x"00",x"01"),
   585 => (x"11",x"27",x"86",x"c8"),
   586 => (x"97",x"00",x"00",x"17"),
   587 => (x"c0",x"c1",x"4a",x"bf"),
   588 => (x"92",x"c0",x"c0",x"c0"),
   589 => (x"92",x"b7",x"c0",x"c4"),
   590 => (x"27",x"1e",x"72",x"4a"),
   591 => (x"00",x"00",x"11",x"dd"),
   592 => (x"01",x"52",x"27",x"1e"),
   593 => (x"c8",x"0f",x"00",x"00"),
   594 => (x"1e",x"c2",x"c1",x"86"),
   595 => (x"00",x"11",x"f6",x"27"),
   596 => (x"52",x"27",x"1e",x"00"),
   597 => (x"0f",x"00",x"00",x"01"),
   598 => (x"38",x"27",x"86",x"c8"),
   599 => (x"bf",x"00",x"00",x"17"),
   600 => (x"12",x"0f",x"27",x"1e"),
   601 => (x"27",x"1e",x"00",x"00"),
   602 => (x"00",x"00",x"01",x"52"),
   603 => (x"c7",x"86",x"c8",x"0f"),
   604 => (x"12",x"28",x"27",x"1e"),
   605 => (x"27",x"1e",x"00",x"00"),
   606 => (x"00",x"00",x"01",x"52"),
   607 => (x"27",x"86",x"c8",x"0f"),
   608 => (x"00",x"00",x"1e",x"3c"),
   609 => (x"41",x"27",x"1e",x"bf"),
   610 => (x"1e",x"00",x"00",x"12"),
   611 => (x"00",x"01",x"52",x"27"),
   612 => (x"86",x"c8",x"0f",x"00"),
   613 => (x"00",x"12",x"5a",x"27"),
   614 => (x"52",x"27",x"1e",x"00"),
   615 => (x"0f",x"00",x"00",x"01"),
   616 => (x"84",x"27",x"86",x"c4"),
   617 => (x"1e",x"00",x"00",x"12"),
   618 => (x"00",x"01",x"52",x"27"),
   619 => (x"86",x"c4",x"0f",x"00"),
   620 => (x"00",x"17",x"00",x"27"),
   621 => (x"1e",x"bf",x"bf",x"00"),
   622 => (x"00",x"12",x"90",x"27"),
   623 => (x"52",x"27",x"1e",x"00"),
   624 => (x"0f",x"00",x"00",x"01"),
   625 => (x"a9",x"27",x"86",x"c8"),
   626 => (x"1e",x"00",x"00",x"12"),
   627 => (x"00",x"01",x"52",x"27"),
   628 => (x"86",x"c4",x"0f",x"00"),
   629 => (x"00",x"17",x"00",x"27"),
   630 => (x"c4",x"4a",x"bf",x"00"),
   631 => (x"27",x"1e",x"6a",x"82"),
   632 => (x"00",x"00",x"12",x"da"),
   633 => (x"01",x"52",x"27",x"1e"),
   634 => (x"c8",x"0f",x"00",x"00"),
   635 => (x"27",x"1e",x"c0",x"86"),
   636 => (x"00",x"00",x"12",x"f3"),
   637 => (x"01",x"52",x"27",x"1e"),
   638 => (x"c8",x"0f",x"00",x"00"),
   639 => (x"17",x"00",x"27",x"86"),
   640 => (x"4a",x"bf",x"00",x"00"),
   641 => (x"1e",x"6a",x"82",x"c8"),
   642 => (x"00",x"13",x"0c",x"27"),
   643 => (x"52",x"27",x"1e",x"00"),
   644 => (x"0f",x"00",x"00",x"01"),
   645 => (x"1e",x"c2",x"86",x"c8"),
   646 => (x"00",x"13",x"25",x"27"),
   647 => (x"52",x"27",x"1e",x"00"),
   648 => (x"0f",x"00",x"00",x"01"),
   649 => (x"00",x"27",x"86",x"c8"),
   650 => (x"bf",x"00",x"00",x"17"),
   651 => (x"6a",x"82",x"cc",x"4a"),
   652 => (x"13",x"3e",x"27",x"1e"),
   653 => (x"27",x"1e",x"00",x"00"),
   654 => (x"00",x"00",x"01",x"52"),
   655 => (x"d1",x"86",x"c8",x"0f"),
   656 => (x"13",x"57",x"27",x"1e"),
   657 => (x"27",x"1e",x"00",x"00"),
   658 => (x"00",x"00",x"01",x"52"),
   659 => (x"27",x"86",x"c8",x"0f"),
   660 => (x"00",x"00",x"17",x"00"),
   661 => (x"82",x"d0",x"4a",x"bf"),
   662 => (x"70",x"27",x"1e",x"72"),
   663 => (x"1e",x"00",x"00",x"13"),
   664 => (x"00",x"01",x"52",x"27"),
   665 => (x"86",x"c8",x"0f",x"00"),
   666 => (x"00",x"13",x"89",x"27"),
   667 => (x"52",x"27",x"1e",x"00"),
   668 => (x"0f",x"00",x"00",x"01"),
   669 => (x"be",x"27",x"86",x"c4"),
   670 => (x"1e",x"00",x"00",x"13"),
   671 => (x"00",x"01",x"52",x"27"),
   672 => (x"86",x"c4",x"0f",x"00"),
   673 => (x"00",x"17",x"04",x"27"),
   674 => (x"1e",x"bf",x"bf",x"00"),
   675 => (x"00",x"13",x"cf",x"27"),
   676 => (x"52",x"27",x"1e",x"00"),
   677 => (x"0f",x"00",x"00",x"01"),
   678 => (x"e8",x"27",x"86",x"c8"),
   679 => (x"1e",x"00",x"00",x"13"),
   680 => (x"00",x"01",x"52",x"27"),
   681 => (x"86",x"c4",x"0f",x"00"),
   682 => (x"00",x"17",x"04",x"27"),
   683 => (x"c4",x"4a",x"bf",x"00"),
   684 => (x"27",x"1e",x"6a",x"82"),
   685 => (x"00",x"00",x"14",x"28"),
   686 => (x"01",x"52",x"27",x"1e"),
   687 => (x"c8",x"0f",x"00",x"00"),
   688 => (x"27",x"1e",x"c0",x"86"),
   689 => (x"00",x"00",x"14",x"41"),
   690 => (x"01",x"52",x"27",x"1e"),
   691 => (x"c8",x"0f",x"00",x"00"),
   692 => (x"17",x"04",x"27",x"86"),
   693 => (x"4a",x"bf",x"00",x"00"),
   694 => (x"1e",x"6a",x"82",x"c8"),
   695 => (x"00",x"14",x"5a",x"27"),
   696 => (x"52",x"27",x"1e",x"00"),
   697 => (x"0f",x"00",x"00",x"01"),
   698 => (x"1e",x"c1",x"86",x"c8"),
   699 => (x"00",x"14",x"73",x"27"),
   700 => (x"52",x"27",x"1e",x"00"),
   701 => (x"0f",x"00",x"00",x"01"),
   702 => (x"04",x"27",x"86",x"c8"),
   703 => (x"bf",x"00",x"00",x"17"),
   704 => (x"6a",x"82",x"cc",x"4a"),
   705 => (x"14",x"8c",x"27",x"1e"),
   706 => (x"27",x"1e",x"00",x"00"),
   707 => (x"00",x"00",x"01",x"52"),
   708 => (x"d2",x"86",x"c8",x"0f"),
   709 => (x"14",x"a5",x"27",x"1e"),
   710 => (x"27",x"1e",x"00",x"00"),
   711 => (x"00",x"00",x"01",x"52"),
   712 => (x"27",x"86",x"c8",x"0f"),
   713 => (x"00",x"00",x"17",x"04"),
   714 => (x"82",x"d0",x"4a",x"bf"),
   715 => (x"be",x"27",x"1e",x"72"),
   716 => (x"1e",x"00",x"00",x"14"),
   717 => (x"00",x"01",x"52",x"27"),
   718 => (x"86",x"c8",x"0f",x"00"),
   719 => (x"00",x"14",x"d7",x"27"),
   720 => (x"52",x"27",x"1e",x"00"),
   721 => (x"0f",x"00",x"00",x"01"),
   722 => (x"1e",x"6e",x"86",x"c4"),
   723 => (x"00",x"15",x"0c",x"27"),
   724 => (x"52",x"27",x"1e",x"00"),
   725 => (x"0f",x"00",x"00",x"01"),
   726 => (x"1e",x"c5",x"86",x"c8"),
   727 => (x"00",x"15",x"25",x"27"),
   728 => (x"52",x"27",x"1e",x"00"),
   729 => (x"0f",x"00",x"00",x"01"),
   730 => (x"1e",x"74",x"86",x"c8"),
   731 => (x"00",x"15",x"3e",x"27"),
   732 => (x"52",x"27",x"1e",x"00"),
   733 => (x"0f",x"00",x"00",x"01"),
   734 => (x"1e",x"cd",x"86",x"c8"),
   735 => (x"00",x"15",x"57",x"27"),
   736 => (x"52",x"27",x"1e",x"00"),
   737 => (x"0f",x"00",x"00",x"01"),
   738 => (x"66",x"cc",x"86",x"c8"),
   739 => (x"15",x"70",x"27",x"1e"),
   740 => (x"27",x"1e",x"00",x"00"),
   741 => (x"00",x"00",x"01",x"52"),
   742 => (x"c7",x"86",x"c8",x"0f"),
   743 => (x"15",x"89",x"27",x"1e"),
   744 => (x"27",x"1e",x"00",x"00"),
   745 => (x"00",x"00",x"01",x"52"),
   746 => (x"c8",x"86",x"c8",x"0f"),
   747 => (x"a2",x"27",x"1e",x"66"),
   748 => (x"1e",x"00",x"00",x"15"),
   749 => (x"00",x"01",x"52",x"27"),
   750 => (x"86",x"c8",x"0f",x"00"),
   751 => (x"bb",x"27",x"1e",x"c1"),
   752 => (x"1e",x"00",x"00",x"15"),
   753 => (x"00",x"01",x"52",x"27"),
   754 => (x"86",x"c8",x"0f",x"00"),
   755 => (x"00",x"3f",x"68",x"27"),
   756 => (x"d4",x"27",x"1e",x"00"),
   757 => (x"1e",x"00",x"00",x"15"),
   758 => (x"00",x"01",x"52",x"27"),
   759 => (x"86",x"c8",x"0f",x"00"),
   760 => (x"00",x"15",x"ed",x"27"),
   761 => (x"52",x"27",x"1e",x"00"),
   762 => (x"0f",x"00",x"00",x"01"),
   763 => (x"88",x"27",x"86",x"c4"),
   764 => (x"1e",x"00",x"00",x"3f"),
   765 => (x"00",x"16",x"22",x"27"),
   766 => (x"52",x"27",x"1e",x"00"),
   767 => (x"0f",x"00",x"00",x"01"),
   768 => (x"3b",x"27",x"86",x"c8"),
   769 => (x"1e",x"00",x"00",x"16"),
   770 => (x"00",x"01",x"52",x"27"),
   771 => (x"86",x"c4",x"0f",x"00"),
   772 => (x"00",x"16",x"70",x"27"),
   773 => (x"52",x"27",x"1e",x"00"),
   774 => (x"0f",x"00",x"00",x"01"),
   775 => (x"f4",x"27",x"86",x"c4"),
   776 => (x"bf",x"00",x"00",x"3e"),
   777 => (x"3e",x"f0",x"27",x"4a"),
   778 => (x"8a",x"bf",x"00",x"00"),
   779 => (x"00",x"3e",x"f8",x"27"),
   780 => (x"79",x"72",x"49",x"00"),
   781 => (x"72",x"27",x"1e",x"72"),
   782 => (x"1e",x"00",x"00",x"16"),
   783 => (x"00",x"01",x"52",x"27"),
   784 => (x"86",x"c8",x"0f",x"00"),
   785 => (x"00",x"3e",x"f8",x"27"),
   786 => (x"c1",x"49",x"bf",x"00"),
   787 => (x"03",x"a9",x"b7",x"f8"),
   788 => (x"27",x"87",x"ea",x"c0"),
   789 => (x"00",x"00",x"0f",x"82"),
   790 => (x"01",x"52",x"27",x"1e"),
   791 => (x"c4",x"0f",x"00",x"00"),
   792 => (x"0f",x"b8",x"27",x"86"),
   793 => (x"27",x"1e",x"00",x"00"),
   794 => (x"00",x"00",x"01",x"52"),
   795 => (x"27",x"86",x"c4",x"0f"),
   796 => (x"00",x"00",x"0f",x"d8"),
   797 => (x"01",x"52",x"27",x"1e"),
   798 => (x"c4",x"0f",x"00",x"00"),
   799 => (x"3e",x"f8",x"27",x"86"),
   800 => (x"4a",x"bf",x"00",x"00"),
   801 => (x"e8",x"cf",x"4b",x"72"),
   802 => (x"72",x"49",x"73",x"93"),
   803 => (x"16",x"88",x"27",x"1e"),
   804 => (x"4a",x"bf",x"00",x"00"),
   805 => (x"00",x"04",x"db",x"27"),
   806 => (x"4a",x"26",x"0f",x"00"),
   807 => (x"00",x"27",x"48",x"70"),
   808 => (x"58",x"00",x"00",x"3f"),
   809 => (x"00",x"16",x"88",x"27"),
   810 => (x"73",x"4b",x"bf",x"00"),
   811 => (x"94",x"e8",x"cf",x"4c"),
   812 => (x"1e",x"72",x"49",x"74"),
   813 => (x"db",x"27",x"4a",x"72"),
   814 => (x"0f",x"00",x"00",x"04"),
   815 => (x"48",x"70",x"4a",x"26"),
   816 => (x"00",x"3f",x"04",x"27"),
   817 => (x"f9",x"c8",x"58",x"00"),
   818 => (x"72",x"49",x"73",x"93"),
   819 => (x"27",x"4a",x"72",x"1e"),
   820 => (x"00",x"00",x"04",x"db"),
   821 => (x"70",x"4a",x"26",x"0f"),
   822 => (x"3f",x"08",x"27",x"48"),
   823 => (x"27",x"58",x"00",x"00"),
   824 => (x"00",x"00",x"0f",x"da"),
   825 => (x"01",x"52",x"27",x"1e"),
   826 => (x"c4",x"0f",x"00",x"00"),
   827 => (x"3e",x"fc",x"27",x"86"),
   828 => (x"1e",x"bf",x"00",x"00"),
   829 => (x"00",x"10",x"07",x"27"),
   830 => (x"52",x"27",x"1e",x"00"),
   831 => (x"0f",x"00",x"00",x"01"),
   832 => (x"0c",x"27",x"86",x"c8"),
   833 => (x"1e",x"00",x"00",x"10"),
   834 => (x"00",x"01",x"52",x"27"),
   835 => (x"86",x"c4",x"0f",x"00"),
   836 => (x"00",x"3f",x"00",x"27"),
   837 => (x"27",x"1e",x"bf",x"00"),
   838 => (x"00",x"00",x"10",x"39"),
   839 => (x"01",x"52",x"27",x"1e"),
   840 => (x"c8",x"0f",x"00",x"00"),
   841 => (x"3f",x"04",x"27",x"86"),
   842 => (x"1e",x"bf",x"00",x"00"),
   843 => (x"00",x"10",x"3e",x"27"),
   844 => (x"52",x"27",x"1e",x"00"),
   845 => (x"0f",x"00",x"00",x"01"),
   846 => (x"5c",x"27",x"86",x"c8"),
   847 => (x"1e",x"00",x"00",x"10"),
   848 => (x"00",x"01",x"52",x"27"),
   849 => (x"86",x"c4",x"0f",x"00"),
   850 => (x"86",x"d0",x"48",x"c0"),
   851 => (x"4c",x"26",x"4d",x"26"),
   852 => (x"4a",x"26",x"4b",x"26"),
   853 => (x"5e",x"0e",x"4f",x"26"),
   854 => (x"5d",x"5c",x"5b",x"5a"),
   855 => (x"bf",x"a6",x"d4",x"0e"),
   856 => (x"4d",x"72",x"4a",x"bf"),
   857 => (x"00",x"17",x"00",x"27"),
   858 => (x"72",x"48",x"bf",x"00"),
   859 => (x"a2",x"f0",x"c0",x"1e"),
   860 => (x"c4",x"7a",x"20",x"49"),
   861 => (x"05",x"a9",x"72",x"82"),
   862 => (x"4a",x"26",x"87",x"f7"),
   863 => (x"cc",x"4c",x"66",x"d4"),
   864 => (x"72",x"7c",x"c5",x"84"),
   865 => (x"6c",x"83",x"cc",x"4b"),
   866 => (x"bf",x"a6",x"d4",x"7b"),
   867 => (x"1e",x"72",x"7a",x"bf"),
   868 => (x"00",x"0e",x"45",x"27"),
   869 => (x"86",x"c4",x"0f",x"00"),
   870 => (x"9a",x"6a",x"82",x"c4"),
   871 => (x"87",x"f4",x"c0",x"05"),
   872 => (x"83",x"c8",x"4b",x"75"),
   873 => (x"82",x"cc",x"4a",x"75"),
   874 => (x"1e",x"73",x"7a",x"c6"),
   875 => (x"c8",x"4b",x"66",x"d8"),
   876 => (x"27",x"1e",x"6b",x"83"),
   877 => (x"00",x"00",x"02",x"a0"),
   878 => (x"27",x"86",x"c8",x"0f"),
   879 => (x"00",x"00",x"17",x"00"),
   880 => (x"72",x"7d",x"bf",x"bf"),
   881 => (x"6a",x"1e",x"ca",x"1e"),
   882 => (x"03",x"17",x"27",x"1e"),
   883 => (x"cc",x"0f",x"00",x"00"),
   884 => (x"87",x"db",x"c0",x"86"),
   885 => (x"bf",x"bf",x"a6",x"d4"),
   886 => (x"bf",x"a6",x"d4",x"4a"),
   887 => (x"1e",x"72",x"48",x"49"),
   888 => (x"4a",x"a1",x"f0",x"c0"),
   889 => (x"81",x"c4",x"79",x"20"),
   890 => (x"f7",x"05",x"aa",x"71"),
   891 => (x"26",x"4a",x"26",x"87"),
   892 => (x"26",x"4c",x"26",x"4d"),
   893 => (x"26",x"4a",x"26",x"4b"),
   894 => (x"5a",x"5e",x"0e",x"4f"),
   895 => (x"0e",x"5d",x"5c",x"5b"),
   896 => (x"d8",x"4d",x"6e",x"1e"),
   897 => (x"4b",x"6c",x"4c",x"66"),
   898 => (x"10",x"27",x"83",x"ca"),
   899 => (x"97",x"00",x"00",x"17"),
   900 => (x"c0",x"c1",x"4a",x"bf"),
   901 => (x"92",x"c0",x"c0",x"c0"),
   902 => (x"92",x"b7",x"c0",x"c4"),
   903 => (x"b7",x"c1",x"c1",x"4a"),
   904 => (x"cf",x"c0",x"05",x"aa"),
   905 => (x"73",x"8b",x"c1",x"87"),
   906 => (x"17",x"08",x"27",x"48"),
   907 => (x"88",x"bf",x"00",x"00"),
   908 => (x"4d",x"c0",x"7c",x"70"),
   909 => (x"ff",x"05",x"9d",x"75"),
   910 => (x"26",x"26",x"87",x"d0"),
   911 => (x"26",x"4c",x"26",x"4d"),
   912 => (x"26",x"4a",x"26",x"4b"),
   913 => (x"1e",x"72",x"1e",x"4f"),
   914 => (x"00",x"17",x"00",x"27"),
   915 => (x"c0",x"02",x"bf",x"00"),
   916 => (x"a6",x"c8",x"87",x"cc"),
   917 => (x"00",x"27",x"49",x"bf"),
   918 => (x"bf",x"00",x"00",x"17"),
   919 => (x"00",x"27",x"79",x"bf"),
   920 => (x"bf",x"00",x"00",x"17"),
   921 => (x"72",x"82",x"cc",x"4a"),
   922 => (x"17",x"08",x"27",x"1e"),
   923 => (x"1e",x"bf",x"00",x"00"),
   924 => (x"17",x"27",x"1e",x"ca"),
   925 => (x"0f",x"00",x"00",x"03"),
   926 => (x"4a",x"26",x"86",x"cc"),
   927 => (x"72",x"1e",x"4f",x"26"),
   928 => (x"17",x"10",x"27",x"1e"),
   929 => (x"bf",x"97",x"00",x"00"),
   930 => (x"c0",x"c0",x"c1",x"4a"),
   931 => (x"c4",x"92",x"c0",x"c0"),
   932 => (x"4a",x"92",x"b7",x"c0"),
   933 => (x"aa",x"b7",x"c1",x"c1"),
   934 => (x"87",x"c5",x"c0",x"02"),
   935 => (x"c2",x"c0",x"4a",x"c0"),
   936 => (x"27",x"4a",x"c1",x"87"),
   937 => (x"00",x"00",x"17",x"0c"),
   938 => (x"b0",x"72",x"48",x"bf"),
   939 => (x"00",x"17",x"10",x"27"),
   940 => (x"11",x"27",x"58",x"00"),
   941 => (x"49",x"00",x"00",x"17"),
   942 => (x"26",x"51",x"c2",x"c1"),
   943 => (x"1e",x"4f",x"26",x"4a"),
   944 => (x"00",x"17",x"10",x"27"),
   945 => (x"c1",x"c1",x"49",x"00"),
   946 => (x"17",x"0c",x"27",x"51"),
   947 => (x"c0",x"49",x"00",x"00"),
   948 => (x"00",x"4f",x"26",x"79"),
   949 => (x"33",x"32",x"31",x"30"),
   950 => (x"37",x"36",x"35",x"34"),
   951 => (x"42",x"41",x"39",x"38"),
   952 => (x"46",x"45",x"44",x"43"),
   953 => (x"6f",x"72",x"50",x"00"),
   954 => (x"6d",x"61",x"72",x"67"),
   955 => (x"6d",x"6f",x"63",x"20"),
   956 => (x"65",x"6c",x"69",x"70"),
   957 => (x"69",x"77",x"20",x"64"),
   958 => (x"27",x"20",x"68",x"74"),
   959 => (x"69",x"67",x"65",x"72"),
   960 => (x"72",x"65",x"74",x"73"),
   961 => (x"74",x"61",x"20",x"27"),
   962 => (x"62",x"69",x"72",x"74"),
   963 => (x"0a",x"65",x"74",x"75"),
   964 => (x"50",x"00",x"0a",x"00"),
   965 => (x"72",x"67",x"6f",x"72"),
   966 => (x"63",x"20",x"6d",x"61"),
   967 => (x"69",x"70",x"6d",x"6f"),
   968 => (x"20",x"64",x"65",x"6c"),
   969 => (x"68",x"74",x"69",x"77"),
   970 => (x"20",x"74",x"75",x"6f"),
   971 => (x"67",x"65",x"72",x"27"),
   972 => (x"65",x"74",x"73",x"69"),
   973 => (x"61",x"20",x"27",x"72"),
   974 => (x"69",x"72",x"74",x"74"),
   975 => (x"65",x"74",x"75",x"62"),
   976 => (x"00",x"0a",x"00",x"0a"),
   977 => (x"59",x"52",x"48",x"44"),
   978 => (x"4e",x"4f",x"54",x"53"),
   979 => (x"52",x"50",x"20",x"45"),
   980 => (x"41",x"52",x"47",x"4f"),
   981 => (x"33",x"20",x"2c",x"4d"),
   982 => (x"20",x"44",x"52",x"27"),
   983 => (x"49",x"52",x"54",x"53"),
   984 => (x"44",x"00",x"47",x"4e"),
   985 => (x"53",x"59",x"52",x"48"),
   986 => (x"45",x"4e",x"4f",x"54"),
   987 => (x"4f",x"52",x"50",x"20"),
   988 => (x"4d",x"41",x"52",x"47"),
   989 => (x"27",x"32",x"20",x"2c"),
   990 => (x"53",x"20",x"44",x"4e"),
   991 => (x"4e",x"49",x"52",x"54"),
   992 => (x"65",x"4d",x"00",x"47"),
   993 => (x"72",x"75",x"73",x"61"),
   994 => (x"74",x"20",x"64",x"65"),
   995 => (x"20",x"65",x"6d",x"69"),
   996 => (x"20",x"6f",x"6f",x"74"),
   997 => (x"6c",x"61",x"6d",x"73"),
   998 => (x"6f",x"74",x"20",x"6c"),
   999 => (x"74",x"62",x"6f",x"20"),
  1000 => (x"20",x"6e",x"69",x"61"),
  1001 => (x"6e",x"61",x"65",x"6d"),
  1002 => (x"66",x"67",x"6e",x"69"),
  1003 => (x"72",x"20",x"6c",x"75"),
  1004 => (x"6c",x"75",x"73",x"65"),
  1005 => (x"00",x"0a",x"73",x"74"),
  1006 => (x"61",x"65",x"6c",x"50"),
  1007 => (x"69",x"20",x"65",x"73"),
  1008 => (x"65",x"72",x"63",x"6e"),
  1009 => (x"20",x"65",x"73",x"61"),
  1010 => (x"62",x"6d",x"75",x"6e"),
  1011 => (x"6f",x"20",x"72",x"65"),
  1012 => (x"75",x"72",x"20",x"66"),
  1013 => (x"00",x"0a",x"73",x"6e"),
  1014 => (x"69",x"4d",x"00",x"0a"),
  1015 => (x"73",x"6f",x"72",x"63"),
  1016 => (x"6e",x"6f",x"63",x"65"),
  1017 => (x"66",x"20",x"73",x"64"),
  1018 => (x"6f",x"20",x"72",x"6f"),
  1019 => (x"72",x"20",x"65",x"6e"),
  1020 => (x"74",x"20",x"6e",x"75"),
  1021 => (x"75",x"6f",x"72",x"68"),
  1022 => (x"44",x"20",x"68",x"67"),
  1023 => (x"73",x"79",x"72",x"68"),
  1024 => (x"65",x"6e",x"6f",x"74"),
  1025 => (x"25",x"00",x"20",x"3a"),
  1026 => (x"00",x"0a",x"20",x"64"),
  1027 => (x"79",x"72",x"68",x"44"),
  1028 => (x"6e",x"6f",x"74",x"73"),
  1029 => (x"70",x"20",x"73",x"65"),
  1030 => (x"53",x"20",x"72",x"65"),
  1031 => (x"6e",x"6f",x"63",x"65"),
  1032 => (x"20",x"20",x"3a",x"64"),
  1033 => (x"20",x"20",x"20",x"20"),
  1034 => (x"20",x"20",x"20",x"20"),
  1035 => (x"20",x"20",x"20",x"20"),
  1036 => (x"20",x"20",x"20",x"20"),
  1037 => (x"20",x"20",x"20",x"20"),
  1038 => (x"20",x"64",x"25",x"00"),
  1039 => (x"41",x"56",x"00",x"0a"),
  1040 => (x"49",x"4d",x"20",x"58"),
  1041 => (x"72",x"20",x"53",x"50"),
  1042 => (x"6e",x"69",x"74",x"61"),
  1043 => (x"20",x"2a",x"20",x"67"),
  1044 => (x"30",x"30",x"30",x"31"),
  1045 => (x"25",x"20",x"3d",x"20"),
  1046 => (x"00",x"0a",x"20",x"64"),
  1047 => (x"48",x"44",x"00",x"0a"),
  1048 => (x"54",x"53",x"59",x"52"),
  1049 => (x"20",x"45",x"4e",x"4f"),
  1050 => (x"47",x"4f",x"52",x"50"),
  1051 => (x"2c",x"4d",x"41",x"52"),
  1052 => (x"4d",x"4f",x"53",x"20"),
  1053 => (x"54",x"53",x"20",x"45"),
  1054 => (x"47",x"4e",x"49",x"52"),
  1055 => (x"52",x"48",x"44",x"00"),
  1056 => (x"4f",x"54",x"53",x"59"),
  1057 => (x"50",x"20",x"45",x"4e"),
  1058 => (x"52",x"47",x"4f",x"52"),
  1059 => (x"20",x"2c",x"4d",x"41"),
  1060 => (x"54",x"53",x"27",x"31"),
  1061 => (x"52",x"54",x"53",x"20"),
  1062 => (x"00",x"47",x"4e",x"49"),
  1063 => (x"68",x"44",x"00",x"0a"),
  1064 => (x"74",x"73",x"79",x"72"),
  1065 => (x"20",x"65",x"6e",x"6f"),
  1066 => (x"63",x"6e",x"65",x"42"),
  1067 => (x"72",x"61",x"6d",x"68"),
  1068 => (x"56",x"20",x"2c",x"6b"),
  1069 => (x"69",x"73",x"72",x"65"),
  1070 => (x"32",x"20",x"6e",x"6f"),
  1071 => (x"28",x"20",x"31",x"2e"),
  1072 => (x"67",x"6e",x"61",x"4c"),
  1073 => (x"65",x"67",x"61",x"75"),
  1074 => (x"29",x"43",x"20",x"3a"),
  1075 => (x"00",x"0a",x"00",x"0a"),
  1076 => (x"63",x"65",x"78",x"45"),
  1077 => (x"6f",x"69",x"74",x"75"),
  1078 => (x"74",x"73",x"20",x"6e"),
  1079 => (x"73",x"74",x"72",x"61"),
  1080 => (x"64",x"25",x"20",x"2c"),
  1081 => (x"6e",x"75",x"72",x"20"),
  1082 => (x"68",x"74",x"20",x"73"),
  1083 => (x"67",x"75",x"6f",x"72"),
  1084 => (x"68",x"44",x"20",x"68"),
  1085 => (x"74",x"73",x"79",x"72"),
  1086 => (x"0a",x"65",x"6e",x"6f"),
  1087 => (x"65",x"78",x"45",x"00"),
  1088 => (x"69",x"74",x"75",x"63"),
  1089 => (x"65",x"20",x"6e",x"6f"),
  1090 => (x"0a",x"73",x"64",x"6e"),
  1091 => (x"46",x"00",x"0a",x"00"),
  1092 => (x"6c",x"61",x"6e",x"69"),
  1093 => (x"6c",x"61",x"76",x"20"),
  1094 => (x"20",x"73",x"65",x"75"),
  1095 => (x"74",x"20",x"66",x"6f"),
  1096 => (x"76",x"20",x"65",x"68"),
  1097 => (x"61",x"69",x"72",x"61"),
  1098 => (x"73",x"65",x"6c",x"62"),
  1099 => (x"65",x"73",x"75",x"20"),
  1100 => (x"6e",x"69",x"20",x"64"),
  1101 => (x"65",x"68",x"74",x"20"),
  1102 => (x"6e",x"65",x"62",x"20"),
  1103 => (x"61",x"6d",x"68",x"63"),
  1104 => (x"0a",x"3a",x"6b",x"72"),
  1105 => (x"49",x"00",x"0a",x"00"),
  1106 => (x"47",x"5f",x"74",x"6e"),
  1107 => (x"3a",x"62",x"6f",x"6c"),
  1108 => (x"20",x"20",x"20",x"20"),
  1109 => (x"20",x"20",x"20",x"20"),
  1110 => (x"20",x"20",x"20",x"20"),
  1111 => (x"00",x"0a",x"64",x"25"),
  1112 => (x"20",x"20",x"20",x"20"),
  1113 => (x"20",x"20",x"20",x"20"),
  1114 => (x"75",x"6f",x"68",x"73"),
  1115 => (x"62",x"20",x"64",x"6c"),
  1116 => (x"20",x"20",x"3a",x"65"),
  1117 => (x"0a",x"64",x"25",x"20"),
  1118 => (x"6f",x"6f",x"42",x"00"),
  1119 => (x"6c",x"47",x"5f",x"6c"),
  1120 => (x"20",x"3a",x"62",x"6f"),
  1121 => (x"20",x"20",x"20",x"20"),
  1122 => (x"20",x"20",x"20",x"20"),
  1123 => (x"64",x"25",x"20",x"20"),
  1124 => (x"20",x"20",x"00",x"0a"),
  1125 => (x"20",x"20",x"20",x"20"),
  1126 => (x"68",x"73",x"20",x"20"),
  1127 => (x"64",x"6c",x"75",x"6f"),
  1128 => (x"3a",x"65",x"62",x"20"),
  1129 => (x"25",x"20",x"20",x"20"),
  1130 => (x"43",x"00",x"0a",x"64"),
  1131 => (x"5f",x"31",x"5f",x"68"),
  1132 => (x"62",x"6f",x"6c",x"47"),
  1133 => (x"20",x"20",x"20",x"3a"),
  1134 => (x"20",x"20",x"20",x"20"),
  1135 => (x"20",x"20",x"20",x"20"),
  1136 => (x"00",x"0a",x"63",x"25"),
  1137 => (x"20",x"20",x"20",x"20"),
  1138 => (x"20",x"20",x"20",x"20"),
  1139 => (x"75",x"6f",x"68",x"73"),
  1140 => (x"62",x"20",x"64",x"6c"),
  1141 => (x"20",x"20",x"3a",x"65"),
  1142 => (x"0a",x"63",x"25",x"20"),
  1143 => (x"5f",x"68",x"43",x"00"),
  1144 => (x"6c",x"47",x"5f",x"32"),
  1145 => (x"20",x"3a",x"62",x"6f"),
  1146 => (x"20",x"20",x"20",x"20"),
  1147 => (x"20",x"20",x"20",x"20"),
  1148 => (x"63",x"25",x"20",x"20"),
  1149 => (x"20",x"20",x"00",x"0a"),
  1150 => (x"20",x"20",x"20",x"20"),
  1151 => (x"68",x"73",x"20",x"20"),
  1152 => (x"64",x"6c",x"75",x"6f"),
  1153 => (x"3a",x"65",x"62",x"20"),
  1154 => (x"25",x"20",x"20",x"20"),
  1155 => (x"41",x"00",x"0a",x"63"),
  1156 => (x"31",x"5f",x"72",x"72"),
  1157 => (x"6f",x"6c",x"47",x"5f"),
  1158 => (x"5d",x"38",x"5b",x"62"),
  1159 => (x"20",x"20",x"20",x"3a"),
  1160 => (x"20",x"20",x"20",x"20"),
  1161 => (x"00",x"0a",x"64",x"25"),
  1162 => (x"20",x"20",x"20",x"20"),
  1163 => (x"20",x"20",x"20",x"20"),
  1164 => (x"75",x"6f",x"68",x"73"),
  1165 => (x"62",x"20",x"64",x"6c"),
  1166 => (x"20",x"20",x"3a",x"65"),
  1167 => (x"0a",x"64",x"25",x"20"),
  1168 => (x"72",x"72",x"41",x"00"),
  1169 => (x"47",x"5f",x"32",x"5f"),
  1170 => (x"5b",x"62",x"6f",x"6c"),
  1171 => (x"37",x"5b",x"5d",x"38"),
  1172 => (x"20",x"20",x"3a",x"5d"),
  1173 => (x"64",x"25",x"20",x"20"),
  1174 => (x"20",x"20",x"00",x"0a"),
  1175 => (x"20",x"20",x"20",x"20"),
  1176 => (x"68",x"73",x"20",x"20"),
  1177 => (x"64",x"6c",x"75",x"6f"),
  1178 => (x"3a",x"65",x"62",x"20"),
  1179 => (x"4e",x"20",x"20",x"20"),
  1180 => (x"65",x"62",x"6d",x"75"),
  1181 => (x"66",x"4f",x"5f",x"72"),
  1182 => (x"6e",x"75",x"52",x"5f"),
  1183 => (x"20",x"2b",x"20",x"73"),
  1184 => (x"00",x"0a",x"30",x"31"),
  1185 => (x"5f",x"72",x"74",x"50"),
  1186 => (x"62",x"6f",x"6c",x"47"),
  1187 => (x"00",x"0a",x"3e",x"2d"),
  1188 => (x"74",x"50",x"20",x"20"),
  1189 => (x"6f",x"43",x"5f",x"72"),
  1190 => (x"20",x"3a",x"70",x"6d"),
  1191 => (x"20",x"20",x"20",x"20"),
  1192 => (x"20",x"20",x"20",x"20"),
  1193 => (x"0a",x"64",x"25",x"20"),
  1194 => (x"20",x"20",x"20",x"00"),
  1195 => (x"20",x"20",x"20",x"20"),
  1196 => (x"6f",x"68",x"73",x"20"),
  1197 => (x"20",x"64",x"6c",x"75"),
  1198 => (x"20",x"3a",x"65",x"62"),
  1199 => (x"69",x"28",x"20",x"20"),
  1200 => (x"65",x"6c",x"70",x"6d"),
  1201 => (x"74",x"6e",x"65",x"6d"),
  1202 => (x"6f",x"69",x"74",x"61"),
  1203 => (x"65",x"64",x"2d",x"6e"),
  1204 => (x"64",x"6e",x"65",x"70"),
  1205 => (x"29",x"74",x"6e",x"65"),
  1206 => (x"20",x"20",x"00",x"0a"),
  1207 => (x"63",x"73",x"69",x"44"),
  1208 => (x"20",x"20",x"3a",x"72"),
  1209 => (x"20",x"20",x"20",x"20"),
  1210 => (x"20",x"20",x"20",x"20"),
  1211 => (x"25",x"20",x"20",x"20"),
  1212 => (x"20",x"00",x"0a",x"64"),
  1213 => (x"20",x"20",x"20",x"20"),
  1214 => (x"73",x"20",x"20",x"20"),
  1215 => (x"6c",x"75",x"6f",x"68"),
  1216 => (x"65",x"62",x"20",x"64"),
  1217 => (x"20",x"20",x"20",x"3a"),
  1218 => (x"00",x"0a",x"64",x"25"),
  1219 => (x"6e",x"45",x"20",x"20"),
  1220 => (x"43",x"5f",x"6d",x"75"),
  1221 => (x"3a",x"70",x"6d",x"6f"),
  1222 => (x"20",x"20",x"20",x"20"),
  1223 => (x"20",x"20",x"20",x"20"),
  1224 => (x"0a",x"64",x"25",x"20"),
  1225 => (x"20",x"20",x"20",x"00"),
  1226 => (x"20",x"20",x"20",x"20"),
  1227 => (x"6f",x"68",x"73",x"20"),
  1228 => (x"20",x"64",x"6c",x"75"),
  1229 => (x"20",x"3a",x"65",x"62"),
  1230 => (x"64",x"25",x"20",x"20"),
  1231 => (x"20",x"20",x"00",x"0a"),
  1232 => (x"5f",x"74",x"6e",x"49"),
  1233 => (x"70",x"6d",x"6f",x"43"),
  1234 => (x"20",x"20",x"20",x"3a"),
  1235 => (x"20",x"20",x"20",x"20"),
  1236 => (x"25",x"20",x"20",x"20"),
  1237 => (x"20",x"00",x"0a",x"64"),
  1238 => (x"20",x"20",x"20",x"20"),
  1239 => (x"73",x"20",x"20",x"20"),
  1240 => (x"6c",x"75",x"6f",x"68"),
  1241 => (x"65",x"62",x"20",x"64"),
  1242 => (x"20",x"20",x"20",x"3a"),
  1243 => (x"00",x"0a",x"64",x"25"),
  1244 => (x"74",x"53",x"20",x"20"),
  1245 => (x"6f",x"43",x"5f",x"72"),
  1246 => (x"20",x"3a",x"70",x"6d"),
  1247 => (x"20",x"20",x"20",x"20"),
  1248 => (x"20",x"20",x"20",x"20"),
  1249 => (x"0a",x"73",x"25",x"20"),
  1250 => (x"20",x"20",x"20",x"00"),
  1251 => (x"20",x"20",x"20",x"20"),
  1252 => (x"6f",x"68",x"73",x"20"),
  1253 => (x"20",x"64",x"6c",x"75"),
  1254 => (x"20",x"3a",x"65",x"62"),
  1255 => (x"48",x"44",x"20",x"20"),
  1256 => (x"54",x"53",x"59",x"52"),
  1257 => (x"20",x"45",x"4e",x"4f"),
  1258 => (x"47",x"4f",x"52",x"50"),
  1259 => (x"2c",x"4d",x"41",x"52"),
  1260 => (x"4d",x"4f",x"53",x"20"),
  1261 => (x"54",x"53",x"20",x"45"),
  1262 => (x"47",x"4e",x"49",x"52"),
  1263 => (x"65",x"4e",x"00",x"0a"),
  1264 => (x"50",x"5f",x"74",x"78"),
  1265 => (x"47",x"5f",x"72",x"74"),
  1266 => (x"2d",x"62",x"6f",x"6c"),
  1267 => (x"20",x"00",x"0a",x"3e"),
  1268 => (x"72",x"74",x"50",x"20"),
  1269 => (x"6d",x"6f",x"43",x"5f"),
  1270 => (x"20",x"20",x"3a",x"70"),
  1271 => (x"20",x"20",x"20",x"20"),
  1272 => (x"20",x"20",x"20",x"20"),
  1273 => (x"00",x"0a",x"64",x"25"),
  1274 => (x"20",x"20",x"20",x"20"),
  1275 => (x"20",x"20",x"20",x"20"),
  1276 => (x"75",x"6f",x"68",x"73"),
  1277 => (x"62",x"20",x"64",x"6c"),
  1278 => (x"20",x"20",x"3a",x"65"),
  1279 => (x"6d",x"69",x"28",x"20"),
  1280 => (x"6d",x"65",x"6c",x"70"),
  1281 => (x"61",x"74",x"6e",x"65"),
  1282 => (x"6e",x"6f",x"69",x"74"),
  1283 => (x"70",x"65",x"64",x"2d"),
  1284 => (x"65",x"64",x"6e",x"65"),
  1285 => (x"2c",x"29",x"74",x"6e"),
  1286 => (x"6d",x"61",x"73",x"20"),
  1287 => (x"73",x"61",x"20",x"65"),
  1288 => (x"6f",x"62",x"61",x"20"),
  1289 => (x"00",x"0a",x"65",x"76"),
  1290 => (x"69",x"44",x"20",x"20"),
  1291 => (x"3a",x"72",x"63",x"73"),
  1292 => (x"20",x"20",x"20",x"20"),
  1293 => (x"20",x"20",x"20",x"20"),
  1294 => (x"20",x"20",x"20",x"20"),
  1295 => (x"0a",x"64",x"25",x"20"),
  1296 => (x"20",x"20",x"20",x"00"),
  1297 => (x"20",x"20",x"20",x"20"),
  1298 => (x"6f",x"68",x"73",x"20"),
  1299 => (x"20",x"64",x"6c",x"75"),
  1300 => (x"20",x"3a",x"65",x"62"),
  1301 => (x"64",x"25",x"20",x"20"),
  1302 => (x"20",x"20",x"00",x"0a"),
  1303 => (x"6d",x"75",x"6e",x"45"),
  1304 => (x"6d",x"6f",x"43",x"5f"),
  1305 => (x"20",x"20",x"3a",x"70"),
  1306 => (x"20",x"20",x"20",x"20"),
  1307 => (x"25",x"20",x"20",x"20"),
  1308 => (x"20",x"00",x"0a",x"64"),
  1309 => (x"20",x"20",x"20",x"20"),
  1310 => (x"73",x"20",x"20",x"20"),
  1311 => (x"6c",x"75",x"6f",x"68"),
  1312 => (x"65",x"62",x"20",x"64"),
  1313 => (x"20",x"20",x"20",x"3a"),
  1314 => (x"00",x"0a",x"64",x"25"),
  1315 => (x"6e",x"49",x"20",x"20"),
  1316 => (x"6f",x"43",x"5f",x"74"),
  1317 => (x"20",x"3a",x"70",x"6d"),
  1318 => (x"20",x"20",x"20",x"20"),
  1319 => (x"20",x"20",x"20",x"20"),
  1320 => (x"0a",x"64",x"25",x"20"),
  1321 => (x"20",x"20",x"20",x"00"),
  1322 => (x"20",x"20",x"20",x"20"),
  1323 => (x"6f",x"68",x"73",x"20"),
  1324 => (x"20",x"64",x"6c",x"75"),
  1325 => (x"20",x"3a",x"65",x"62"),
  1326 => (x"64",x"25",x"20",x"20"),
  1327 => (x"20",x"20",x"00",x"0a"),
  1328 => (x"5f",x"72",x"74",x"53"),
  1329 => (x"70",x"6d",x"6f",x"43"),
  1330 => (x"20",x"20",x"20",x"3a"),
  1331 => (x"20",x"20",x"20",x"20"),
  1332 => (x"25",x"20",x"20",x"20"),
  1333 => (x"20",x"00",x"0a",x"73"),
  1334 => (x"20",x"20",x"20",x"20"),
  1335 => (x"73",x"20",x"20",x"20"),
  1336 => (x"6c",x"75",x"6f",x"68"),
  1337 => (x"65",x"62",x"20",x"64"),
  1338 => (x"20",x"20",x"20",x"3a"),
  1339 => (x"59",x"52",x"48",x"44"),
  1340 => (x"4e",x"4f",x"54",x"53"),
  1341 => (x"52",x"50",x"20",x"45"),
  1342 => (x"41",x"52",x"47",x"4f"),
  1343 => (x"53",x"20",x"2c",x"4d"),
  1344 => (x"20",x"45",x"4d",x"4f"),
  1345 => (x"49",x"52",x"54",x"53"),
  1346 => (x"00",x"0a",x"47",x"4e"),
  1347 => (x"5f",x"74",x"6e",x"49"),
  1348 => (x"6f",x"4c",x"5f",x"31"),
  1349 => (x"20",x"20",x"3a",x"63"),
  1350 => (x"20",x"20",x"20",x"20"),
  1351 => (x"20",x"20",x"20",x"20"),
  1352 => (x"0a",x"64",x"25",x"20"),
  1353 => (x"20",x"20",x"20",x"00"),
  1354 => (x"20",x"20",x"20",x"20"),
  1355 => (x"6f",x"68",x"73",x"20"),
  1356 => (x"20",x"64",x"6c",x"75"),
  1357 => (x"20",x"3a",x"65",x"62"),
  1358 => (x"64",x"25",x"20",x"20"),
  1359 => (x"6e",x"49",x"00",x"0a"),
  1360 => (x"5f",x"32",x"5f",x"74"),
  1361 => (x"3a",x"63",x"6f",x"4c"),
  1362 => (x"20",x"20",x"20",x"20"),
  1363 => (x"20",x"20",x"20",x"20"),
  1364 => (x"25",x"20",x"20",x"20"),
  1365 => (x"20",x"00",x"0a",x"64"),
  1366 => (x"20",x"20",x"20",x"20"),
  1367 => (x"73",x"20",x"20",x"20"),
  1368 => (x"6c",x"75",x"6f",x"68"),
  1369 => (x"65",x"62",x"20",x"64"),
  1370 => (x"20",x"20",x"20",x"3a"),
  1371 => (x"00",x"0a",x"64",x"25"),
  1372 => (x"5f",x"74",x"6e",x"49"),
  1373 => (x"6f",x"4c",x"5f",x"33"),
  1374 => (x"20",x"20",x"3a",x"63"),
  1375 => (x"20",x"20",x"20",x"20"),
  1376 => (x"20",x"20",x"20",x"20"),
  1377 => (x"0a",x"64",x"25",x"20"),
  1378 => (x"20",x"20",x"20",x"00"),
  1379 => (x"20",x"20",x"20",x"20"),
  1380 => (x"6f",x"68",x"73",x"20"),
  1381 => (x"20",x"64",x"6c",x"75"),
  1382 => (x"20",x"3a",x"65",x"62"),
  1383 => (x"64",x"25",x"20",x"20"),
  1384 => (x"6e",x"45",x"00",x"0a"),
  1385 => (x"4c",x"5f",x"6d",x"75"),
  1386 => (x"20",x"3a",x"63",x"6f"),
  1387 => (x"20",x"20",x"20",x"20"),
  1388 => (x"20",x"20",x"20",x"20"),
  1389 => (x"25",x"20",x"20",x"20"),
  1390 => (x"20",x"00",x"0a",x"64"),
  1391 => (x"20",x"20",x"20",x"20"),
  1392 => (x"73",x"20",x"20",x"20"),
  1393 => (x"6c",x"75",x"6f",x"68"),
  1394 => (x"65",x"62",x"20",x"64"),
  1395 => (x"20",x"20",x"20",x"3a"),
  1396 => (x"00",x"0a",x"64",x"25"),
  1397 => (x"5f",x"72",x"74",x"53"),
  1398 => (x"6f",x"4c",x"5f",x"31"),
  1399 => (x"20",x"20",x"3a",x"63"),
  1400 => (x"20",x"20",x"20",x"20"),
  1401 => (x"20",x"20",x"20",x"20"),
  1402 => (x"0a",x"73",x"25",x"20"),
  1403 => (x"20",x"20",x"20",x"00"),
  1404 => (x"20",x"20",x"20",x"20"),
  1405 => (x"6f",x"68",x"73",x"20"),
  1406 => (x"20",x"64",x"6c",x"75"),
  1407 => (x"20",x"3a",x"65",x"62"),
  1408 => (x"48",x"44",x"20",x"20"),
  1409 => (x"54",x"53",x"59",x"52"),
  1410 => (x"20",x"45",x"4e",x"4f"),
  1411 => (x"47",x"4f",x"52",x"50"),
  1412 => (x"2c",x"4d",x"41",x"52"),
  1413 => (x"53",x"27",x"31",x"20"),
  1414 => (x"54",x"53",x"20",x"54"),
  1415 => (x"47",x"4e",x"49",x"52"),
  1416 => (x"74",x"53",x"00",x"0a"),
  1417 => (x"5f",x"32",x"5f",x"72"),
  1418 => (x"3a",x"63",x"6f",x"4c"),
  1419 => (x"20",x"20",x"20",x"20"),
  1420 => (x"20",x"20",x"20",x"20"),
  1421 => (x"25",x"20",x"20",x"20"),
  1422 => (x"20",x"00",x"0a",x"73"),
  1423 => (x"20",x"20",x"20",x"20"),
  1424 => (x"73",x"20",x"20",x"20"),
  1425 => (x"6c",x"75",x"6f",x"68"),
  1426 => (x"65",x"62",x"20",x"64"),
  1427 => (x"20",x"20",x"20",x"3a"),
  1428 => (x"59",x"52",x"48",x"44"),
  1429 => (x"4e",x"4f",x"54",x"53"),
  1430 => (x"52",x"50",x"20",x"45"),
  1431 => (x"41",x"52",x"47",x"4f"),
  1432 => (x"32",x"20",x"2c",x"4d"),
  1433 => (x"20",x"44",x"4e",x"27"),
  1434 => (x"49",x"52",x"54",x"53"),
  1435 => (x"00",x"0a",x"47",x"4e"),
  1436 => (x"73",x"55",x"00",x"0a"),
  1437 => (x"74",x"20",x"72",x"65"),
  1438 => (x"3a",x"65",x"6d",x"69"),
  1439 => (x"0a",x"64",x"25",x"20"),
  1440 => (x"00",x"00",x"00",x"00"),
  1441 => (x"00",x"00",x"00",x"00"),
  1442 => (x"00",x"00",x"61",x"a8"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
