
package Toplevel_Config is
	constant Toplevel_UseUART : boolean := true;
	constant Toplevel_UseVGA : boolean := true;
	constant Toplevel_UseAudio : boolean := false;
	constant Toplevel_Frequency : integer := 100;
	constant Toplevel_SDRAMWidth : integer := 16;
end package;
