
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of OSDBoot_832_ROM is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"d4",x"01"),
     1 => (x"18",x"0e",x"87",x"d7"),
     2 => (x"3e",x"27",x"0e",x"1e"),
     3 => (x"0f",x"00",x"00",x"00"),
     4 => (x"80",x"ff",x"48",x"26"),
     5 => (x"27",x"4f",x"08",x"26"),
     6 => (x"00",x"00",x"00",x"23"),
     7 => (x"00",x"30",x"27",x"4f"),
     8 => (x"c2",x"4f",x"00",x"00"),
     9 => (x"27",x"4e",x"c0",x"c0"),
    10 => (x"00",x"00",x"02",x"dc"),
    11 => (x"87",x"fd",x"00",x"0f"),
    12 => (x"4e",x"c0",x"f0",x"c1"),
    13 => (x"00",x"00",x"3d",x"27"),
    14 => (x"fd",x"00",x"0f",x"00"),
    15 => (x"0e",x"4f",x"4f",x"87"),
    16 => (x"5c",x"5b",x"5a",x"5e"),
    17 => (x"d8",x"1e",x"0e",x"5d"),
    18 => (x"49",x"76",x"4d",x"66"),
    19 => (x"b7",x"c0",x"79",x"c0"),
    20 => (x"cd",x"c0",x"03",x"ad"),
    21 => (x"1e",x"ed",x"c0",x"87"),
    22 => (x"00",x"13",x"cb",x"27"),
    23 => (x"86",x"c4",x"0f",x"00"),
    24 => (x"9d",x"75",x"8d",x"0d"),
    25 => (x"87",x"c2",x"c1",x"02"),
    26 => (x"4a",x"75",x"4c",x"c0"),
    27 => (x"72",x"2a",x"b7",x"dc"),
    28 => (x"c4",x"9b",x"cf",x"4b"),
    29 => (x"02",x"9b",x"73",x"35"),
    30 => (x"76",x"87",x"c4",x"c0"),
    31 => (x"c9",x"79",x"c1",x"49"),
    32 => (x"c0",x"06",x"ab",x"b7"),
    33 => (x"f7",x"c0",x"87",x"c6"),
    34 => (x"87",x"c3",x"c0",x"83"),
    35 => (x"6e",x"83",x"f0",x"c0"),
    36 => (x"87",x"ca",x"c0",x"02"),
    37 => (x"cb",x"27",x"1e",x"73"),
    38 => (x"0f",x"00",x"00",x"13"),
    39 => (x"84",x"c1",x"86",x"c4"),
    40 => (x"04",x"ac",x"b7",x"c8"),
    41 => (x"c0",x"87",x"c3",x"ff"),
    42 => (x"f0",x"c0",x"87",x"cb"),
    43 => (x"13",x"cb",x"27",x"1e"),
    44 => (x"c4",x"0f",x"00",x"00"),
    45 => (x"26",x"48",x"c0",x"86"),
    46 => (x"4c",x"26",x"4d",x"26"),
    47 => (x"4a",x"26",x"4b",x"26"),
    48 => (x"5e",x"0e",x"4f",x"26"),
    49 => (x"5d",x"5c",x"5b",x"5a"),
    50 => (x"4c",x"c0",x"1e",x"0e"),
    51 => (x"79",x"c0",x"49",x"76"),
    52 => (x"d8",x"4b",x"a6",x"dc"),
    53 => (x"66",x"d8",x"4a",x"66"),
    54 => (x"dc",x"80",x"c1",x"48"),
    55 => (x"4d",x"12",x"58",x"a6"),
    56 => (x"c0",x"c0",x"c0",x"c1"),
    57 => (x"c0",x"c4",x"95",x"c0"),
    58 => (x"75",x"4d",x"95",x"b7"),
    59 => (x"d2",x"c4",x"02",x"9d"),
    60 => (x"c3",x"02",x"6e",x"87"),
    61 => (x"49",x"76",x"87",x"d7"),
    62 => (x"4a",x"75",x"79",x"c0"),
    63 => (x"02",x"ad",x"e3",x"c1"),
    64 => (x"c1",x"87",x"dd",x"c2"),
    65 => (x"c0",x"02",x"aa",x"e4"),
    66 => (x"ec",x"c1",x"87",x"d8"),
    67 => (x"c8",x"c2",x"02",x"aa"),
    68 => (x"aa",x"f3",x"c1",x"87"),
    69 => (x"87",x"e8",x"c1",x"02"),
    70 => (x"02",x"aa",x"f8",x"c1"),
    71 => (x"c2",x"87",x"f2",x"c0"),
    72 => (x"1e",x"ca",x"87",x"d3"),
    73 => (x"00",x"16",x"e8",x"27"),
    74 => (x"83",x"c4",x"1e",x"00"),
    75 => (x"8a",x"c4",x"4a",x"73"),
    76 => (x"3f",x"27",x"1e",x"6a"),
    77 => (x"0f",x"00",x"00",x"00"),
    78 => (x"4a",x"70",x"86",x"cc"),
    79 => (x"84",x"72",x"4c",x"74"),
    80 => (x"00",x"16",x"e8",x"27"),
    81 => (x"fa",x"27",x"1e",x"00"),
    82 => (x"0f",x"00",x"00",x"13"),
    83 => (x"d4",x"c2",x"86",x"c4"),
    84 => (x"27",x"1e",x"d0",x"87"),
    85 => (x"00",x"00",x"16",x"e8"),
    86 => (x"73",x"83",x"c4",x"1e"),
    87 => (x"6a",x"8a",x"c4",x"4a"),
    88 => (x"00",x"3f",x"27",x"1e"),
    89 => (x"cc",x"0f",x"00",x"00"),
    90 => (x"74",x"4a",x"70",x"86"),
    91 => (x"27",x"84",x"72",x"4c"),
    92 => (x"00",x"00",x"16",x"e8"),
    93 => (x"13",x"fa",x"27",x"1e"),
    94 => (x"c4",x"0f",x"00",x"00"),
    95 => (x"87",x"e5",x"c1",x"86"),
    96 => (x"4a",x"73",x"83",x"c4"),
    97 => (x"1e",x"6a",x"8a",x"c4"),
    98 => (x"00",x"13",x"fa",x"27"),
    99 => (x"86",x"c4",x"0f",x"00"),
   100 => (x"4c",x"74",x"4a",x"70"),
   101 => (x"cc",x"c1",x"84",x"72"),
   102 => (x"c1",x"49",x"76",x"87"),
   103 => (x"87",x"c5",x"c1",x"79"),
   104 => (x"4a",x"73",x"83",x"c4"),
   105 => (x"1e",x"6a",x"8a",x"c4"),
   106 => (x"00",x"13",x"cb",x"27"),
   107 => (x"86",x"c4",x"0f",x"00"),
   108 => (x"f0",x"c0",x"84",x"c1"),
   109 => (x"1e",x"e5",x"c0",x"87"),
   110 => (x"00",x"13",x"cb",x"27"),
   111 => (x"86",x"c4",x"0f",x"00"),
   112 => (x"cb",x"27",x"1e",x"75"),
   113 => (x"0f",x"00",x"00",x"13"),
   114 => (x"d8",x"c0",x"86",x"c4"),
   115 => (x"ad",x"e5",x"c0",x"87"),
   116 => (x"87",x"c7",x"c0",x"05"),
   117 => (x"79",x"c1",x"49",x"76"),
   118 => (x"75",x"87",x"ca",x"c0"),
   119 => (x"13",x"cb",x"27",x"1e"),
   120 => (x"c4",x"0f",x"00",x"00"),
   121 => (x"4a",x"66",x"d8",x"86"),
   122 => (x"c1",x"48",x"66",x"d8"),
   123 => (x"58",x"a6",x"dc",x"80"),
   124 => (x"c0",x"c1",x"4d",x"12"),
   125 => (x"95",x"c0",x"c0",x"c0"),
   126 => (x"95",x"b7",x"c0",x"c4"),
   127 => (x"05",x"9d",x"75",x"4d"),
   128 => (x"74",x"87",x"ee",x"fb"),
   129 => (x"4d",x"26",x"26",x"48"),
   130 => (x"4b",x"26",x"4c",x"26"),
   131 => (x"4f",x"26",x"4a",x"26"),
   132 => (x"5b",x"5a",x"5e",x"0e"),
   133 => (x"4a",x"66",x"cc",x"0e"),
   134 => (x"ff",x"c3",x"2a",x"d8"),
   135 => (x"4b",x"66",x"cc",x"9a"),
   136 => (x"fc",x"cf",x"2b",x"c8"),
   137 => (x"4a",x"72",x"9b",x"c0"),
   138 => (x"66",x"cc",x"b2",x"73"),
   139 => (x"c0",x"33",x"c8",x"4b"),
   140 => (x"c0",x"c0",x"f0",x"ff"),
   141 => (x"73",x"4a",x"72",x"9b"),
   142 => (x"4b",x"66",x"cc",x"b2"),
   143 => (x"fc",x"cf",x"33",x"d8"),
   144 => (x"9b",x"c0",x"c0",x"c0"),
   145 => (x"b2",x"73",x"4a",x"72"),
   146 => (x"4b",x"26",x"48",x"72"),
   147 => (x"4f",x"26",x"4a",x"26"),
   148 => (x"5b",x"5a",x"5e",x"0e"),
   149 => (x"4a",x"66",x"cc",x"0e"),
   150 => (x"ff",x"c3",x"2a",x"c8"),
   151 => (x"4b",x"66",x"cc",x"9a"),
   152 => (x"fc",x"cf",x"33",x"c8"),
   153 => (x"4a",x"72",x"9b",x"c0"),
   154 => (x"48",x"72",x"b2",x"73"),
   155 => (x"4a",x"26",x"4b",x"26"),
   156 => (x"5e",x"0e",x"4f",x"26"),
   157 => (x"cc",x"0e",x"5b",x"5a"),
   158 => (x"2a",x"d0",x"4a",x"66"),
   159 => (x"9a",x"ff",x"ff",x"cf"),
   160 => (x"4b",x"66",x"cc",x"4a"),
   161 => (x"c0",x"f0",x"33",x"d0"),
   162 => (x"4a",x"72",x"9b",x"c0"),
   163 => (x"48",x"72",x"b2",x"73"),
   164 => (x"4a",x"26",x"4b",x"26"),
   165 => (x"5e",x"0e",x"4f",x"26"),
   166 => (x"5d",x"5c",x"5b",x"5a"),
   167 => (x"4d",x"66",x"d8",x"0e"),
   168 => (x"66",x"d4",x"4c",x"c0"),
   169 => (x"2a",x"b7",x"dc",x"4a"),
   170 => (x"9b",x"cf",x"4b",x"72"),
   171 => (x"c4",x"48",x"66",x"d4"),
   172 => (x"58",x"a6",x"d8",x"30"),
   173 => (x"06",x"ab",x"b7",x"c9"),
   174 => (x"c0",x"87",x"c6",x"c0"),
   175 => (x"c3",x"c0",x"83",x"f7"),
   176 => (x"83",x"f0",x"c0",x"87"),
   177 => (x"c1",x"7d",x"97",x"73"),
   178 => (x"c8",x"84",x"c1",x"85"),
   179 => (x"ff",x"04",x"ac",x"b7"),
   180 => (x"4d",x"26",x"87",x"d0"),
   181 => (x"4b",x"26",x"4c",x"26"),
   182 => (x"4f",x"26",x"4a",x"26"),
   183 => (x"5b",x"5a",x"5e",x"0e"),
   184 => (x"cc",x"0e",x"5d",x"5c"),
   185 => (x"15",x"04",x"27",x"8e"),
   186 => (x"27",x"1e",x"00",x"00"),
   187 => (x"00",x"00",x"13",x"fa"),
   188 => (x"27",x"86",x"c4",x"0f"),
   189 => (x"00",x"00",x"12",x"2e"),
   190 => (x"72",x"4a",x"70",x"0f"),
   191 => (x"cf",x"c4",x"02",x"9a"),
   192 => (x"14",x"ed",x"27",x"87"),
   193 => (x"27",x"1e",x"00",x"00"),
   194 => (x"00",x"00",x"13",x"fa"),
   195 => (x"27",x"86",x"c4",x"0f"),
   196 => (x"00",x"00",x"04",x"7c"),
   197 => (x"72",x"4a",x"70",x"0f"),
   198 => (x"e5",x"c3",x"02",x"9a"),
   199 => (x"20",x"00",x"27",x"87"),
   200 => (x"27",x"1e",x"00",x"00"),
   201 => (x"00",x"00",x"14",x"c5"),
   202 => (x"0b",x"3b",x"27",x"1e"),
   203 => (x"c8",x"0f",x"00",x"00"),
   204 => (x"73",x"4b",x"70",x"86"),
   205 => (x"d7",x"c3",x"02",x"9b"),
   206 => (x"49",x"a6",x"c4",x"87"),
   207 => (x"00",x"20",x"00",x"27"),
   208 => (x"4d",x"c0",x"79",x"00"),
   209 => (x"9b",x"fc",x"83",x"c3"),
   210 => (x"00",x"20",x"00",x"27"),
   211 => (x"84",x"73",x"4c",x"00"),
   212 => (x"b9",x"27",x"1e",x"74"),
   213 => (x"1e",x"00",x"00",x"14"),
   214 => (x"00",x"0b",x"3b",x"27"),
   215 => (x"86",x"c8",x"0f",x"00"),
   216 => (x"9a",x"72",x"4a",x"70"),
   217 => (x"87",x"e8",x"c2",x"02"),
   218 => (x"ab",x"b7",x"ff",x"c7"),
   219 => (x"87",x"e0",x"c2",x"06"),
   220 => (x"c8",x"1e",x"c0",x"c8"),
   221 => (x"82",x"75",x"4a",x"66"),
   222 => (x"2e",x"27",x"1e",x"72"),
   223 => (x"0f",x"00",x"00",x"14"),
   224 => (x"4a",x"70",x"86",x"c8"),
   225 => (x"72",x"49",x"a6",x"c8"),
   226 => (x"24",x"49",x"76",x"79"),
   227 => (x"85",x"c0",x"c8",x"79"),
   228 => (x"c8",x"8b",x"c0",x"c8"),
   229 => (x"b7",x"6e",x"49",x"66"),
   230 => (x"da",x"c1",x"02",x"a9"),
   231 => (x"17",x"08",x"27",x"87"),
   232 => (x"75",x"1e",x"00",x"00"),
   233 => (x"02",x"96",x"27",x"1e"),
   234 => (x"c8",x"0f",x"00",x"00"),
   235 => (x"17",x"10",x"27",x"86"),
   236 => (x"c0",x"49",x"00",x"00"),
   237 => (x"11",x"27",x"51",x"e0"),
   238 => (x"1e",x"00",x"00",x"17"),
   239 => (x"27",x"1e",x"66",x"cc"),
   240 => (x"00",x"00",x"02",x"96"),
   241 => (x"27",x"86",x"c8",x"0f"),
   242 => (x"00",x"00",x"17",x"19"),
   243 => (x"51",x"e0",x"c0",x"49"),
   244 => (x"00",x"17",x"1a",x"27"),
   245 => (x"66",x"c4",x"1e",x"00"),
   246 => (x"02",x"96",x"27",x"1e"),
   247 => (x"c8",x"0f",x"00",x"00"),
   248 => (x"17",x"22",x"27",x"86"),
   249 => (x"c0",x"49",x"00",x"00"),
   250 => (x"17",x"08",x"27",x"51"),
   251 => (x"27",x"1e",x"00",x"00"),
   252 => (x"00",x"00",x"0c",x"a1"),
   253 => (x"c7",x"86",x"c4",x"0f"),
   254 => (x"01",x"ab",x"b7",x"ff"),
   255 => (x"c0",x"87",x"f1",x"fd"),
   256 => (x"d1",x"27",x"87",x"ce"),
   257 => (x"1e",x"00",x"00",x"14"),
   258 => (x"00",x"13",x"fa",x"27"),
   259 => (x"86",x"c4",x"0f",x"00"),
   260 => (x"cc",x"87",x"fd",x"ff"),
   261 => (x"26",x"4d",x"26",x"86"),
   262 => (x"26",x"4b",x"26",x"4c"),
   263 => (x"0e",x"4f",x"26",x"4a"),
   264 => (x"5c",x"5b",x"5a",x"5e"),
   265 => (x"66",x"d4",x"0e",x"5d"),
   266 => (x"dc",x"4c",x"c0",x"4d"),
   267 => (x"b7",x"c0",x"49",x"66"),
   268 => (x"fb",x"c0",x"06",x"a9"),
   269 => (x"c1",x"4b",x"15",x"87"),
   270 => (x"c0",x"c0",x"c0",x"c0"),
   271 => (x"b7",x"c0",x"c4",x"93"),
   272 => (x"66",x"d8",x"4b",x"93"),
   273 => (x"c1",x"4a",x"bf",x"97"),
   274 => (x"c0",x"c0",x"c0",x"c0"),
   275 => (x"b7",x"c0",x"c4",x"92"),
   276 => (x"66",x"d8",x"4a",x"92"),
   277 => (x"dc",x"80",x"c1",x"48"),
   278 => (x"b7",x"72",x"58",x"a6"),
   279 => (x"c5",x"c0",x"02",x"ab"),
   280 => (x"c0",x"48",x"c1",x"87"),
   281 => (x"84",x"c1",x"87",x"cc"),
   282 => (x"ac",x"b7",x"66",x"dc"),
   283 => (x"87",x"c5",x"ff",x"04"),
   284 => (x"4d",x"26",x"48",x"c0"),
   285 => (x"4b",x"26",x"4c",x"26"),
   286 => (x"4f",x"26",x"4a",x"26"),
   287 => (x"5b",x"5a",x"5e",x"0e"),
   288 => (x"27",x"0e",x"5d",x"5c"),
   289 => (x"00",x"00",x"19",x"30"),
   290 => (x"27",x"79",x"c0",x"49"),
   291 => (x"00",x"00",x"15",x"ee"),
   292 => (x"13",x"fa",x"27",x"1e"),
   293 => (x"c4",x"0f",x"00",x"00"),
   294 => (x"17",x"28",x"27",x"86"),
   295 => (x"c0",x"1e",x"00",x"00"),
   296 => (x"12",x"cf",x"27",x"1e"),
   297 => (x"c8",x"0f",x"00",x"00"),
   298 => (x"72",x"4a",x"70",x"86"),
   299 => (x"d3",x"c0",x"05",x"9a"),
   300 => (x"15",x"1a",x"27",x"87"),
   301 => (x"27",x"1e",x"00",x"00"),
   302 => (x"00",x"00",x"13",x"fa"),
   303 => (x"c0",x"86",x"c4",x"0f"),
   304 => (x"87",x"d8",x"cf",x"48"),
   305 => (x"00",x"15",x"fb",x"27"),
   306 => (x"fa",x"27",x"1e",x"00"),
   307 => (x"0f",x"00",x"00",x"13"),
   308 => (x"4c",x"c0",x"86",x"c4"),
   309 => (x"00",x"19",x"5c",x"27"),
   310 => (x"79",x"c1",x"49",x"00"),
   311 => (x"12",x"27",x"1e",x"c8"),
   312 => (x"1e",x"00",x"00",x"16"),
   313 => (x"00",x"17",x"5e",x"27"),
   314 => (x"1f",x"27",x"1e",x"00"),
   315 => (x"0f",x"00",x"00",x"04"),
   316 => (x"4a",x"70",x"86",x"cc"),
   317 => (x"c0",x"05",x"9a",x"72"),
   318 => (x"5c",x"27",x"87",x"c8"),
   319 => (x"49",x"00",x"00",x"19"),
   320 => (x"1e",x"c8",x"79",x"c0"),
   321 => (x"00",x"16",x"1b",x"27"),
   322 => (x"7a",x"27",x"1e",x"00"),
   323 => (x"1e",x"00",x"00",x"17"),
   324 => (x"00",x"04",x"1f",x"27"),
   325 => (x"86",x"cc",x"0f",x"00"),
   326 => (x"9a",x"72",x"4a",x"70"),
   327 => (x"87",x"c8",x"c0",x"05"),
   328 => (x"00",x"19",x"5c",x"27"),
   329 => (x"79",x"c0",x"49",x"00"),
   330 => (x"00",x"19",x"5c",x"27"),
   331 => (x"27",x"1e",x"bf",x"00"),
   332 => (x"00",x"00",x"16",x"24"),
   333 => (x"00",x"c2",x"27",x"1e"),
   334 => (x"c8",x"0f",x"00",x"00"),
   335 => (x"19",x"5c",x"27",x"86"),
   336 => (x"02",x"bf",x"00",x"00"),
   337 => (x"27",x"87",x"c0",x"c3"),
   338 => (x"00",x"00",x"17",x"28"),
   339 => (x"18",x"e6",x"27",x"4d"),
   340 => (x"27",x"4b",x"00",x"00"),
   341 => (x"00",x"00",x"19",x"26"),
   342 => (x"72",x"4a",x"bf",x"9f"),
   343 => (x"19",x"26",x"27",x"1e"),
   344 => (x"27",x"4a",x"00",x"00"),
   345 => (x"00",x"00",x"17",x"28"),
   346 => (x"d0",x"1e",x"72",x"8a"),
   347 => (x"1e",x"c0",x"c8",x"1e"),
   348 => (x"00",x"15",x"4c",x"27"),
   349 => (x"c2",x"27",x"1e",x"00"),
   350 => (x"0f",x"00",x"00",x"00"),
   351 => (x"4a",x"73",x"86",x"d4"),
   352 => (x"4c",x"6a",x"82",x"c8"),
   353 => (x"00",x"19",x"26",x"27"),
   354 => (x"4a",x"bf",x"9f",x"00"),
   355 => (x"b7",x"ea",x"d6",x"c5"),
   356 => (x"d3",x"c0",x"05",x"aa"),
   357 => (x"c8",x"4a",x"73",x"87"),
   358 => (x"27",x"1e",x"6a",x"82"),
   359 => (x"00",x"00",x"02",x"10"),
   360 => (x"70",x"86",x"c4",x"0f"),
   361 => (x"87",x"e4",x"c0",x"4c"),
   362 => (x"fe",x"c7",x"4a",x"75"),
   363 => (x"4a",x"6a",x"9f",x"82"),
   364 => (x"b7",x"d5",x"e9",x"ca"),
   365 => (x"d3",x"c0",x"02",x"aa"),
   366 => (x"15",x"2e",x"27",x"87"),
   367 => (x"27",x"1e",x"00",x"00"),
   368 => (x"00",x"00",x"13",x"fa"),
   369 => (x"c0",x"86",x"c4",x"0f"),
   370 => (x"87",x"d0",x"cb",x"48"),
   371 => (x"89",x"27",x"1e",x"74"),
   372 => (x"1e",x"00",x"00",x"15"),
   373 => (x"00",x"00",x"c2",x"27"),
   374 => (x"86",x"c8",x"0f",x"00"),
   375 => (x"00",x"17",x"28",x"27"),
   376 => (x"1e",x"74",x"1e",x"00"),
   377 => (x"00",x"12",x"cf",x"27"),
   378 => (x"86",x"c8",x"0f",x"00"),
   379 => (x"9a",x"72",x"4a",x"70"),
   380 => (x"87",x"c5",x"c0",x"05"),
   381 => (x"e3",x"ca",x"48",x"c0"),
   382 => (x"15",x"a1",x"27",x"87"),
   383 => (x"27",x"1e",x"00",x"00"),
   384 => (x"00",x"00",x"13",x"fa"),
   385 => (x"27",x"86",x"c4",x"0f"),
   386 => (x"00",x"00",x"16",x"37"),
   387 => (x"00",x"c2",x"27",x"1e"),
   388 => (x"c4",x"0f",x"00",x"00"),
   389 => (x"27",x"1e",x"c8",x"86"),
   390 => (x"00",x"00",x"16",x"4f"),
   391 => (x"17",x"7a",x"27",x"1e"),
   392 => (x"27",x"1e",x"00",x"00"),
   393 => (x"00",x"00",x"04",x"1f"),
   394 => (x"70",x"86",x"cc",x"0f"),
   395 => (x"05",x"9a",x"72",x"4a"),
   396 => (x"27",x"87",x"cb",x"c0"),
   397 => (x"00",x"00",x"19",x"30"),
   398 => (x"c0",x"79",x"c1",x"49"),
   399 => (x"1e",x"c8",x"87",x"f1"),
   400 => (x"00",x"16",x"58",x"27"),
   401 => (x"5e",x"27",x"1e",x"00"),
   402 => (x"1e",x"00",x"00",x"17"),
   403 => (x"00",x"04",x"1f",x"27"),
   404 => (x"86",x"cc",x"0f",x"00"),
   405 => (x"9a",x"72",x"4a",x"70"),
   406 => (x"87",x"d3",x"c0",x"02"),
   407 => (x"00",x"15",x"c8",x"27"),
   408 => (x"c2",x"27",x"1e",x"00"),
   409 => (x"0f",x"00",x"00",x"00"),
   410 => (x"48",x"c0",x"86",x"c4"),
   411 => (x"27",x"87",x"ed",x"c8"),
   412 => (x"00",x"00",x"19",x"26"),
   413 => (x"c1",x"4a",x"bf",x"97"),
   414 => (x"05",x"aa",x"b7",x"d5"),
   415 => (x"27",x"87",x"d0",x"c0"),
   416 => (x"00",x"00",x"19",x"27"),
   417 => (x"c2",x"4a",x"bf",x"97"),
   418 => (x"02",x"aa",x"b7",x"ea"),
   419 => (x"c0",x"87",x"c5",x"c0"),
   420 => (x"87",x"c8",x"c8",x"48"),
   421 => (x"00",x"17",x"28",x"27"),
   422 => (x"4a",x"bf",x"97",x"00"),
   423 => (x"aa",x"b7",x"e9",x"c3"),
   424 => (x"87",x"d5",x"c0",x"02"),
   425 => (x"00",x"17",x"28",x"27"),
   426 => (x"4a",x"bf",x"97",x"00"),
   427 => (x"aa",x"b7",x"eb",x"c3"),
   428 => (x"87",x"c5",x"c0",x"02"),
   429 => (x"e3",x"c7",x"48",x"c0"),
   430 => (x"17",x"33",x"27",x"87"),
   431 => (x"bf",x"97",x"00",x"00"),
   432 => (x"05",x"9a",x"72",x"4a"),
   433 => (x"27",x"87",x"cf",x"c0"),
   434 => (x"00",x"00",x"17",x"34"),
   435 => (x"c2",x"4a",x"bf",x"97"),
   436 => (x"c0",x"02",x"aa",x"b7"),
   437 => (x"48",x"c0",x"87",x"c5"),
   438 => (x"27",x"87",x"c1",x"c7"),
   439 => (x"00",x"00",x"17",x"35"),
   440 => (x"27",x"48",x"bf",x"97"),
   441 => (x"00",x"00",x"19",x"2c"),
   442 => (x"19",x"28",x"27",x"58"),
   443 => (x"4a",x"bf",x"00",x"00"),
   444 => (x"8b",x"c1",x"4b",x"72"),
   445 => (x"00",x"19",x"2c",x"27"),
   446 => (x"79",x"73",x"49",x"00"),
   447 => (x"1e",x"72",x"1e",x"73"),
   448 => (x"00",x"16",x"61",x"27"),
   449 => (x"c2",x"27",x"1e",x"00"),
   450 => (x"0f",x"00",x"00",x"00"),
   451 => (x"36",x"27",x"86",x"cc"),
   452 => (x"97",x"00",x"00",x"17"),
   453 => (x"82",x"74",x"4a",x"bf"),
   454 => (x"00",x"17",x"37",x"27"),
   455 => (x"4b",x"bf",x"97",x"00"),
   456 => (x"48",x"73",x"33",x"c8"),
   457 => (x"40",x"27",x"80",x"72"),
   458 => (x"58",x"00",x"00",x"19"),
   459 => (x"00",x"17",x"38",x"27"),
   460 => (x"48",x"bf",x"97",x"00"),
   461 => (x"00",x"19",x"54",x"27"),
   462 => (x"30",x"27",x"58",x"00"),
   463 => (x"bf",x"00",x"00",x"19"),
   464 => (x"87",x"df",x"c3",x"02"),
   465 => (x"e5",x"27",x"1e",x"c8"),
   466 => (x"1e",x"00",x"00",x"15"),
   467 => (x"00",x"17",x"7a",x"27"),
   468 => (x"1f",x"27",x"1e",x"00"),
   469 => (x"0f",x"00",x"00",x"04"),
   470 => (x"4a",x"70",x"86",x"cc"),
   471 => (x"c0",x"02",x"9a",x"72"),
   472 => (x"48",x"c0",x"87",x"c5"),
   473 => (x"27",x"87",x"f5",x"c4"),
   474 => (x"00",x"00",x"19",x"28"),
   475 => (x"48",x"73",x"4b",x"bf"),
   476 => (x"58",x"27",x"30",x"c4"),
   477 => (x"58",x"00",x"00",x"19"),
   478 => (x"00",x"19",x"4c",x"27"),
   479 => (x"79",x"73",x"49",x"00"),
   480 => (x"00",x"17",x"4d",x"27"),
   481 => (x"4a",x"bf",x"97",x"00"),
   482 => (x"4c",x"27",x"32",x"c8"),
   483 => (x"97",x"00",x"00",x"17"),
   484 => (x"4a",x"72",x"4c",x"bf"),
   485 => (x"4e",x"27",x"82",x"74"),
   486 => (x"97",x"00",x"00",x"17"),
   487 => (x"34",x"d0",x"4c",x"bf"),
   488 => (x"82",x"74",x"4a",x"72"),
   489 => (x"00",x"17",x"4f",x"27"),
   490 => (x"4c",x"bf",x"97",x"00"),
   491 => (x"4a",x"72",x"34",x"d8"),
   492 => (x"58",x"27",x"82",x"74"),
   493 => (x"49",x"00",x"00",x"19"),
   494 => (x"4a",x"72",x"79",x"72"),
   495 => (x"00",x"19",x"50",x"27"),
   496 => (x"72",x"92",x"bf",x"00"),
   497 => (x"19",x"3c",x"27",x"4a"),
   498 => (x"82",x"bf",x"00",x"00"),
   499 => (x"00",x"19",x"40",x"27"),
   500 => (x"79",x"72",x"49",x"00"),
   501 => (x"00",x"17",x"55",x"27"),
   502 => (x"4c",x"bf",x"97",x"00"),
   503 => (x"54",x"27",x"34",x"c8"),
   504 => (x"97",x"00",x"00",x"17"),
   505 => (x"4c",x"74",x"4d",x"bf"),
   506 => (x"56",x"27",x"84",x"75"),
   507 => (x"97",x"00",x"00",x"17"),
   508 => (x"35",x"d0",x"4d",x"bf"),
   509 => (x"84",x"75",x"4c",x"74"),
   510 => (x"00",x"17",x"57",x"27"),
   511 => (x"4d",x"bf",x"97",x"00"),
   512 => (x"35",x"d8",x"9d",x"cf"),
   513 => (x"84",x"75",x"4c",x"74"),
   514 => (x"00",x"19",x"44",x"27"),
   515 => (x"79",x"74",x"49",x"00"),
   516 => (x"4b",x"73",x"8c",x"c2"),
   517 => (x"48",x"73",x"93",x"74"),
   518 => (x"4c",x"27",x"80",x"72"),
   519 => (x"58",x"00",x"00",x"19"),
   520 => (x"27",x"87",x"f7",x"c1"),
   521 => (x"00",x"00",x"17",x"3a"),
   522 => (x"c8",x"4a",x"bf",x"97"),
   523 => (x"17",x"39",x"27",x"32"),
   524 => (x"bf",x"97",x"00",x"00"),
   525 => (x"73",x"4a",x"72",x"4b"),
   526 => (x"19",x"54",x"27",x"82"),
   527 => (x"72",x"49",x"00",x"00"),
   528 => (x"c7",x"32",x"c5",x"79"),
   529 => (x"2a",x"c9",x"82",x"ff"),
   530 => (x"00",x"19",x"4c",x"27"),
   531 => (x"79",x"72",x"49",x"00"),
   532 => (x"00",x"17",x"3f",x"27"),
   533 => (x"4b",x"bf",x"97",x"00"),
   534 => (x"3e",x"27",x"33",x"c8"),
   535 => (x"97",x"00",x"00",x"17"),
   536 => (x"4b",x"73",x"4c",x"bf"),
   537 => (x"58",x"27",x"83",x"74"),
   538 => (x"49",x"00",x"00",x"19"),
   539 => (x"4b",x"73",x"79",x"73"),
   540 => (x"00",x"19",x"50",x"27"),
   541 => (x"73",x"93",x"bf",x"00"),
   542 => (x"19",x"3c",x"27",x"4b"),
   543 => (x"83",x"bf",x"00",x"00"),
   544 => (x"00",x"19",x"48",x"27"),
   545 => (x"79",x"73",x"49",x"00"),
   546 => (x"00",x"19",x"44",x"27"),
   547 => (x"79",x"c0",x"49",x"00"),
   548 => (x"80",x"72",x"48",x"73"),
   549 => (x"00",x"19",x"44",x"27"),
   550 => (x"48",x"c1",x"58",x"00"),
   551 => (x"4c",x"26",x"4d",x"26"),
   552 => (x"4a",x"26",x"4b",x"26"),
   553 => (x"5e",x"0e",x"4f",x"26"),
   554 => (x"5d",x"5c",x"5b",x"5a"),
   555 => (x"19",x"30",x"27",x"0e"),
   556 => (x"02",x"bf",x"00",x"00"),
   557 => (x"d4",x"87",x"cf",x"c0"),
   558 => (x"b7",x"c7",x"4c",x"66"),
   559 => (x"4b",x"66",x"d4",x"2c"),
   560 => (x"c0",x"9b",x"ff",x"c1"),
   561 => (x"66",x"d4",x"87",x"cc"),
   562 => (x"2c",x"b7",x"c8",x"4c"),
   563 => (x"c3",x"4b",x"66",x"d4"),
   564 => (x"28",x"27",x"9b",x"ff"),
   565 => (x"1e",x"00",x"00",x"17"),
   566 => (x"00",x"19",x"3c",x"27"),
   567 => (x"74",x"4a",x"bf",x"00"),
   568 => (x"27",x"1e",x"72",x"82"),
   569 => (x"00",x"00",x"12",x"cf"),
   570 => (x"70",x"86",x"c8",x"0f"),
   571 => (x"05",x"9a",x"72",x"4a"),
   572 => (x"c0",x"87",x"c5",x"c0"),
   573 => (x"87",x"f2",x"c0",x"48"),
   574 => (x"00",x"19",x"30",x"27"),
   575 => (x"c0",x"02",x"bf",x"00"),
   576 => (x"4a",x"73",x"87",x"d7"),
   577 => (x"4a",x"72",x"92",x"c4"),
   578 => (x"00",x"17",x"28",x"27"),
   579 => (x"4d",x"6a",x"82",x"00"),
   580 => (x"ff",x"ff",x"ff",x"cf"),
   581 => (x"cf",x"c0",x"9d",x"ff"),
   582 => (x"c2",x"4a",x"73",x"87"),
   583 => (x"27",x"4a",x"72",x"92"),
   584 => (x"00",x"00",x"17",x"28"),
   585 => (x"4d",x"6a",x"9f",x"82"),
   586 => (x"4d",x"26",x"48",x"75"),
   587 => (x"4b",x"26",x"4c",x"26"),
   588 => (x"4f",x"26",x"4a",x"26"),
   589 => (x"5b",x"5a",x"5e",x"0e"),
   590 => (x"cc",x"0e",x"5d",x"5c"),
   591 => (x"ff",x"ff",x"cf",x"8e"),
   592 => (x"c0",x"4d",x"f8",x"ff"),
   593 => (x"27",x"49",x"76",x"4c"),
   594 => (x"00",x"00",x"19",x"44"),
   595 => (x"a6",x"c4",x"79",x"bf"),
   596 => (x"19",x"48",x"27",x"49"),
   597 => (x"79",x"bf",x"00",x"00"),
   598 => (x"00",x"19",x"30",x"27"),
   599 => (x"c0",x"02",x"bf",x"00"),
   600 => (x"28",x"27",x"87",x"cc"),
   601 => (x"bf",x"00",x"00",x"19"),
   602 => (x"c0",x"32",x"c4",x"4a"),
   603 => (x"4c",x"27",x"87",x"c9"),
   604 => (x"bf",x"00",x"00",x"19"),
   605 => (x"c8",x"32",x"c4",x"4a"),
   606 => (x"79",x"72",x"49",x"a6"),
   607 => (x"66",x"c8",x"4b",x"c0"),
   608 => (x"06",x"a9",x"c0",x"49"),
   609 => (x"73",x"87",x"d0",x"c3"),
   610 => (x"72",x"9a",x"cf",x"4a"),
   611 => (x"e4",x"c0",x"05",x"9a"),
   612 => (x"17",x"28",x"27",x"87"),
   613 => (x"c8",x"1e",x"00",x"00"),
   614 => (x"66",x"c8",x"4a",x"66"),
   615 => (x"cc",x"80",x"c1",x"48"),
   616 => (x"1e",x"72",x"58",x"a6"),
   617 => (x"00",x"12",x"cf",x"27"),
   618 => (x"86",x"c8",x"0f",x"00"),
   619 => (x"00",x"17",x"28",x"27"),
   620 => (x"c3",x"c0",x"4c",x"00"),
   621 => (x"84",x"e0",x"c0",x"87"),
   622 => (x"72",x"4a",x"6c",x"97"),
   623 => (x"cd",x"c2",x"02",x"9a"),
   624 => (x"4a",x"6c",x"97",x"87"),
   625 => (x"aa",x"b7",x"e5",x"c3"),
   626 => (x"87",x"c2",x"c2",x"02"),
   627 => (x"82",x"cb",x"4a",x"74"),
   628 => (x"d8",x"4a",x"6a",x"97"),
   629 => (x"05",x"9a",x"72",x"9a"),
   630 => (x"74",x"87",x"f3",x"c1"),
   631 => (x"13",x"fa",x"27",x"1e"),
   632 => (x"c4",x"0f",x"00",x"00"),
   633 => (x"c0",x"1e",x"cb",x"86"),
   634 => (x"74",x"1e",x"66",x"e8"),
   635 => (x"04",x"1f",x"27",x"1e"),
   636 => (x"cc",x"0f",x"00",x"00"),
   637 => (x"72",x"4a",x"70",x"86"),
   638 => (x"d1",x"c1",x"05",x"9a"),
   639 => (x"dc",x"4b",x"74",x"87"),
   640 => (x"66",x"e0",x"c0",x"83"),
   641 => (x"6b",x"82",x"c4",x"4a"),
   642 => (x"da",x"4b",x"74",x"7a"),
   643 => (x"66",x"e0",x"c0",x"83"),
   644 => (x"9f",x"82",x"c8",x"4a"),
   645 => (x"7a",x"70",x"48",x"6b"),
   646 => (x"30",x"27",x"4d",x"72"),
   647 => (x"bf",x"00",x"00",x"19"),
   648 => (x"87",x"d5",x"c0",x"02"),
   649 => (x"82",x"d4",x"4a",x"74"),
   650 => (x"c0",x"4a",x"6a",x"9f"),
   651 => (x"72",x"9a",x"ff",x"ff"),
   652 => (x"c4",x"30",x"d0",x"48"),
   653 => (x"c4",x"c0",x"58",x"a6"),
   654 => (x"c0",x"49",x"76",x"87"),
   655 => (x"6d",x"48",x"6e",x"79"),
   656 => (x"c0",x"7d",x"70",x"80"),
   657 => (x"c0",x"49",x"66",x"e0"),
   658 => (x"c1",x"48",x"c1",x"79"),
   659 => (x"83",x"c1",x"87",x"ce"),
   660 => (x"04",x"ab",x"66",x"c8"),
   661 => (x"cf",x"87",x"f0",x"fc"),
   662 => (x"f8",x"ff",x"ff",x"ff"),
   663 => (x"19",x"30",x"27",x"4d"),
   664 => (x"02",x"bf",x"00",x"00"),
   665 => (x"6e",x"87",x"f3",x"c0"),
   666 => (x"08",x"a6",x"27",x"1e"),
   667 => (x"c4",x"0f",x"00",x"00"),
   668 => (x"58",x"a6",x"c4",x"86"),
   669 => (x"9a",x"75",x"4a",x"6e"),
   670 => (x"c0",x"02",x"aa",x"75"),
   671 => (x"4a",x"6e",x"87",x"dc"),
   672 => (x"4a",x"72",x"8a",x"c2"),
   673 => (x"00",x"19",x"28",x"27"),
   674 => (x"27",x"92",x"bf",x"00"),
   675 => (x"00",x"00",x"19",x"40"),
   676 => (x"80",x"72",x"48",x"bf"),
   677 => (x"fb",x"58",x"a6",x"c8"),
   678 => (x"48",x"c0",x"87",x"e2"),
   679 => (x"ff",x"ff",x"ff",x"cf"),
   680 => (x"86",x"cc",x"4d",x"f8"),
   681 => (x"4c",x"26",x"4d",x"26"),
   682 => (x"4a",x"26",x"4b",x"26"),
   683 => (x"5e",x"0e",x"4f",x"26"),
   684 => (x"cc",x"0e",x"5b",x"5a"),
   685 => (x"c1",x"4a",x"bf",x"66"),
   686 => (x"49",x"66",x"cc",x"82"),
   687 => (x"4a",x"72",x"79",x"72"),
   688 => (x"00",x"19",x"2c",x"27"),
   689 => (x"72",x"9a",x"bf",x"00"),
   690 => (x"d3",x"c0",x"05",x"9a"),
   691 => (x"4a",x"66",x"cc",x"87"),
   692 => (x"1e",x"6a",x"82",x"c8"),
   693 => (x"00",x"08",x"a6",x"27"),
   694 => (x"86",x"c4",x"0f",x"00"),
   695 => (x"7a",x"73",x"4b",x"70"),
   696 => (x"4b",x"26",x"48",x"c1"),
   697 => (x"4f",x"26",x"4a",x"26"),
   698 => (x"5b",x"5a",x"5e",x"0e"),
   699 => (x"19",x"40",x"27",x"0e"),
   700 => (x"4a",x"bf",x"00",x"00"),
   701 => (x"c8",x"4b",x"66",x"cc"),
   702 => (x"c2",x"4b",x"6b",x"83"),
   703 => (x"27",x"4b",x"73",x"8b"),
   704 => (x"00",x"00",x"19",x"28"),
   705 => (x"4a",x"72",x"93",x"bf"),
   706 => (x"2c",x"27",x"82",x"73"),
   707 => (x"bf",x"00",x"00",x"19"),
   708 => (x"bf",x"66",x"cc",x"4b"),
   709 => (x"73",x"4a",x"72",x"9b"),
   710 => (x"1e",x"66",x"d0",x"82"),
   711 => (x"cf",x"27",x"1e",x"72"),
   712 => (x"0f",x"00",x"00",x"12"),
   713 => (x"4a",x"70",x"86",x"c8"),
   714 => (x"c0",x"05",x"9a",x"72"),
   715 => (x"48",x"c0",x"87",x"c5"),
   716 => (x"c1",x"87",x"c2",x"c0"),
   717 => (x"26",x"4b",x"26",x"48"),
   718 => (x"0e",x"4f",x"26",x"4a"),
   719 => (x"5c",x"5b",x"5a",x"5e"),
   720 => (x"66",x"d8",x"0e",x"5d"),
   721 => (x"1e",x"66",x"d4",x"4c"),
   722 => (x"00",x"19",x"60",x"27"),
   723 => (x"34",x"27",x"1e",x"00"),
   724 => (x"0f",x"00",x"00",x"09"),
   725 => (x"4a",x"70",x"86",x"c8"),
   726 => (x"c1",x"02",x"9a",x"72"),
   727 => (x"64",x"27",x"87",x"df"),
   728 => (x"bf",x"00",x"00",x"19"),
   729 => (x"82",x"ff",x"c7",x"4a"),
   730 => (x"4d",x"72",x"2a",x"c9"),
   731 => (x"df",x"27",x"4b",x"c0"),
   732 => (x"1e",x"00",x"00",x"0b"),
   733 => (x"00",x"13",x"fa",x"27"),
   734 => (x"86",x"c4",x"0f",x"00"),
   735 => (x"06",x"ad",x"b7",x"c0"),
   736 => (x"74",x"87",x"d0",x"c1"),
   737 => (x"19",x"60",x"27",x"1e"),
   738 => (x"27",x"1e",x"00",x"00"),
   739 => (x"00",x"00",x"0a",x"e8"),
   740 => (x"70",x"86",x"c8",x"0f"),
   741 => (x"05",x"9a",x"72",x"4a"),
   742 => (x"c0",x"87",x"c5",x"c0"),
   743 => (x"87",x"f5",x"c0",x"48"),
   744 => (x"00",x"19",x"60",x"27"),
   745 => (x"ae",x"27",x"1e",x"00"),
   746 => (x"0f",x"00",x"00",x"0a"),
   747 => (x"c0",x"c8",x"86",x"c4"),
   748 => (x"75",x"83",x"c1",x"84"),
   749 => (x"ff",x"04",x"ab",x"b7"),
   750 => (x"d6",x"c0",x"87",x"c9"),
   751 => (x"1e",x"66",x"d4",x"87"),
   752 => (x"00",x"0b",x"f8",x"27"),
   753 => (x"c2",x"27",x"1e",x"00"),
   754 => (x"0f",x"00",x"00",x"00"),
   755 => (x"48",x"c0",x"86",x"c8"),
   756 => (x"c1",x"87",x"c2",x"c0"),
   757 => (x"26",x"4d",x"26",x"48"),
   758 => (x"26",x"4b",x"26",x"4c"),
   759 => (x"4f",x"4f",x"26",x"4a"),
   760 => (x"65",x"6e",x"65",x"70"),
   761 => (x"69",x"66",x"20",x"64"),
   762 => (x"20",x"2c",x"65",x"6c"),
   763 => (x"64",x"61",x"6f",x"6c"),
   764 => (x"2e",x"67",x"6e",x"69"),
   765 => (x"00",x"0a",x"2e",x"2e"),
   766 => (x"27",x"6e",x"61",x"43"),
   767 => (x"70",x"6f",x"20",x"74"),
   768 => (x"25",x"20",x"6e",x"65"),
   769 => (x"1e",x"00",x"0a",x"73"),
   770 => (x"66",x"c8",x"1e",x"72"),
   771 => (x"87",x"d1",x"c0",x"02"),
   772 => (x"00",x"19",x"6c",x"27"),
   773 => (x"66",x"c8",x"49",x"00"),
   774 => (x"19",x"74",x"27",x"79"),
   775 => (x"c0",x"49",x"00",x"00"),
   776 => (x"19",x"74",x"27",x"79"),
   777 => (x"c0",x"05",x"00",x"00"),
   778 => (x"6c",x"27",x"87",x"db"),
   779 => (x"4a",x"00",x"00",x"19"),
   780 => (x"80",x"c4",x"48",x"72"),
   781 => (x"00",x"19",x"70",x"27"),
   782 => (x"70",x"27",x"58",x"00"),
   783 => (x"49",x"00",x"00",x"19"),
   784 => (x"ce",x"c0",x"79",x"6a"),
   785 => (x"19",x"70",x"27",x"87"),
   786 => (x"c8",x"48",x"00",x"00"),
   787 => (x"19",x"74",x"27",x"30"),
   788 => (x"27",x"58",x"00",x"00"),
   789 => (x"00",x"00",x"19",x"74"),
   790 => (x"72",x"82",x"c1",x"4a"),
   791 => (x"27",x"98",x"c3",x"48"),
   792 => (x"00",x"00",x"19",x"78"),
   793 => (x"19",x"70",x"27",x"58"),
   794 => (x"d8",x"4a",x"00",x"00"),
   795 => (x"48",x"72",x"2a",x"b7"),
   796 => (x"4f",x"26",x"4a",x"26"),
   797 => (x"5b",x"5a",x"5e",x"0e"),
   798 => (x"1e",x"66",x"cc",x"0e"),
   799 => (x"c4",x"87",x"c8",x"fe"),
   800 => (x"c0",x"4b",x"70",x"86"),
   801 => (x"02",x"9b",x"73",x"4a"),
   802 => (x"c1",x"87",x"ce",x"c0"),
   803 => (x"fd",x"1e",x"c0",x"82"),
   804 => (x"86",x"c4",x"87",x"f5"),
   805 => (x"ec",x"ff",x"4b",x"70"),
   806 => (x"26",x"48",x"72",x"87"),
   807 => (x"26",x"4a",x"26",x"4b"),
   808 => (x"5a",x"5e",x"0e",x"4f"),
   809 => (x"0e",x"5d",x"5c",x"5b"),
   810 => (x"f6",x"c0",x"8e",x"c8"),
   811 => (x"4c",x"c4",x"c0",x"e4"),
   812 => (x"c0",x"e4",x"f6",x"c0"),
   813 => (x"66",x"dc",x"4b",x"c0"),
   814 => (x"87",x"f8",x"fe",x"1e"),
   815 => (x"4a",x"70",x"86",x"c4"),
   816 => (x"85",x"c2",x"4d",x"72"),
   817 => (x"79",x"c1",x"49",x"76"),
   818 => (x"c1",x"7c",x"9f",x"d0"),
   819 => (x"7b",x"9f",x"c1",x"c0"),
   820 => (x"c0",x"4a",x"6b",x"9f"),
   821 => (x"9f",x"c0",x"7b",x"9f"),
   822 => (x"48",x"6b",x"9f",x"7b"),
   823 => (x"c4",x"58",x"a6",x"c8"),
   824 => (x"9a",x"72",x"9a",x"c0"),
   825 => (x"87",x"fd",x"c1",x"02"),
   826 => (x"e6",x"c0",x"02",x"6e"),
   827 => (x"49",x"66",x"c4",x"87"),
   828 => (x"a9",x"c6",x"c0",x"c8"),
   829 => (x"87",x"ed",x"c1",x"05"),
   830 => (x"79",x"c0",x"49",x"76"),
   831 => (x"9f",x"ca",x"eb",x"fa"),
   832 => (x"7b",x"9f",x"c1",x"7b"),
   833 => (x"75",x"7b",x"9f",x"c0"),
   834 => (x"9f",x"c0",x"7b",x"9f"),
   835 => (x"7b",x"9f",x"c0",x"7b"),
   836 => (x"75",x"87",x"d2",x"c1"),
   837 => (x"c8",x"2a",x"c1",x"4a"),
   838 => (x"c4",x"b2",x"c0",x"c0"),
   839 => (x"a9",x"72",x"49",x"66"),
   840 => (x"87",x"c1",x"c1",x"05"),
   841 => (x"fb",x"1e",x"66",x"dc"),
   842 => (x"86",x"c4",x"87",x"dd"),
   843 => (x"75",x"58",x"a6",x"c4"),
   844 => (x"72",x"8d",x"c1",x"4a"),
   845 => (x"de",x"c0",x"02",x"9a"),
   846 => (x"74",x"4c",x"6e",x"87"),
   847 => (x"9c",x"74",x"7b",x"97"),
   848 => (x"87",x"c9",x"c0",x"02"),
   849 => (x"fe",x"fa",x"1e",x"c0"),
   850 => (x"70",x"86",x"c4",x"87"),
   851 => (x"c1",x"4a",x"75",x"4c"),
   852 => (x"05",x"9a",x"72",x"8d"),
   853 => (x"c0",x"87",x"e4",x"ff"),
   854 => (x"c4",x"c0",x"e4",x"f6"),
   855 => (x"7c",x"9f",x"d1",x"4c"),
   856 => (x"c6",x"c0",x"48",x"c1"),
   857 => (x"7c",x"9f",x"d1",x"87"),
   858 => (x"c8",x"87",x"dd",x"fd"),
   859 => (x"26",x"4d",x"26",x"86"),
   860 => (x"26",x"4b",x"26",x"4c"),
   861 => (x"0e",x"4f",x"26",x"4a"),
   862 => (x"5c",x"5b",x"5a",x"5e"),
   863 => (x"8e",x"e4",x"c0",x"0e"),
   864 => (x"c0",x"4c",x"ff",x"c3"),
   865 => (x"c0",x"c0",x"e4",x"f6"),
   866 => (x"6b",x"7b",x"74",x"4b"),
   867 => (x"74",x"9a",x"74",x"4a"),
   868 => (x"74",x"48",x"6b",x"7b"),
   869 => (x"58",x"a6",x"c4",x"98"),
   870 => (x"30",x"c8",x"48",x"6e"),
   871 => (x"c8",x"58",x"a6",x"c8"),
   872 => (x"79",x"72",x"49",x"a6"),
   873 => (x"66",x"c4",x"4a",x"72"),
   874 => (x"6b",x"7b",x"74",x"b2"),
   875 => (x"d0",x"98",x"74",x"48"),
   876 => (x"66",x"cc",x"58",x"a6"),
   877 => (x"d4",x"30",x"d0",x"48"),
   878 => (x"a6",x"d4",x"58",x"a6"),
   879 => (x"72",x"79",x"72",x"49"),
   880 => (x"b2",x"66",x"d0",x"4a"),
   881 => (x"48",x"6b",x"7b",x"74"),
   882 => (x"a6",x"dc",x"98",x"74"),
   883 => (x"48",x"66",x"d8",x"58"),
   884 => (x"e0",x"c0",x"30",x"d8"),
   885 => (x"e0",x"c0",x"58",x"a6"),
   886 => (x"79",x"72",x"49",x"a6"),
   887 => (x"66",x"dc",x"4a",x"72"),
   888 => (x"c0",x"48",x"72",x"b2"),
   889 => (x"4c",x"26",x"86",x"e4"),
   890 => (x"4a",x"26",x"4b",x"26"),
   891 => (x"5e",x"0e",x"4f",x"26"),
   892 => (x"0e",x"5c",x"5b",x"5a"),
   893 => (x"ff",x"c3",x"8e",x"d8"),
   894 => (x"e4",x"f6",x"c0",x"4c"),
   895 => (x"74",x"4b",x"c0",x"c0"),
   896 => (x"74",x"4a",x"6b",x"7b"),
   897 => (x"c8",x"7b",x"74",x"9a"),
   898 => (x"74",x"48",x"6b",x"32"),
   899 => (x"58",x"a6",x"c4",x"98"),
   900 => (x"72",x"49",x"a6",x"c4"),
   901 => (x"6e",x"4a",x"72",x"79"),
   902 => (x"c8",x"7b",x"74",x"b2"),
   903 => (x"74",x"48",x"6b",x"32"),
   904 => (x"58",x"a6",x"cc",x"98"),
   905 => (x"72",x"49",x"a6",x"cc"),
   906 => (x"c8",x"4a",x"72",x"79"),
   907 => (x"7b",x"74",x"b2",x"66"),
   908 => (x"48",x"6b",x"32",x"c8"),
   909 => (x"a6",x"d4",x"98",x"74"),
   910 => (x"49",x"a6",x"d4",x"58"),
   911 => (x"4a",x"72",x"79",x"72"),
   912 => (x"72",x"b2",x"66",x"d0"),
   913 => (x"26",x"86",x"d8",x"48"),
   914 => (x"26",x"4b",x"26",x"4c"),
   915 => (x"0e",x"4f",x"26",x"4a"),
   916 => (x"5c",x"5b",x"5a",x"5e"),
   917 => (x"f6",x"c0",x"0e",x"5d"),
   918 => (x"4b",x"c0",x"c0",x"e4"),
   919 => (x"c3",x"48",x"66",x"d4"),
   920 => (x"7b",x"70",x"98",x"ff"),
   921 => (x"00",x"19",x"78",x"27"),
   922 => (x"c0",x"05",x"bf",x"00"),
   923 => (x"66",x"d8",x"87",x"c8"),
   924 => (x"dc",x"30",x"c9",x"48"),
   925 => (x"66",x"d8",x"58",x"a6"),
   926 => (x"72",x"2a",x"d8",x"4a"),
   927 => (x"98",x"ff",x"c3",x"48"),
   928 => (x"66",x"d8",x"7b",x"70"),
   929 => (x"72",x"2a",x"d0",x"4a"),
   930 => (x"98",x"ff",x"c3",x"48"),
   931 => (x"66",x"d8",x"7b",x"70"),
   932 => (x"72",x"2a",x"c8",x"4a"),
   933 => (x"98",x"ff",x"c3",x"48"),
   934 => (x"66",x"d8",x"7b",x"70"),
   935 => (x"98",x"ff",x"c3",x"48"),
   936 => (x"66",x"d4",x"7b",x"70"),
   937 => (x"72",x"2a",x"d0",x"4a"),
   938 => (x"98",x"ff",x"c3",x"48"),
   939 => (x"4d",x"6b",x"7b",x"70"),
   940 => (x"c9",x"9d",x"ff",x"c3"),
   941 => (x"c3",x"4c",x"ff",x"f0"),
   942 => (x"05",x"ad",x"b7",x"ff"),
   943 => (x"c3",x"87",x"d8",x"c0"),
   944 => (x"7b",x"72",x"4a",x"ff"),
   945 => (x"9d",x"72",x"4d",x"6b"),
   946 => (x"9c",x"74",x"8c",x"c1"),
   947 => (x"87",x"c7",x"c0",x"02"),
   948 => (x"02",x"ad",x"b7",x"72"),
   949 => (x"75",x"87",x"eb",x"ff"),
   950 => (x"16",x"85",x"27",x"1e"),
   951 => (x"27",x"1e",x"00",x"00"),
   952 => (x"00",x"00",x"00",x"c2"),
   953 => (x"75",x"86",x"c8",x"0f"),
   954 => (x"26",x"4d",x"26",x"48"),
   955 => (x"26",x"4b",x"26",x"4c"),
   956 => (x"0e",x"4f",x"26",x"4a"),
   957 => (x"0e",x"5b",x"5a",x"5e"),
   958 => (x"c0",x"e4",x"f6",x"c0"),
   959 => (x"4a",x"c0",x"4b",x"c0"),
   960 => (x"c1",x"7b",x"ff",x"c3"),
   961 => (x"b7",x"c8",x"c3",x"82"),
   962 => (x"f3",x"ff",x"04",x"aa"),
   963 => (x"26",x"4b",x"26",x"87"),
   964 => (x"0e",x"4f",x"26",x"4a"),
   965 => (x"5c",x"5b",x"5a",x"5e"),
   966 => (x"c0",x"c1",x"0e",x"5d"),
   967 => (x"c0",x"c0",x"c0",x"c0"),
   968 => (x"e4",x"f6",x"c0",x"4c"),
   969 => (x"27",x"4b",x"c0",x"c0"),
   970 => (x"00",x"00",x"0e",x"f3"),
   971 => (x"df",x"f8",x"c4",x"0f"),
   972 => (x"c0",x"1e",x"c0",x"4d"),
   973 => (x"f7",x"c1",x"f0",x"ff"),
   974 => (x"0e",x"4f",x"27",x"1e"),
   975 => (x"c8",x"0f",x"00",x"00"),
   976 => (x"c1",x"4a",x"70",x"86"),
   977 => (x"c1",x"05",x"aa",x"b7"),
   978 => (x"1e",x"72",x"87",x"dc"),
   979 => (x"00",x"0f",x"d4",x"27"),
   980 => (x"c2",x"27",x"1e",x"00"),
   981 => (x"0f",x"00",x"00",x"00"),
   982 => (x"ff",x"c3",x"86",x"c8"),
   983 => (x"c0",x"1e",x"74",x"7b"),
   984 => (x"e9",x"c1",x"f0",x"e1"),
   985 => (x"0e",x"4f",x"27",x"1e"),
   986 => (x"c8",x"0f",x"00",x"00"),
   987 => (x"72",x"4a",x"70",x"86"),
   988 => (x"d8",x"c0",x"05",x"9a"),
   989 => (x"27",x"1e",x"72",x"87"),
   990 => (x"00",x"00",x"0f",x"ca"),
   991 => (x"00",x"c2",x"27",x"1e"),
   992 => (x"c8",x"0f",x"00",x"00"),
   993 => (x"7b",x"ff",x"c3",x"86"),
   994 => (x"f3",x"c0",x"48",x"c1"),
   995 => (x"27",x"1e",x"72",x"87"),
   996 => (x"00",x"00",x"0f",x"de"),
   997 => (x"00",x"c2",x"27",x"1e"),
   998 => (x"c8",x"0f",x"00",x"00"),
   999 => (x"0e",x"f3",x"27",x"86"),
  1000 => (x"c0",x"0f",x"00",x"00"),
  1001 => (x"1e",x"72",x"87",x"d0"),
  1002 => (x"00",x"0f",x"e8",x"27"),
  1003 => (x"c2",x"27",x"1e",x"00"),
  1004 => (x"0f",x"00",x"00",x"00"),
  1005 => (x"8d",x"c1",x"86",x"c8"),
  1006 => (x"fd",x"05",x"9d",x"75"),
  1007 => (x"48",x"c0",x"87",x"f3"),
  1008 => (x"4c",x"26",x"4d",x"26"),
  1009 => (x"4a",x"26",x"4b",x"26"),
  1010 => (x"4d",x"43",x"4f",x"26"),
  1011 => (x"20",x"31",x"34",x"44"),
  1012 => (x"00",x"0a",x"64",x"25"),
  1013 => (x"35",x"44",x"4d",x"43"),
  1014 => (x"64",x"25",x"20",x"35"),
  1015 => (x"4d",x"43",x"00",x"0a"),
  1016 => (x"20",x"31",x"34",x"44"),
  1017 => (x"00",x"0a",x"64",x"25"),
  1018 => (x"35",x"44",x"4d",x"43"),
  1019 => (x"64",x"25",x"20",x"35"),
  1020 => (x"5e",x"0e",x"00",x"0a"),
  1021 => (x"5d",x"5c",x"5b",x"5a"),
  1022 => (x"f0",x"ff",x"c0",x"0e"),
  1023 => (x"c0",x"4d",x"c1",x"c1"),
  1024 => (x"c0",x"c0",x"e4",x"f6"),
  1025 => (x"7b",x"ff",x"c3",x"4b"),
  1026 => (x"00",x"10",x"84",x"27"),
  1027 => (x"fa",x"27",x"1e",x"00"),
  1028 => (x"0f",x"00",x"00",x"13"),
  1029 => (x"4c",x"d3",x"86",x"c4"),
  1030 => (x"1e",x"75",x"1e",x"c0"),
  1031 => (x"00",x"0e",x"4f",x"27"),
  1032 => (x"86",x"c8",x"0f",x"00"),
  1033 => (x"9a",x"72",x"4a",x"70"),
  1034 => (x"87",x"d8",x"c0",x"05"),
  1035 => (x"6e",x"27",x"1e",x"72"),
  1036 => (x"1e",x"00",x"00",x"10"),
  1037 => (x"00",x"00",x"c2",x"27"),
  1038 => (x"86",x"c8",x"0f",x"00"),
  1039 => (x"c1",x"7b",x"ff",x"c3"),
  1040 => (x"87",x"e0",x"c0",x"48"),
  1041 => (x"79",x"27",x"1e",x"72"),
  1042 => (x"1e",x"00",x"00",x"10"),
  1043 => (x"00",x"00",x"c2",x"27"),
  1044 => (x"86",x"c8",x"0f",x"00"),
  1045 => (x"00",x"0e",x"f3",x"27"),
  1046 => (x"8c",x"c1",x"0f",x"00"),
  1047 => (x"fe",x"05",x"9c",x"74"),
  1048 => (x"48",x"c0",x"87",x"f6"),
  1049 => (x"4c",x"26",x"4d",x"26"),
  1050 => (x"4a",x"26",x"4b",x"26"),
  1051 => (x"6e",x"69",x"4f",x"26"),
  1052 => (x"25",x"20",x"74",x"69"),
  1053 => (x"20",x"20",x"0a",x"64"),
  1054 => (x"69",x"6e",x"69",x"00"),
  1055 => (x"64",x"25",x"20",x"74"),
  1056 => (x"00",x"20",x"20",x"0a"),
  1057 => (x"5f",x"64",x"6d",x"43"),
  1058 => (x"74",x"69",x"6e",x"69"),
  1059 => (x"5e",x"0e",x"00",x"0a"),
  1060 => (x"5d",x"5c",x"5b",x"5a"),
  1061 => (x"ff",x"c3",x"1e",x"0e"),
  1062 => (x"e4",x"f6",x"c0",x"4d"),
  1063 => (x"27",x"4b",x"c0",x"c0"),
  1064 => (x"00",x"00",x"0e",x"f3"),
  1065 => (x"1e",x"ea",x"c6",x"0f"),
  1066 => (x"c1",x"f0",x"e1",x"c0"),
  1067 => (x"4f",x"27",x"1e",x"c8"),
  1068 => (x"0f",x"00",x"00",x"0e"),
  1069 => (x"4a",x"70",x"86",x"c8"),
  1070 => (x"17",x"27",x"1e",x"72"),
  1071 => (x"1e",x"00",x"00",x"12"),
  1072 => (x"00",x"00",x"c2",x"27"),
  1073 => (x"86",x"c8",x"0f",x"00"),
  1074 => (x"02",x"aa",x"b7",x"c1"),
  1075 => (x"27",x"87",x"cb",x"c0"),
  1076 => (x"00",x"00",x"0f",x"f2"),
  1077 => (x"c3",x"48",x"c0",x"0f"),
  1078 => (x"ee",x"27",x"87",x"db"),
  1079 => (x"0f",x"00",x"00",x"0d"),
  1080 => (x"4a",x"74",x"4c",x"70"),
  1081 => (x"9a",x"ff",x"ff",x"cf"),
  1082 => (x"aa",x"b7",x"ea",x"c6"),
  1083 => (x"87",x"db",x"c0",x"02"),
  1084 => (x"c0",x"27",x"1e",x"74"),
  1085 => (x"1e",x"00",x"00",x"11"),
  1086 => (x"00",x"00",x"c2",x"27"),
  1087 => (x"86",x"c8",x"0f",x"00"),
  1088 => (x"00",x"0f",x"f2",x"27"),
  1089 => (x"48",x"c0",x"0f",x"00"),
  1090 => (x"75",x"87",x"ea",x"c2"),
  1091 => (x"c0",x"49",x"76",x"7b"),
  1092 => (x"13",x"27",x"79",x"f1"),
  1093 => (x"0f",x"00",x"00",x"0f"),
  1094 => (x"9a",x"72",x"4a",x"70"),
  1095 => (x"87",x"eb",x"c1",x"02"),
  1096 => (x"ff",x"c0",x"1e",x"c0"),
  1097 => (x"1e",x"fa",x"c1",x"f0"),
  1098 => (x"00",x"0e",x"4f",x"27"),
  1099 => (x"86",x"c8",x"0f",x"00"),
  1100 => (x"9c",x"74",x"4c",x"70"),
  1101 => (x"87",x"c3",x"c1",x"05"),
  1102 => (x"d5",x"27",x"1e",x"74"),
  1103 => (x"1e",x"00",x"00",x"11"),
  1104 => (x"00",x"00",x"c2",x"27"),
  1105 => (x"86",x"c8",x"0f",x"00"),
  1106 => (x"4c",x"6b",x"7b",x"75"),
  1107 => (x"1e",x"74",x"9c",x"75"),
  1108 => (x"00",x"11",x"e1",x"27"),
  1109 => (x"c2",x"27",x"1e",x"00"),
  1110 => (x"0f",x"00",x"00",x"00"),
  1111 => (x"7b",x"75",x"86",x"c8"),
  1112 => (x"7b",x"75",x"7b",x"75"),
  1113 => (x"4a",x"74",x"7b",x"75"),
  1114 => (x"72",x"9a",x"c0",x"c1"),
  1115 => (x"c5",x"c0",x"02",x"9a"),
  1116 => (x"c0",x"48",x"c1",x"87"),
  1117 => (x"48",x"c0",x"87",x"ff"),
  1118 => (x"74",x"87",x"fa",x"c0"),
  1119 => (x"11",x"ef",x"27",x"1e"),
  1120 => (x"27",x"1e",x"00",x"00"),
  1121 => (x"00",x"00",x"00",x"c2"),
  1122 => (x"6e",x"86",x"c8",x"0f"),
  1123 => (x"a9",x"b7",x"c2",x"49"),
  1124 => (x"87",x"d3",x"c0",x"05"),
  1125 => (x"00",x"11",x"fb",x"27"),
  1126 => (x"c2",x"27",x"1e",x"00"),
  1127 => (x"0f",x"00",x"00",x"00"),
  1128 => (x"48",x"c0",x"86",x"c4"),
  1129 => (x"6e",x"87",x"ce",x"c0"),
  1130 => (x"c4",x"88",x"c1",x"48"),
  1131 => (x"05",x"6e",x"58",x"a6"),
  1132 => (x"c0",x"87",x"df",x"fd"),
  1133 => (x"4d",x"26",x"26",x"48"),
  1134 => (x"4b",x"26",x"4c",x"26"),
  1135 => (x"4f",x"26",x"4a",x"26"),
  1136 => (x"38",x"44",x"4d",x"43"),
  1137 => (x"72",x"20",x"34",x"5f"),
  1138 => (x"6f",x"70",x"73",x"65"),
  1139 => (x"3a",x"65",x"73",x"6e"),
  1140 => (x"0a",x"64",x"25",x"20"),
  1141 => (x"44",x"4d",x"43",x"00"),
  1142 => (x"25",x"20",x"38",x"35"),
  1143 => (x"20",x"20",x"0a",x"64"),
  1144 => (x"44",x"4d",x"43",x"00"),
  1145 => (x"32",x"5f",x"38",x"35"),
  1146 => (x"0a",x"64",x"25",x"20"),
  1147 => (x"43",x"00",x"20",x"20"),
  1148 => (x"38",x"35",x"44",x"4d"),
  1149 => (x"0a",x"64",x"25",x"20"),
  1150 => (x"53",x"00",x"20",x"20"),
  1151 => (x"20",x"43",x"48",x"44"),
  1152 => (x"74",x"69",x"6e",x"49"),
  1153 => (x"69",x"6c",x"61",x"69"),
  1154 => (x"69",x"74",x"61",x"7a"),
  1155 => (x"65",x"20",x"6e",x"6f"),
  1156 => (x"72",x"6f",x"72",x"72"),
  1157 => (x"63",x"00",x"0a",x"21"),
  1158 => (x"43",x"5f",x"64",x"6d"),
  1159 => (x"20",x"38",x"44",x"4d"),
  1160 => (x"70",x"73",x"65",x"72"),
  1161 => (x"65",x"73",x"6e",x"6f"),
  1162 => (x"64",x"25",x"20",x"3a"),
  1163 => (x"5e",x"0e",x"00",x"0a"),
  1164 => (x"5d",x"5c",x"5b",x"5a"),
  1165 => (x"e4",x"f6",x"c0",x"0e"),
  1166 => (x"c0",x"4d",x"c0",x"c0"),
  1167 => (x"c4",x"c0",x"e4",x"f6"),
  1168 => (x"19",x"78",x"27",x"4b"),
  1169 => (x"c1",x"49",x"00",x"00"),
  1170 => (x"e4",x"f6",x"c0",x"79"),
  1171 => (x"c0",x"49",x"c8",x"c0"),
  1172 => (x"4c",x"c7",x"79",x"e0"),
  1173 => (x"f3",x"27",x"7b",x"c3"),
  1174 => (x"0f",x"00",x"00",x"0e"),
  1175 => (x"ff",x"c3",x"7b",x"c2"),
  1176 => (x"c0",x"1e",x"c0",x"7d"),
  1177 => (x"c0",x"c1",x"d0",x"e5"),
  1178 => (x"0e",x"4f",x"27",x"1e"),
  1179 => (x"c8",x"0f",x"00",x"00"),
  1180 => (x"c1",x"4a",x"70",x"86"),
  1181 => (x"c0",x"05",x"aa",x"b7"),
  1182 => (x"4c",x"c1",x"87",x"c2"),
  1183 => (x"05",x"ac",x"b7",x"c2"),
  1184 => (x"c0",x"87",x"c5",x"c0"),
  1185 => (x"87",x"f8",x"c0",x"48"),
  1186 => (x"9c",x"74",x"8c",x"c1"),
  1187 => (x"87",x"c4",x"ff",x"05"),
  1188 => (x"00",x"10",x"8e",x"27"),
  1189 => (x"7c",x"27",x"0f",x"00"),
  1190 => (x"58",x"00",x"00",x"19"),
  1191 => (x"00",x"19",x"78",x"27"),
  1192 => (x"c0",x"05",x"bf",x"00"),
  1193 => (x"1e",x"c1",x"87",x"d0"),
  1194 => (x"c1",x"f0",x"ff",x"c0"),
  1195 => (x"4f",x"27",x"1e",x"d0"),
  1196 => (x"0f",x"00",x"00",x"0e"),
  1197 => (x"ff",x"c3",x"86",x"c8"),
  1198 => (x"c3",x"7b",x"c3",x"7d"),
  1199 => (x"48",x"c1",x"7d",x"ff"),
  1200 => (x"4c",x"26",x"4d",x"26"),
  1201 => (x"4a",x"26",x"4b",x"26"),
  1202 => (x"c0",x"1e",x"4f",x"26"),
  1203 => (x"0e",x"4f",x"26",x"48"),
  1204 => (x"5c",x"5b",x"5a",x"5e"),
  1205 => (x"8e",x"c8",x"0e",x"5d"),
  1206 => (x"4d",x"66",x"e0",x"c0"),
  1207 => (x"c0",x"e4",x"f6",x"c0"),
  1208 => (x"49",x"76",x"4b",x"c0"),
  1209 => (x"1e",x"75",x"79",x"c0"),
  1210 => (x"1e",x"66",x"e0",x"c0"),
  1211 => (x"00",x"13",x"b4",x"27"),
  1212 => (x"c2",x"27",x"1e",x"00"),
  1213 => (x"0f",x"00",x"00",x"00"),
  1214 => (x"ff",x"c3",x"86",x"cc"),
  1215 => (x"e4",x"f6",x"c0",x"7b"),
  1216 => (x"c2",x"49",x"c4",x"c0"),
  1217 => (x"e4",x"f6",x"c0",x"79"),
  1218 => (x"c1",x"49",x"c8",x"c0"),
  1219 => (x"7b",x"ff",x"c3",x"79"),
  1220 => (x"c0",x"1e",x"66",x"dc"),
  1221 => (x"d1",x"c1",x"f0",x"ff"),
  1222 => (x"0e",x"4f",x"27",x"1e"),
  1223 => (x"c8",x"0f",x"00",x"00"),
  1224 => (x"58",x"a6",x"c8",x"86"),
  1225 => (x"c0",x"02",x"66",x"c4"),
  1226 => (x"66",x"c4",x"87",x"d8"),
  1227 => (x"66",x"e0",x"c0",x"1e"),
  1228 => (x"13",x"94",x"27",x"1e"),
  1229 => (x"27",x"1e",x"00",x"00"),
  1230 => (x"00",x"00",x"00",x"c2"),
  1231 => (x"c1",x"86",x"cc",x"0f"),
  1232 => (x"ee",x"c5",x"87",x"c4"),
  1233 => (x"c3",x"4c",x"df",x"cd"),
  1234 => (x"4a",x"6b",x"7b",x"ff"),
  1235 => (x"c3",x"9a",x"ff",x"c3"),
  1236 => (x"05",x"aa",x"b7",x"fe"),
  1237 => (x"c0",x"87",x"dc",x"c0"),
  1238 => (x"0d",x"77",x"27",x"4a"),
  1239 => (x"70",x"0f",x"00",x"00"),
  1240 => (x"c1",x"85",x"c4",x"7d"),
  1241 => (x"b7",x"c0",x"c2",x"82"),
  1242 => (x"ec",x"ff",x"04",x"aa"),
  1243 => (x"76",x"4c",x"c1",x"87"),
  1244 => (x"c1",x"79",x"c1",x"49"),
  1245 => (x"05",x"9c",x"74",x"8c"),
  1246 => (x"c3",x"87",x"cc",x"ff"),
  1247 => (x"f6",x"c0",x"7b",x"ff"),
  1248 => (x"49",x"c4",x"c0",x"e4"),
  1249 => (x"48",x"6e",x"79",x"c3"),
  1250 => (x"4d",x"26",x"86",x"c8"),
  1251 => (x"4b",x"26",x"4c",x"26"),
  1252 => (x"4f",x"26",x"4a",x"26"),
  1253 => (x"64",x"61",x"65",x"52"),
  1254 => (x"6d",x"6f",x"63",x"20"),
  1255 => (x"64",x"6e",x"61",x"6d"),
  1256 => (x"69",x"61",x"66",x"20"),
  1257 => (x"20",x"64",x"65",x"6c"),
  1258 => (x"25",x"20",x"74",x"61"),
  1259 => (x"25",x"28",x"20",x"64"),
  1260 => (x"00",x"0a",x"29",x"64"),
  1261 => (x"72",x"5f",x"64",x"73"),
  1262 => (x"5f",x"64",x"61",x"65"),
  1263 => (x"74",x"63",x"65",x"73"),
  1264 => (x"25",x"20",x"72",x"6f"),
  1265 => (x"25",x"20",x"2c",x"64"),
  1266 => (x"1e",x"00",x"0a",x"64"),
  1267 => (x"c0",x"1e",x"1e",x"72"),
  1268 => (x"c0",x"c0",x"e8",x"f6"),
  1269 => (x"c4",x"48",x"6a",x"4a"),
  1270 => (x"a6",x"c4",x"98",x"c0"),
  1271 => (x"c0",x"05",x"6e",x"58"),
  1272 => (x"48",x"6a",x"87",x"cd"),
  1273 => (x"c4",x"98",x"c0",x"c4"),
  1274 => (x"02",x"6e",x"58",x"a6"),
  1275 => (x"cc",x"87",x"f3",x"ff"),
  1276 => (x"66",x"cc",x"7a",x"66"),
  1277 => (x"4a",x"26",x"26",x"48"),
  1278 => (x"5e",x"0e",x"4f",x"26"),
  1279 => (x"0e",x"5c",x"5b",x"5a"),
  1280 => (x"c0",x"4b",x"66",x"d0"),
  1281 => (x"c1",x"4a",x"13",x"4c"),
  1282 => (x"c0",x"c0",x"c0",x"c0"),
  1283 => (x"b7",x"c0",x"c4",x"92"),
  1284 => (x"1e",x"72",x"4a",x"92"),
  1285 => (x"00",x"13",x"cb",x"27"),
  1286 => (x"86",x"c4",x"0f",x"00"),
  1287 => (x"9a",x"72",x"84",x"c1"),
  1288 => (x"87",x"e1",x"ff",x"05"),
  1289 => (x"4c",x"26",x"48",x"74"),
  1290 => (x"4a",x"26",x"4b",x"26"),
  1291 => (x"5e",x"0e",x"4f",x"26"),
  1292 => (x"5d",x"5c",x"5b",x"5a"),
  1293 => (x"c0",x"8e",x"c8",x"0e"),
  1294 => (x"dc",x"4c",x"66",x"e0"),
  1295 => (x"49",x"76",x"4a",x"66"),
  1296 => (x"b7",x"c0",x"79",x"c0"),
  1297 => (x"e2",x"c1",x"06",x"ac"),
  1298 => (x"c8",x"4b",x"12",x"87"),
  1299 => (x"c0",x"8c",x"c1",x"33"),
  1300 => (x"c0",x"06",x"ac",x"b7"),
  1301 => (x"48",x"12",x"87",x"c8"),
  1302 => (x"c0",x"58",x"a6",x"c8"),
  1303 => (x"a6",x"c4",x"87",x"c5"),
  1304 => (x"73",x"79",x"c0",x"49"),
  1305 => (x"b3",x"66",x"c4",x"4b"),
  1306 => (x"8c",x"c1",x"33",x"c8"),
  1307 => (x"06",x"ac",x"b7",x"c0"),
  1308 => (x"12",x"87",x"c5",x"c0"),
  1309 => (x"87",x"c2",x"c0",x"4d"),
  1310 => (x"4b",x"73",x"4d",x"c0"),
  1311 => (x"33",x"c8",x"b3",x"75"),
  1312 => (x"b7",x"c0",x"8c",x"c1"),
  1313 => (x"c8",x"c0",x"06",x"ac"),
  1314 => (x"c8",x"48",x"12",x"87"),
  1315 => (x"c5",x"c0",x"58",x"a6"),
  1316 => (x"49",x"a6",x"c4",x"87"),
  1317 => (x"4b",x"73",x"79",x"c0"),
  1318 => (x"73",x"b3",x"66",x"c4"),
  1319 => (x"c4",x"80",x"6e",x"48"),
  1320 => (x"8c",x"c1",x"58",x"a6"),
  1321 => (x"01",x"ac",x"b7",x"c0"),
  1322 => (x"6e",x"87",x"de",x"fe"),
  1323 => (x"26",x"86",x"c8",x"48"),
  1324 => (x"26",x"4c",x"26",x"4d"),
  1325 => (x"26",x"4a",x"26",x"4b"),
  1326 => (x"45",x"48",x"43",x"4f"),
  1327 => (x"55",x"53",x"4b",x"43"),
  1328 => (x"4e",x"49",x"42",x"4d"),
  1329 => (x"44",x"53",x"4f",x"00"),
  1330 => (x"30",x"32",x"33",x"38"),
  1331 => (x"53",x"59",x"53",x"31"),
  1332 => (x"61",x"6e",x"55",x"00"),
  1333 => (x"20",x"65",x"6c",x"62"),
  1334 => (x"6c",x"20",x"6f",x"74"),
  1335 => (x"74",x"61",x"63",x"6f"),
  1336 => (x"61",x"70",x"20",x"65"),
  1337 => (x"74",x"69",x"74",x"72"),
  1338 => (x"0a",x"6e",x"6f",x"69"),
  1339 => (x"6e",x"75",x"48",x"00"),
  1340 => (x"67",x"6e",x"69",x"74"),
  1341 => (x"72",x"6f",x"66",x"20"),
  1342 => (x"72",x"61",x"70",x"20"),
  1343 => (x"69",x"74",x"69",x"74"),
  1344 => (x"00",x"0a",x"6e",x"6f"),
  1345 => (x"74",x"69",x"6e",x"49"),
  1346 => (x"69",x"6c",x"61",x"69"),
  1347 => (x"67",x"6e",x"69",x"7a"),
  1348 => (x"20",x"44",x"53",x"20"),
  1349 => (x"64",x"72",x"61",x"63"),
  1350 => (x"65",x"52",x"00",x"0a"),
  1351 => (x"6f",x"20",x"64",x"61"),
  1352 => (x"42",x"4d",x"20",x"66"),
  1353 => (x"61",x"66",x"20",x"52"),
  1354 => (x"64",x"65",x"6c",x"69"),
  1355 => (x"6f",x"4e",x"00",x"0a"),
  1356 => (x"72",x"61",x"70",x"20"),
  1357 => (x"69",x"74",x"69",x"74"),
  1358 => (x"73",x"20",x"6e",x"6f"),
  1359 => (x"61",x"6e",x"67",x"69"),
  1360 => (x"65",x"72",x"75",x"74"),
  1361 => (x"75",x"6f",x"66",x"20"),
  1362 => (x"00",x"0a",x"64",x"6e"),
  1363 => (x"73",x"52",x"42",x"4d"),
  1364 => (x"3a",x"65",x"7a",x"69"),
  1365 => (x"2c",x"64",x"25",x"20"),
  1366 => (x"72",x"61",x"70",x"20"),
  1367 => (x"69",x"74",x"69",x"74"),
  1368 => (x"69",x"73",x"6e",x"6f"),
  1369 => (x"20",x"3a",x"65",x"7a"),
  1370 => (x"20",x"2c",x"64",x"25"),
  1371 => (x"73",x"66",x"66",x"6f"),
  1372 => (x"6f",x"20",x"74",x"65"),
  1373 => (x"69",x"73",x"20",x"66"),
  1374 => (x"25",x"20",x"3a",x"67"),
  1375 => (x"73",x"20",x"2c",x"64"),
  1376 => (x"30",x"20",x"67",x"69"),
  1377 => (x"0a",x"78",x"25",x"78"),
  1378 => (x"61",x"65",x"52",x"00"),
  1379 => (x"67",x"6e",x"69",x"64"),
  1380 => (x"6f",x"6f",x"62",x"20"),
  1381 => (x"65",x"73",x"20",x"74"),
  1382 => (x"72",x"6f",x"74",x"63"),
  1383 => (x"0a",x"64",x"25",x"20"),
  1384 => (x"61",x"65",x"52",x"00"),
  1385 => (x"6f",x"62",x"20",x"64"),
  1386 => (x"73",x"20",x"74",x"6f"),
  1387 => (x"6f",x"74",x"63",x"65"),
  1388 => (x"72",x"66",x"20",x"72"),
  1389 => (x"66",x"20",x"6d",x"6f"),
  1390 => (x"74",x"73",x"72",x"69"),
  1391 => (x"72",x"61",x"70",x"20"),
  1392 => (x"69",x"74",x"69",x"74"),
  1393 => (x"00",x"0a",x"6e",x"6f"),
  1394 => (x"75",x"73",x"6e",x"55"),
  1395 => (x"72",x"6f",x"70",x"70"),
  1396 => (x"20",x"64",x"65",x"74"),
  1397 => (x"74",x"72",x"61",x"70"),
  1398 => (x"6f",x"69",x"74",x"69"),
  1399 => (x"79",x"74",x"20",x"6e"),
  1400 => (x"0d",x"21",x"65",x"70"),
  1401 => (x"54",x"41",x"46",x"00"),
  1402 => (x"20",x"20",x"32",x"33"),
  1403 => (x"65",x"52",x"00",x"20"),
  1404 => (x"6e",x"69",x"64",x"61"),
  1405 => (x"42",x"4d",x"20",x"67"),
  1406 => (x"4d",x"00",x"0a",x"52"),
  1407 => (x"73",x"20",x"52",x"42"),
  1408 => (x"65",x"63",x"63",x"75"),
  1409 => (x"75",x"66",x"73",x"73"),
  1410 => (x"20",x"79",x"6c",x"6c"),
  1411 => (x"64",x"61",x"65",x"72"),
  1412 => (x"41",x"46",x"00",x"0a"),
  1413 => (x"20",x"36",x"31",x"54"),
  1414 => (x"46",x"00",x"20",x"20"),
  1415 => (x"32",x"33",x"54",x"41"),
  1416 => (x"00",x"20",x"20",x"20"),
  1417 => (x"74",x"72",x"61",x"50"),
  1418 => (x"6f",x"69",x"74",x"69"),
  1419 => (x"75",x"6f",x"63",x"6e"),
  1420 => (x"25",x"20",x"74",x"6e"),
  1421 => (x"48",x"00",x"0a",x"64"),
  1422 => (x"69",x"74",x"6e",x"75"),
  1423 => (x"66",x"20",x"67",x"6e"),
  1424 => (x"66",x"20",x"72",x"6f"),
  1425 => (x"73",x"65",x"6c",x"69"),
  1426 => (x"65",x"74",x"73",x"79"),
  1427 => (x"46",x"00",x"0a",x"6d"),
  1428 => (x"32",x"33",x"54",x"41"),
  1429 => (x"00",x"20",x"20",x"20"),
  1430 => (x"31",x"54",x"41",x"46"),
  1431 => (x"20",x"20",x"20",x"36"),
  1432 => (x"75",x"6c",x"43",x"00"),
  1433 => (x"72",x"65",x"74",x"73"),
  1434 => (x"7a",x"69",x"73",x"20"),
  1435 => (x"25",x"20",x"3a",x"65"),
  1436 => (x"43",x"20",x"2c",x"64"),
  1437 => (x"74",x"73",x"75",x"6c"),
  1438 => (x"6d",x"20",x"72",x"65"),
  1439 => (x"2c",x"6b",x"73",x"61"),
  1440 => (x"0a",x"64",x"25",x"20"),
  1441 => (x"74",x"6f",x"47",x"00"),
  1442 => (x"73",x"65",x"72",x"20"),
  1443 => (x"20",x"74",x"6c",x"75"),
  1444 => (x"0a",x"20",x"64",x"25"),
  1445 => (x"0a",x"20",x"64",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
