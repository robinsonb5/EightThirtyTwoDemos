
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"3b",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"38"),
    10 => (x"20",x"00",x"27",x"4f"),
    11 => (x"27",x"4e",x"00",x"00"),
    12 => (x"00",x"00",x"13",x"64"),
    13 => (x"87",x"fd",x"00",x"0f"),
    14 => (x"4f",x"87",x"fd",x"00"),
    15 => (x"ff",x"86",x"fc",x"1e"),
    16 => (x"48",x"69",x"49",x"c0"),
    17 => (x"c4",x"98",x"c0",x"c4"),
    18 => (x"02",x"6e",x"58",x"a6"),
    19 => (x"66",x"c8",x"87",x"f4"),
    20 => (x"8e",x"fc",x"48",x"79"),
    21 => (x"5e",x"0e",x"4f",x"26"),
    22 => (x"cc",x"0e",x"5c",x"5b"),
    23 => (x"4c",x"c0",x"4b",x"66"),
    24 => (x"ff",x"c3",x"4a",x"13"),
    25 => (x"02",x"9a",x"72",x"9a"),
    26 => (x"49",x"72",x"87",x"d5"),
    27 => (x"cb",x"ff",x"1e",x"71"),
    28 => (x"c1",x"86",x"c4",x"87"),
    29 => (x"c3",x"4a",x"13",x"84"),
    30 => (x"9a",x"72",x"9a",x"ff"),
    31 => (x"74",x"87",x"eb",x"05"),
    32 => (x"26",x"4c",x"26",x"48"),
    33 => (x"0e",x"4f",x"26",x"4b"),
    34 => (x"5d",x"5c",x"5b",x"5e"),
    35 => (x"c0",x"86",x"f0",x"0e"),
    36 => (x"48",x"a6",x"c4",x"4b"),
    37 => (x"e4",x"c0",x"78",x"c0"),
    38 => (x"e0",x"c0",x"4c",x"a6"),
    39 => (x"c1",x"48",x"49",x"66"),
    40 => (x"a6",x"e4",x"c0",x"80"),
    41 => (x"fe",x"4a",x"11",x"58"),
    42 => (x"72",x"ba",x"82",x"c0"),
    43 => (x"d3",x"c4",x"02",x"9a"),
    44 => (x"02",x"66",x"c4",x"87"),
    45 => (x"c4",x"87",x"e2",x"c3"),
    46 => (x"78",x"c0",x"48",x"a6"),
    47 => (x"f0",x"c0",x"49",x"72"),
    48 => (x"f2",x"c2",x"02",x"aa"),
    49 => (x"a9",x"e3",x"c1",x"87"),
    50 => (x"87",x"f3",x"c2",x"02"),
    51 => (x"02",x"a9",x"e4",x"c1"),
    52 => (x"c1",x"87",x"e1",x"c0"),
    53 => (x"c2",x"02",x"a9",x"ec"),
    54 => (x"f0",x"c1",x"87",x"dd"),
    55 => (x"87",x"d4",x"02",x"a9"),
    56 => (x"02",x"a9",x"f3",x"c1"),
    57 => (x"c1",x"87",x"fc",x"c1"),
    58 => (x"c7",x"02",x"a9",x"f5"),
    59 => (x"a9",x"f8",x"c1",x"87"),
    60 => (x"87",x"dc",x"c2",x"05"),
    61 => (x"49",x"74",x"84",x"c4"),
    62 => (x"48",x"76",x"89",x"c4"),
    63 => (x"02",x"6e",x"78",x"69"),
    64 => (x"c8",x"87",x"d3",x"c1"),
    65 => (x"cc",x"78",x"c0",x"80"),
    66 => (x"78",x"c0",x"48",x"a6"),
    67 => (x"b7",x"dc",x"49",x"6e"),
    68 => (x"cf",x"4a",x"71",x"29"),
    69 => (x"c4",x"48",x"6e",x"9a"),
    70 => (x"58",x"a6",x"c4",x"30"),
    71 => (x"c5",x"02",x"9a",x"72"),
    72 => (x"48",x"a6",x"c8",x"87"),
    73 => (x"aa",x"c9",x"78",x"c1"),
    74 => (x"c0",x"87",x"c5",x"06"),
    75 => (x"87",x"c3",x"82",x"f7"),
    76 => (x"c8",x"82",x"f0",x"c0"),
    77 => (x"87",x"c9",x"02",x"66"),
    78 => (x"ff",x"fb",x"1e",x"72"),
    79 => (x"c1",x"86",x"c4",x"87"),
    80 => (x"48",x"66",x"cc",x"83"),
    81 => (x"a6",x"d0",x"80",x"c1"),
    82 => (x"48",x"66",x"cc",x"58"),
    83 => (x"04",x"a8",x"b7",x"c8"),
    84 => (x"c1",x"87",x"f9",x"fe"),
    85 => (x"f0",x"c0",x"87",x"d7"),
    86 => (x"87",x"e0",x"fb",x"1e"),
    87 => (x"83",x"c1",x"86",x"c4"),
    88 => (x"c4",x"87",x"ca",x"c1"),
    89 => (x"c4",x"49",x"74",x"84"),
    90 => (x"fb",x"1e",x"69",x"89"),
    91 => (x"86",x"c4",x"87",x"e8"),
    92 => (x"83",x"71",x"49",x"70"),
    93 => (x"c4",x"87",x"f6",x"c0"),
    94 => (x"78",x"c1",x"48",x"a6"),
    95 => (x"c4",x"87",x"ee",x"c0"),
    96 => (x"c4",x"49",x"74",x"84"),
    97 => (x"fa",x"1e",x"69",x"89"),
    98 => (x"86",x"c4",x"87",x"f2"),
    99 => (x"87",x"dd",x"83",x"c1"),
   100 => (x"e7",x"fa",x"1e",x"72"),
   101 => (x"d4",x"86",x"c4",x"87"),
   102 => (x"aa",x"e5",x"c0",x"87"),
   103 => (x"c4",x"87",x"c7",x"05"),
   104 => (x"78",x"c1",x"48",x"a6"),
   105 => (x"1e",x"72",x"87",x"c7"),
   106 => (x"c4",x"87",x"d1",x"fa"),
   107 => (x"66",x"e0",x"c0",x"86"),
   108 => (x"80",x"c1",x"48",x"49"),
   109 => (x"58",x"a6",x"e4",x"c0"),
   110 => (x"c0",x"fe",x"4a",x"11"),
   111 => (x"9a",x"72",x"ba",x"82"),
   112 => (x"87",x"ed",x"fb",x"05"),
   113 => (x"8e",x"f0",x"48",x"73"),
   114 => (x"4c",x"26",x"4d",x"26"),
   115 => (x"4f",x"26",x"4b",x"26"),
   116 => (x"e8",x"0e",x"5e",x"0e"),
   117 => (x"4a",x"d4",x"ff",x"86"),
   118 => (x"6a",x"7a",x"ff",x"c3"),
   119 => (x"7a",x"ff",x"c3",x"49"),
   120 => (x"30",x"c8",x"48",x"6a"),
   121 => (x"c8",x"58",x"a6",x"c4"),
   122 => (x"b1",x"6e",x"59",x"a6"),
   123 => (x"6a",x"7a",x"ff",x"c3"),
   124 => (x"cc",x"30",x"d0",x"48"),
   125 => (x"a6",x"d0",x"58",x"a6"),
   126 => (x"b1",x"66",x"c8",x"59"),
   127 => (x"6a",x"7a",x"ff",x"c3"),
   128 => (x"d4",x"30",x"d8",x"48"),
   129 => (x"a6",x"d8",x"58",x"a6"),
   130 => (x"b1",x"66",x"d0",x"59"),
   131 => (x"8e",x"e8",x"48",x"71"),
   132 => (x"5e",x"0e",x"4f",x"26"),
   133 => (x"ff",x"86",x"f4",x"0e"),
   134 => (x"ff",x"c3",x"4a",x"d4"),
   135 => (x"c3",x"49",x"6a",x"7a"),
   136 => (x"48",x"71",x"7a",x"ff"),
   137 => (x"a6",x"c4",x"30",x"c8"),
   138 => (x"6e",x"49",x"6a",x"58"),
   139 => (x"7a",x"ff",x"c3",x"b1"),
   140 => (x"30",x"c8",x"48",x"71"),
   141 => (x"6a",x"58",x"a6",x"c8"),
   142 => (x"b1",x"66",x"c4",x"49"),
   143 => (x"71",x"7a",x"ff",x"c3"),
   144 => (x"cc",x"30",x"c8",x"48"),
   145 => (x"49",x"6a",x"58",x"a6"),
   146 => (x"71",x"b1",x"66",x"c8"),
   147 => (x"26",x"8e",x"f4",x"48"),
   148 => (x"5b",x"5e",x"0e",x"4f"),
   149 => (x"c3",x"0e",x"5d",x"5c"),
   150 => (x"d4",x"ff",x"4d",x"ff"),
   151 => (x"48",x"66",x"d0",x"4c"),
   152 => (x"70",x"98",x"ff",x"c3"),
   153 => (x"c0",x"d2",x"c1",x"7c"),
   154 => (x"87",x"c8",x"05",x"bf"),
   155 => (x"c9",x"48",x"66",x"d4"),
   156 => (x"58",x"a6",x"d8",x"30"),
   157 => (x"d8",x"49",x"66",x"d4"),
   158 => (x"c3",x"48",x"71",x"29"),
   159 => (x"7c",x"70",x"98",x"ff"),
   160 => (x"d0",x"49",x"66",x"d4"),
   161 => (x"c3",x"48",x"71",x"29"),
   162 => (x"7c",x"70",x"98",x"ff"),
   163 => (x"c8",x"49",x"66",x"d4"),
   164 => (x"c3",x"48",x"71",x"29"),
   165 => (x"7c",x"70",x"98",x"ff"),
   166 => (x"c3",x"48",x"66",x"d4"),
   167 => (x"7c",x"70",x"98",x"ff"),
   168 => (x"d0",x"49",x"66",x"d0"),
   169 => (x"c3",x"48",x"71",x"29"),
   170 => (x"7c",x"70",x"98",x"ff"),
   171 => (x"f0",x"c9",x"4b",x"6c"),
   172 => (x"ab",x"75",x"4a",x"ff"),
   173 => (x"75",x"87",x"ce",x"05"),
   174 => (x"c1",x"4b",x"6c",x"7c"),
   175 => (x"87",x"c5",x"02",x"8a"),
   176 => (x"f2",x"02",x"ab",x"75"),
   177 => (x"26",x"48",x"73",x"87"),
   178 => (x"26",x"4c",x"26",x"4d"),
   179 => (x"1e",x"4f",x"26",x"4b"),
   180 => (x"d4",x"ff",x"49",x"c0"),
   181 => (x"78",x"ff",x"c3",x"48"),
   182 => (x"c8",x"c3",x"81",x"c1"),
   183 => (x"f1",x"04",x"a9",x"b7"),
   184 => (x"0e",x"4f",x"26",x"87"),
   185 => (x"5d",x"5c",x"5b",x"5e"),
   186 => (x"f0",x"ff",x"c0",x"0e"),
   187 => (x"c1",x"4d",x"f7",x"c1"),
   188 => (x"c0",x"c0",x"c0",x"c0"),
   189 => (x"d6",x"ff",x"4b",x"c0"),
   190 => (x"df",x"f8",x"c4",x"87"),
   191 => (x"75",x"1e",x"c0",x"4c"),
   192 => (x"87",x"cd",x"fd",x"1e"),
   193 => (x"a8",x"c1",x"86",x"c8"),
   194 => (x"87",x"e5",x"c0",x"05"),
   195 => (x"c3",x"48",x"d4",x"ff"),
   196 => (x"1e",x"73",x"78",x"ff"),
   197 => (x"c1",x"f0",x"e1",x"c0"),
   198 => (x"f4",x"fc",x"1e",x"e9"),
   199 => (x"70",x"86",x"c8",x"87"),
   200 => (x"87",x"ca",x"05",x"98"),
   201 => (x"c3",x"48",x"d4",x"ff"),
   202 => (x"48",x"c1",x"78",x"ff"),
   203 => (x"de",x"fe",x"87",x"cb"),
   204 => (x"05",x"8c",x"c1",x"87"),
   205 => (x"c0",x"87",x"c6",x"ff"),
   206 => (x"26",x"4d",x"26",x"48"),
   207 => (x"26",x"4b",x"26",x"4c"),
   208 => (x"5b",x"5e",x"0e",x"4f"),
   209 => (x"ff",x"c0",x"0e",x"5c"),
   210 => (x"4c",x"c1",x"c1",x"f0"),
   211 => (x"c3",x"48",x"d4",x"ff"),
   212 => (x"e5",x"c0",x"78",x"ff"),
   213 => (x"fd",x"f3",x"1e",x"d8"),
   214 => (x"d3",x"86",x"c4",x"87"),
   215 => (x"74",x"1e",x"c0",x"4b"),
   216 => (x"87",x"ed",x"fb",x"1e"),
   217 => (x"98",x"70",x"86",x"c8"),
   218 => (x"ff",x"87",x"ca",x"05"),
   219 => (x"ff",x"c3",x"48",x"d4"),
   220 => (x"cb",x"48",x"c1",x"78"),
   221 => (x"87",x"d7",x"fd",x"87"),
   222 => (x"ff",x"05",x"8b",x"c1"),
   223 => (x"48",x"c0",x"87",x"df"),
   224 => (x"4b",x"26",x"4c",x"26"),
   225 => (x"5e",x"0e",x"4f",x"26"),
   226 => (x"0e",x"5d",x"5c",x"5b"),
   227 => (x"fc",x"4c",x"d4",x"ff"),
   228 => (x"ea",x"c6",x"87",x"fd"),
   229 => (x"f0",x"e1",x"c0",x"1e"),
   230 => (x"fa",x"1e",x"c8",x"c1"),
   231 => (x"86",x"c8",x"87",x"f3"),
   232 => (x"1e",x"73",x"4b",x"70"),
   233 => (x"f3",x"1e",x"d2",x"d2"),
   234 => (x"86",x"c8",x"87",x"dd"),
   235 => (x"c8",x"02",x"ab",x"c1"),
   236 => (x"87",x"cd",x"fe",x"87"),
   237 => (x"cf",x"c2",x"48",x"c0"),
   238 => (x"87",x"d6",x"f9",x"87"),
   239 => (x"ff",x"cf",x"49",x"70"),
   240 => (x"ea",x"c6",x"99",x"ff"),
   241 => (x"87",x"c8",x"02",x"a9"),
   242 => (x"c0",x"87",x"f6",x"fd"),
   243 => (x"87",x"f8",x"c1",x"48"),
   244 => (x"c0",x"7c",x"ff",x"c3"),
   245 => (x"ca",x"fc",x"4d",x"f1"),
   246 => (x"02",x"98",x"70",x"87"),
   247 => (x"c0",x"87",x"d0",x"c1"),
   248 => (x"f0",x"ff",x"c0",x"1e"),
   249 => (x"f9",x"1e",x"fa",x"c1"),
   250 => (x"86",x"c8",x"87",x"e7"),
   251 => (x"9b",x"73",x"4b",x"70"),
   252 => (x"87",x"f1",x"c0",x"05"),
   253 => (x"d0",x"d1",x"1e",x"73"),
   254 => (x"87",x"cb",x"f2",x"1e"),
   255 => (x"ff",x"c3",x"86",x"c8"),
   256 => (x"73",x"4b",x"6c",x"7c"),
   257 => (x"1e",x"dc",x"d1",x"1e"),
   258 => (x"c8",x"87",x"fc",x"f1"),
   259 => (x"7c",x"ff",x"c3",x"86"),
   260 => (x"73",x"7c",x"7c",x"7c"),
   261 => (x"99",x"c0",x"c1",x"49"),
   262 => (x"c1",x"87",x"c5",x"02"),
   263 => (x"87",x"e8",x"c0",x"48"),
   264 => (x"e3",x"c0",x"48",x"c0"),
   265 => (x"d1",x"1e",x"73",x"87"),
   266 => (x"da",x"f1",x"1e",x"ea"),
   267 => (x"c2",x"86",x"c8",x"87"),
   268 => (x"87",x"cc",x"05",x"ad"),
   269 => (x"f1",x"1e",x"f6",x"d1"),
   270 => (x"86",x"c4",x"87",x"cd"),
   271 => (x"87",x"c8",x"48",x"c0"),
   272 => (x"fe",x"05",x"8d",x"c1"),
   273 => (x"48",x"c0",x"87",x"d0"),
   274 => (x"4c",x"26",x"4d",x"26"),
   275 => (x"4f",x"26",x"4b",x"26"),
   276 => (x"35",x"44",x"4d",x"43"),
   277 => (x"64",x"25",x"20",x"38"),
   278 => (x"00",x"20",x"20",x"0a"),
   279 => (x"35",x"44",x"4d",x"43"),
   280 => (x"20",x"32",x"5f",x"38"),
   281 => (x"20",x"0a",x"64",x"25"),
   282 => (x"4d",x"43",x"00",x"20"),
   283 => (x"20",x"38",x"35",x"44"),
   284 => (x"20",x"0a",x"64",x"25"),
   285 => (x"44",x"53",x"00",x"20"),
   286 => (x"49",x"20",x"43",x"48"),
   287 => (x"69",x"74",x"69",x"6e"),
   288 => (x"7a",x"69",x"6c",x"61"),
   289 => (x"6f",x"69",x"74",x"61"),
   290 => (x"72",x"65",x"20",x"6e"),
   291 => (x"21",x"72",x"6f",x"72"),
   292 => (x"6d",x"63",x"00",x"0a"),
   293 => (x"4d",x"43",x"5f",x"64"),
   294 => (x"72",x"20",x"38",x"44"),
   295 => (x"6f",x"70",x"73",x"65"),
   296 => (x"3a",x"65",x"73",x"6e"),
   297 => (x"0a",x"64",x"25",x"20"),
   298 => (x"5b",x"5e",x"0e",x"00"),
   299 => (x"fc",x"0e",x"5d",x"5c"),
   300 => (x"4c",x"d0",x"ff",x"86"),
   301 => (x"4b",x"c0",x"c0",x"c8"),
   302 => (x"48",x"c0",x"d2",x"c1"),
   303 => (x"d2",x"d6",x"78",x"c1"),
   304 => (x"87",x"d2",x"ee",x"1e"),
   305 => (x"4d",x"c7",x"86",x"c4"),
   306 => (x"98",x"73",x"48",x"6c"),
   307 => (x"6e",x"58",x"a6",x"c4"),
   308 => (x"6c",x"87",x"cc",x"02"),
   309 => (x"c4",x"98",x"73",x"48"),
   310 => (x"05",x"6e",x"58",x"a6"),
   311 => (x"c0",x"87",x"f4",x"ff"),
   312 => (x"87",x"eb",x"f7",x"7c"),
   313 => (x"98",x"73",x"48",x"6c"),
   314 => (x"6e",x"58",x"a6",x"c4"),
   315 => (x"6c",x"87",x"cc",x"02"),
   316 => (x"c4",x"98",x"73",x"48"),
   317 => (x"05",x"6e",x"58",x"a6"),
   318 => (x"c1",x"87",x"f4",x"ff"),
   319 => (x"c0",x"1e",x"c0",x"7c"),
   320 => (x"c0",x"c1",x"d0",x"e5"),
   321 => (x"87",x"c9",x"f5",x"1e"),
   322 => (x"a8",x"c1",x"86",x"c8"),
   323 => (x"87",x"c2",x"c0",x"05"),
   324 => (x"ad",x"c2",x"4d",x"c1"),
   325 => (x"87",x"cd",x"c0",x"05"),
   326 => (x"ec",x"1e",x"cd",x"d6"),
   327 => (x"86",x"c4",x"87",x"f8"),
   328 => (x"de",x"c1",x"48",x"c0"),
   329 => (x"05",x"8d",x"c1",x"87"),
   330 => (x"f9",x"87",x"dd",x"fe"),
   331 => (x"d2",x"c1",x"87",x"d8"),
   332 => (x"d2",x"c1",x"58",x"c4"),
   333 => (x"c0",x"05",x"bf",x"c0"),
   334 => (x"1e",x"c1",x"87",x"cd"),
   335 => (x"c1",x"f0",x"ff",x"c0"),
   336 => (x"cc",x"f4",x"1e",x"d0"),
   337 => (x"ff",x"86",x"c8",x"87"),
   338 => (x"ff",x"c3",x"48",x"d4"),
   339 => (x"87",x"ca",x"ca",x"78"),
   340 => (x"58",x"c8",x"d2",x"c1"),
   341 => (x"bf",x"c4",x"d2",x"c1"),
   342 => (x"1e",x"d6",x"d6",x"1e"),
   343 => (x"c8",x"87",x"e8",x"ec"),
   344 => (x"73",x"48",x"6c",x"86"),
   345 => (x"58",x"a6",x"c4",x"98"),
   346 => (x"cc",x"c0",x"02",x"6e"),
   347 => (x"73",x"48",x"6c",x"87"),
   348 => (x"58",x"a6",x"c4",x"98"),
   349 => (x"f4",x"ff",x"05",x"6e"),
   350 => (x"ff",x"7c",x"c0",x"87"),
   351 => (x"ff",x"c3",x"48",x"d4"),
   352 => (x"fc",x"48",x"c1",x"78"),
   353 => (x"26",x"4d",x"26",x"8e"),
   354 => (x"26",x"4b",x"26",x"4c"),
   355 => (x"52",x"45",x"49",x"4f"),
   356 => (x"50",x"53",x"00",x"52"),
   357 => (x"44",x"53",x"00",x"49"),
   358 => (x"72",x"61",x"63",x"20"),
   359 => (x"69",x"73",x"20",x"64"),
   360 => (x"69",x"20",x"65",x"7a"),
   361 => (x"64",x"25",x"20",x"73"),
   362 => (x"5e",x"0e",x"00",x"0a"),
   363 => (x"0e",x"5d",x"5c",x"5b"),
   364 => (x"c0",x"c8",x"86",x"fc"),
   365 => (x"ff",x"c3",x"4d",x"c0"),
   366 => (x"4b",x"d4",x"ff",x"4c"),
   367 => (x"d0",x"ff",x"7b",x"74"),
   368 => (x"98",x"75",x"48",x"bf"),
   369 => (x"6e",x"58",x"a6",x"c4"),
   370 => (x"87",x"ce",x"c0",x"02"),
   371 => (x"48",x"bf",x"d0",x"ff"),
   372 => (x"a6",x"c4",x"98",x"75"),
   373 => (x"ff",x"05",x"6e",x"58"),
   374 => (x"d0",x"ff",x"87",x"f2"),
   375 => (x"78",x"c1",x"c4",x"48"),
   376 => (x"66",x"d4",x"7b",x"74"),
   377 => (x"f0",x"ff",x"c0",x"1e"),
   378 => (x"f1",x"1e",x"d8",x"c1"),
   379 => (x"86",x"c8",x"87",x"e3"),
   380 => (x"c0",x"02",x"98",x"70"),
   381 => (x"d2",x"da",x"87",x"cd"),
   382 => (x"87",x"da",x"e9",x"1e"),
   383 => (x"48",x"c1",x"86",x"c4"),
   384 => (x"74",x"87",x"c5",x"c2"),
   385 => (x"7b",x"fe",x"c3",x"7b"),
   386 => (x"78",x"c0",x"48",x"76"),
   387 => (x"25",x"4d",x"66",x"d8"),
   388 => (x"d8",x"4a",x"71",x"49"),
   389 => (x"48",x"72",x"2a",x"b7"),
   390 => (x"7b",x"70",x"98",x"74"),
   391 => (x"b7",x"d0",x"4a",x"71"),
   392 => (x"74",x"48",x"72",x"2a"),
   393 => (x"71",x"7b",x"70",x"98"),
   394 => (x"2a",x"b7",x"c8",x"4a"),
   395 => (x"98",x"74",x"48",x"72"),
   396 => (x"48",x"71",x"7b",x"70"),
   397 => (x"7b",x"70",x"98",x"74"),
   398 => (x"80",x"c1",x"48",x"6e"),
   399 => (x"6e",x"58",x"a6",x"c4"),
   400 => (x"b7",x"c0",x"c2",x"48"),
   401 => (x"c6",x"ff",x"04",x"a8"),
   402 => (x"c0",x"c0",x"c8",x"87"),
   403 => (x"74",x"7b",x"74",x"4d"),
   404 => (x"d8",x"7b",x"74",x"7b"),
   405 => (x"74",x"49",x"e0",x"da"),
   406 => (x"c0",x"05",x"6b",x"7b"),
   407 => (x"89",x"c1",x"87",x"c6"),
   408 => (x"87",x"f3",x"ff",x"05"),
   409 => (x"d0",x"ff",x"7b",x"74"),
   410 => (x"98",x"75",x"48",x"bf"),
   411 => (x"6e",x"58",x"a6",x"c4"),
   412 => (x"87",x"ce",x"c0",x"02"),
   413 => (x"48",x"bf",x"d0",x"ff"),
   414 => (x"a6",x"c4",x"98",x"75"),
   415 => (x"ff",x"05",x"6e",x"58"),
   416 => (x"d0",x"ff",x"87",x"f2"),
   417 => (x"48",x"78",x"c0",x"48"),
   418 => (x"4d",x"26",x"8e",x"fc"),
   419 => (x"4b",x"26",x"4c",x"26"),
   420 => (x"72",x"57",x"4f",x"26"),
   421 => (x"20",x"65",x"74",x"69"),
   422 => (x"6c",x"69",x"61",x"66"),
   423 => (x"00",x"0a",x"64",x"65"),
   424 => (x"5c",x"5b",x"5e",x"0e"),
   425 => (x"d4",x"ff",x"0e",x"5d"),
   426 => (x"4c",x"66",x"d4",x"4d"),
   427 => (x"c0",x"4b",x"66",x"d0"),
   428 => (x"cd",x"ee",x"c5",x"4a"),
   429 => (x"ff",x"c3",x"49",x"df"),
   430 => (x"c3",x"48",x"6d",x"7d"),
   431 => (x"c1",x"05",x"a8",x"fe"),
   432 => (x"d1",x"c1",x"87",x"d4"),
   433 => (x"78",x"c0",x"48",x"fc"),
   434 => (x"04",x"ac",x"b7",x"c4"),
   435 => (x"eb",x"87",x"dc",x"c0"),
   436 => (x"49",x"70",x"87",x"fe"),
   437 => (x"83",x"c4",x"7b",x"71"),
   438 => (x"bf",x"fc",x"d1",x"c1"),
   439 => (x"c1",x"80",x"71",x"48"),
   440 => (x"c4",x"58",x"c0",x"d2"),
   441 => (x"03",x"ac",x"b7",x"8c"),
   442 => (x"c0",x"87",x"e4",x"ff"),
   443 => (x"c0",x"06",x"ac",x"b7"),
   444 => (x"ff",x"c3",x"87",x"e1"),
   445 => (x"71",x"49",x"6d",x"7d"),
   446 => (x"ff",x"c3",x"7b",x"97"),
   447 => (x"c1",x"83",x"c1",x"98"),
   448 => (x"48",x"bf",x"fc",x"d1"),
   449 => (x"d2",x"c1",x"80",x"71"),
   450 => (x"8c",x"c1",x"58",x"c0"),
   451 => (x"01",x"ac",x"b7",x"c0"),
   452 => (x"c1",x"87",x"df",x"ff"),
   453 => (x"89",x"c1",x"4a",x"49"),
   454 => (x"87",x"da",x"fe",x"05"),
   455 => (x"72",x"7d",x"ff",x"c3"),
   456 => (x"26",x"4d",x"26",x"48"),
   457 => (x"26",x"4b",x"26",x"4c"),
   458 => (x"5b",x"5e",x"0e",x"4f"),
   459 => (x"fc",x"0e",x"5d",x"5c"),
   460 => (x"4c",x"d0",x"ff",x"86"),
   461 => (x"4b",x"c0",x"c0",x"c8"),
   462 => (x"d4",x"ff",x"4d",x"c0"),
   463 => (x"78",x"ff",x"c3",x"48"),
   464 => (x"98",x"73",x"48",x"6c"),
   465 => (x"6e",x"58",x"a6",x"c4"),
   466 => (x"87",x"cc",x"c0",x"02"),
   467 => (x"98",x"73",x"48",x"6c"),
   468 => (x"6e",x"58",x"a6",x"c4"),
   469 => (x"87",x"f4",x"ff",x"05"),
   470 => (x"ff",x"7c",x"c1",x"c4"),
   471 => (x"ff",x"c3",x"48",x"d4"),
   472 => (x"1e",x"66",x"d4",x"78"),
   473 => (x"c1",x"f0",x"ff",x"c0"),
   474 => (x"e4",x"eb",x"1e",x"d1"),
   475 => (x"70",x"86",x"c8",x"87"),
   476 => (x"02",x"99",x"71",x"49"),
   477 => (x"71",x"87",x"d0",x"c0"),
   478 => (x"1e",x"66",x"d8",x"1e"),
   479 => (x"e4",x"1e",x"fa",x"de"),
   480 => (x"86",x"cc",x"87",x"c5"),
   481 => (x"c8",x"87",x"e7",x"c0"),
   482 => (x"66",x"dc",x"1e",x"c0"),
   483 => (x"87",x"d0",x"fc",x"1e"),
   484 => (x"4d",x"70",x"86",x"c8"),
   485 => (x"98",x"73",x"48",x"6c"),
   486 => (x"6e",x"58",x"a6",x"c4"),
   487 => (x"87",x"cc",x"c0",x"02"),
   488 => (x"98",x"73",x"48",x"6c"),
   489 => (x"6e",x"58",x"a6",x"c4"),
   490 => (x"87",x"f4",x"ff",x"05"),
   491 => (x"48",x"75",x"7c",x"c0"),
   492 => (x"4d",x"26",x"8e",x"fc"),
   493 => (x"4b",x"26",x"4c",x"26"),
   494 => (x"65",x"52",x"4f",x"26"),
   495 => (x"63",x"20",x"64",x"61"),
   496 => (x"61",x"6d",x"6d",x"6f"),
   497 => (x"66",x"20",x"64",x"6e"),
   498 => (x"65",x"6c",x"69",x"61"),
   499 => (x"74",x"61",x"20",x"64"),
   500 => (x"20",x"64",x"25",x"20"),
   501 => (x"29",x"64",x"25",x"28"),
   502 => (x"5e",x"0e",x"00",x"0a"),
   503 => (x"0e",x"5d",x"5c",x"5b"),
   504 => (x"1e",x"c0",x"86",x"fc"),
   505 => (x"c1",x"f0",x"ff",x"c0"),
   506 => (x"e4",x"e9",x"1e",x"c9"),
   507 => (x"d2",x"86",x"c8",x"87"),
   508 => (x"ce",x"d2",x"c1",x"1e"),
   509 => (x"87",x"e8",x"fa",x"1e"),
   510 => (x"4d",x"c0",x"86",x"c8"),
   511 => (x"b7",x"d2",x"85",x"c1"),
   512 => (x"f7",x"ff",x"04",x"ad"),
   513 => (x"ce",x"d2",x"c1",x"87"),
   514 => (x"c3",x"49",x"bf",x"97"),
   515 => (x"c0",x"c1",x"99",x"c0"),
   516 => (x"e8",x"c0",x"05",x"a9"),
   517 => (x"d5",x"d2",x"c1",x"87"),
   518 => (x"d0",x"49",x"bf",x"97"),
   519 => (x"d6",x"d2",x"c1",x"31"),
   520 => (x"c8",x"4a",x"bf",x"97"),
   521 => (x"c1",x"b1",x"72",x"32"),
   522 => (x"bf",x"97",x"d7",x"d2"),
   523 => (x"cf",x"b1",x"72",x"4a"),
   524 => (x"99",x"ff",x"ff",x"ff"),
   525 => (x"85",x"c1",x"4d",x"71"),
   526 => (x"eb",x"c2",x"35",x"ca"),
   527 => (x"d7",x"d2",x"c1",x"87"),
   528 => (x"c1",x"4b",x"bf",x"97"),
   529 => (x"c1",x"9b",x"c6",x"33"),
   530 => (x"bf",x"97",x"d8",x"d2"),
   531 => (x"29",x"b7",x"c7",x"49"),
   532 => (x"d2",x"c1",x"b3",x"71"),
   533 => (x"49",x"bf",x"97",x"d3"),
   534 => (x"98",x"cf",x"48",x"71"),
   535 => (x"c1",x"58",x"a6",x"c4"),
   536 => (x"bf",x"97",x"d4",x"d2"),
   537 => (x"ca",x"9c",x"c3",x"4c"),
   538 => (x"d5",x"d2",x"c1",x"34"),
   539 => (x"c2",x"49",x"bf",x"97"),
   540 => (x"c1",x"b4",x"71",x"31"),
   541 => (x"bf",x"97",x"d6",x"d2"),
   542 => (x"99",x"c0",x"c3",x"49"),
   543 => (x"71",x"29",x"b7",x"c6"),
   544 => (x"c4",x"1e",x"74",x"b4"),
   545 => (x"1e",x"73",x"1e",x"66"),
   546 => (x"1e",x"f4",x"e3",x"c0"),
   547 => (x"87",x"f7",x"df",x"ff"),
   548 => (x"83",x"c2",x"86",x"d0"),
   549 => (x"30",x"73",x"48",x"c1"),
   550 => (x"1e",x"73",x"4b",x"70"),
   551 => (x"1e",x"e1",x"e4",x"c0"),
   552 => (x"87",x"e3",x"df",x"ff"),
   553 => (x"48",x"c1",x"86",x"c8"),
   554 => (x"a6",x"c4",x"30",x"6e"),
   555 => (x"c1",x"49",x"74",x"58"),
   556 => (x"73",x"4d",x"71",x"81"),
   557 => (x"1e",x"6e",x"95",x"b7"),
   558 => (x"e4",x"c0",x"1e",x"75"),
   559 => (x"df",x"ff",x"1e",x"ea"),
   560 => (x"86",x"cc",x"87",x"c5"),
   561 => (x"c0",x"c8",x"48",x"6e"),
   562 => (x"c0",x"06",x"a8",x"b7"),
   563 => (x"4b",x"6e",x"87",x"ce"),
   564 => (x"2b",x"b7",x"35",x"c1"),
   565 => (x"ab",x"b7",x"c0",x"c8"),
   566 => (x"87",x"f4",x"ff",x"01"),
   567 => (x"e5",x"c0",x"1e",x"75"),
   568 => (x"de",x"ff",x"1e",x"c0"),
   569 => (x"86",x"c8",x"87",x"e1"),
   570 => (x"8e",x"fc",x"48",x"75"),
   571 => (x"4c",x"26",x"4d",x"26"),
   572 => (x"4f",x"26",x"4b",x"26"),
   573 => (x"69",x"73",x"5f",x"63"),
   574 => (x"6d",x"5f",x"65",x"7a"),
   575 => (x"3a",x"74",x"6c",x"75"),
   576 => (x"2c",x"64",x"25",x"20"),
   577 => (x"61",x"65",x"72",x"20"),
   578 => (x"6c",x"62",x"5f",x"64"),
   579 => (x"6e",x"65",x"6c",x"5f"),
   580 => (x"64",x"25",x"20",x"3a"),
   581 => (x"73",x"63",x"20",x"2c"),
   582 => (x"3a",x"65",x"7a",x"69"),
   583 => (x"0a",x"64",x"25",x"20"),
   584 => (x"6c",x"75",x"4d",x"00"),
   585 => (x"64",x"25",x"20",x"74"),
   586 => (x"64",x"25",x"00",x"0a"),
   587 => (x"6f",x"6c",x"62",x"20"),
   588 => (x"20",x"73",x"6b",x"63"),
   589 => (x"73",x"20",x"66",x"6f"),
   590 => (x"20",x"65",x"7a",x"69"),
   591 => (x"00",x"0a",x"64",x"25"),
   592 => (x"62",x"20",x"64",x"25"),
   593 => (x"6b",x"63",x"6f",x"6c"),
   594 => (x"66",x"6f",x"20",x"73"),
   595 => (x"32",x"31",x"35",x"20"),
   596 => (x"74",x"79",x"62",x"20"),
   597 => (x"00",x"0a",x"73",x"65"),
   598 => (x"00",x"44",x"4d",x"43"),
   599 => (x"0e",x"5b",x"5e",x"0e"),
   600 => (x"66",x"d0",x"4b",x"c0"),
   601 => (x"a8",x"b7",x"c0",x"48"),
   602 => (x"87",x"f6",x"c0",x"06"),
   603 => (x"bf",x"97",x"66",x"c8"),
   604 => (x"82",x"c0",x"fe",x"4a"),
   605 => (x"48",x"66",x"c8",x"ba"),
   606 => (x"a6",x"cc",x"80",x"c1"),
   607 => (x"97",x"66",x"cc",x"58"),
   608 => (x"c0",x"fe",x"49",x"bf"),
   609 => (x"66",x"cc",x"b9",x"81"),
   610 => (x"d0",x"80",x"c1",x"48"),
   611 => (x"b7",x"71",x"58",x"a6"),
   612 => (x"87",x"c4",x"02",x"aa"),
   613 => (x"87",x"cc",x"48",x"c1"),
   614 => (x"66",x"d0",x"83",x"c1"),
   615 => (x"ff",x"04",x"ab",x"b7"),
   616 => (x"48",x"c0",x"87",x"ca"),
   617 => (x"4d",x"26",x"87",x"c4"),
   618 => (x"4b",x"26",x"4c",x"26"),
   619 => (x"5e",x"0e",x"4f",x"26"),
   620 => (x"0e",x"5d",x"5c",x"5b"),
   621 => (x"48",x"e8",x"da",x"c1"),
   622 => (x"f6",x"c0",x"78",x"c0"),
   623 => (x"da",x"ff",x"1e",x"d0"),
   624 => (x"86",x"c4",x"87",x"d4"),
   625 => (x"1e",x"e0",x"d2",x"c1"),
   626 => (x"dc",x"f5",x"1e",x"c0"),
   627 => (x"70",x"86",x"c8",x"87"),
   628 => (x"87",x"cf",x"05",x"98"),
   629 => (x"1e",x"fc",x"f2",x"c0"),
   630 => (x"87",x"fa",x"d9",x"ff"),
   631 => (x"48",x"c0",x"86",x"c4"),
   632 => (x"c0",x"87",x"d6",x"cb"),
   633 => (x"ff",x"1e",x"dd",x"f6"),
   634 => (x"c4",x"87",x"eb",x"d9"),
   635 => (x"c1",x"4b",x"c0",x"86"),
   636 => (x"c1",x"48",x"d4",x"db"),
   637 => (x"c0",x"1e",x"c8",x"78"),
   638 => (x"c1",x"1e",x"f4",x"f6"),
   639 => (x"fd",x"1e",x"d6",x"d3"),
   640 => (x"86",x"cc",x"87",x"da"),
   641 => (x"c6",x"05",x"98",x"70"),
   642 => (x"d4",x"db",x"c1",x"87"),
   643 => (x"c8",x"78",x"c0",x"48"),
   644 => (x"fd",x"f6",x"c0",x"1e"),
   645 => (x"f2",x"d3",x"c1",x"1e"),
   646 => (x"87",x"c0",x"fd",x"1e"),
   647 => (x"98",x"70",x"86",x"cc"),
   648 => (x"c1",x"87",x"c6",x"05"),
   649 => (x"c0",x"48",x"d4",x"db"),
   650 => (x"d4",x"db",x"c1",x"78"),
   651 => (x"f7",x"c0",x"1e",x"bf"),
   652 => (x"d9",x"ff",x"1e",x"c6"),
   653 => (x"86",x"c8",x"87",x"d1"),
   654 => (x"bf",x"d4",x"db",x"c1"),
   655 => (x"87",x"d8",x"c2",x"02"),
   656 => (x"4d",x"e0",x"d2",x"c1"),
   657 => (x"4c",x"de",x"d9",x"c1"),
   658 => (x"9f",x"de",x"da",x"c1"),
   659 => (x"1e",x"71",x"49",x"bf"),
   660 => (x"49",x"de",x"da",x"c1"),
   661 => (x"89",x"e0",x"d2",x"c1"),
   662 => (x"1e",x"d0",x"1e",x"71"),
   663 => (x"c0",x"1e",x"c0",x"c8"),
   664 => (x"ff",x"1e",x"ee",x"f3"),
   665 => (x"d4",x"87",x"e0",x"d8"),
   666 => (x"c8",x"49",x"74",x"86"),
   667 => (x"c1",x"4b",x"69",x"81"),
   668 => (x"bf",x"9f",x"de",x"da"),
   669 => (x"ea",x"d6",x"c5",x"49"),
   670 => (x"d0",x"c0",x"05",x"a9"),
   671 => (x"c8",x"49",x"74",x"87"),
   672 => (x"d9",x"1e",x"69",x"81"),
   673 => (x"86",x"c4",x"87",x"c2"),
   674 => (x"df",x"c0",x"4b",x"70"),
   675 => (x"c7",x"49",x"75",x"87"),
   676 => (x"69",x"9f",x"81",x"fe"),
   677 => (x"d5",x"e9",x"ca",x"49"),
   678 => (x"cf",x"c0",x"02",x"a9"),
   679 => (x"d0",x"f3",x"c0",x"87"),
   680 => (x"f1",x"d6",x"ff",x"1e"),
   681 => (x"c0",x"86",x"c4",x"87"),
   682 => (x"87",x"cd",x"c8",x"48"),
   683 => (x"f4",x"c0",x"1e",x"73"),
   684 => (x"d7",x"ff",x"1e",x"eb"),
   685 => (x"86",x"c8",x"87",x"d1"),
   686 => (x"1e",x"e0",x"d2",x"c1"),
   687 => (x"e8",x"f1",x"1e",x"73"),
   688 => (x"70",x"86",x"c8",x"87"),
   689 => (x"c5",x"c0",x"05",x"98"),
   690 => (x"c7",x"48",x"c0",x"87"),
   691 => (x"f5",x"c0",x"87",x"eb"),
   692 => (x"d6",x"ff",x"1e",x"c3"),
   693 => (x"86",x"c4",x"87",x"c0"),
   694 => (x"1e",x"d9",x"f7",x"c0"),
   695 => (x"87",x"e7",x"d6",x"ff"),
   696 => (x"1e",x"c8",x"86",x"c4"),
   697 => (x"1e",x"f1",x"f7",x"c0"),
   698 => (x"1e",x"f2",x"d3",x"c1"),
   699 => (x"cc",x"87",x"ed",x"f9"),
   700 => (x"05",x"98",x"70",x"86"),
   701 => (x"c1",x"87",x"c9",x"c0"),
   702 => (x"c1",x"48",x"e8",x"da"),
   703 => (x"87",x"e4",x"c0",x"78"),
   704 => (x"f7",x"c0",x"1e",x"c8"),
   705 => (x"d3",x"c1",x"1e",x"fa"),
   706 => (x"cf",x"f9",x"1e",x"d6"),
   707 => (x"70",x"86",x"cc",x"87"),
   708 => (x"cf",x"c0",x"02",x"98"),
   709 => (x"ea",x"f5",x"c0",x"87"),
   710 => (x"ea",x"d5",x"ff",x"1e"),
   711 => (x"c0",x"86",x"c4",x"87"),
   712 => (x"87",x"d5",x"c6",x"48"),
   713 => (x"97",x"de",x"da",x"c1"),
   714 => (x"d5",x"c1",x"49",x"bf"),
   715 => (x"cd",x"c0",x"05",x"a9"),
   716 => (x"df",x"da",x"c1",x"87"),
   717 => (x"c2",x"49",x"bf",x"97"),
   718 => (x"c0",x"02",x"a9",x"ea"),
   719 => (x"48",x"c0",x"87",x"c5"),
   720 => (x"c1",x"87",x"f6",x"c5"),
   721 => (x"bf",x"97",x"e0",x"d2"),
   722 => (x"a9",x"e9",x"c3",x"49"),
   723 => (x"87",x"d2",x"c0",x"02"),
   724 => (x"97",x"e0",x"d2",x"c1"),
   725 => (x"eb",x"c3",x"49",x"bf"),
   726 => (x"c5",x"c0",x"02",x"a9"),
   727 => (x"c5",x"48",x"c0",x"87"),
   728 => (x"d2",x"c1",x"87",x"d7"),
   729 => (x"49",x"bf",x"97",x"eb"),
   730 => (x"c0",x"05",x"99",x"71"),
   731 => (x"d2",x"c1",x"87",x"cc"),
   732 => (x"49",x"bf",x"97",x"ec"),
   733 => (x"c0",x"02",x"a9",x"c2"),
   734 => (x"48",x"c0",x"87",x"c5"),
   735 => (x"c1",x"87",x"fa",x"c4"),
   736 => (x"bf",x"97",x"ed",x"d2"),
   737 => (x"e4",x"da",x"c1",x"48"),
   738 => (x"e0",x"da",x"c1",x"58"),
   739 => (x"4a",x"71",x"49",x"bf"),
   740 => (x"da",x"c1",x"8a",x"c1"),
   741 => (x"1e",x"72",x"5a",x"e8"),
   742 => (x"f8",x"c0",x"1e",x"71"),
   743 => (x"d3",x"ff",x"1e",x"c3"),
   744 => (x"86",x"cc",x"87",x"e5"),
   745 => (x"97",x"ee",x"d2",x"c1"),
   746 => (x"81",x"73",x"49",x"bf"),
   747 => (x"97",x"ef",x"d2",x"c1"),
   748 => (x"32",x"c8",x"4a",x"bf"),
   749 => (x"80",x"71",x"48",x"72"),
   750 => (x"58",x"f8",x"da",x"c1"),
   751 => (x"97",x"f0",x"d2",x"c1"),
   752 => (x"db",x"c1",x"48",x"bf"),
   753 => (x"da",x"c1",x"58",x"cc"),
   754 => (x"c2",x"02",x"bf",x"e8"),
   755 => (x"1e",x"c8",x"87",x"da"),
   756 => (x"1e",x"c7",x"f6",x"c0"),
   757 => (x"1e",x"f2",x"d3",x"c1"),
   758 => (x"cc",x"87",x"c1",x"f6"),
   759 => (x"02",x"98",x"70",x"86"),
   760 => (x"c0",x"87",x"c5",x"c0"),
   761 => (x"87",x"d1",x"c3",x"48"),
   762 => (x"bf",x"e0",x"da",x"c1"),
   763 => (x"c4",x"48",x"72",x"4a"),
   764 => (x"d0",x"db",x"c1",x"30"),
   765 => (x"c8",x"db",x"c1",x"58"),
   766 => (x"c5",x"d3",x"c1",x"5a"),
   767 => (x"c8",x"49",x"bf",x"97"),
   768 => (x"c4",x"d3",x"c1",x"31"),
   769 => (x"73",x"4b",x"bf",x"97"),
   770 => (x"c6",x"d3",x"c1",x"81"),
   771 => (x"d0",x"4b",x"bf",x"97"),
   772 => (x"c1",x"81",x"73",x"33"),
   773 => (x"bf",x"97",x"c7",x"d3"),
   774 => (x"73",x"33",x"d8",x"4b"),
   775 => (x"d4",x"db",x"c1",x"81"),
   776 => (x"c8",x"db",x"c1",x"59"),
   777 => (x"da",x"c1",x"91",x"bf"),
   778 => (x"c1",x"81",x"bf",x"f4"),
   779 => (x"c1",x"59",x"fc",x"da"),
   780 => (x"bf",x"97",x"cd",x"d3"),
   781 => (x"c1",x"33",x"c8",x"4b"),
   782 => (x"bf",x"97",x"cc",x"d3"),
   783 => (x"c1",x"83",x"74",x"4c"),
   784 => (x"bf",x"97",x"ce",x"d3"),
   785 => (x"74",x"34",x"d0",x"4c"),
   786 => (x"cf",x"d3",x"c1",x"83"),
   787 => (x"cf",x"4c",x"bf",x"97"),
   788 => (x"74",x"34",x"d8",x"9c"),
   789 => (x"c0",x"db",x"c1",x"83"),
   790 => (x"73",x"8b",x"c2",x"5b"),
   791 => (x"71",x"48",x"72",x"92"),
   792 => (x"c4",x"db",x"c1",x"80"),
   793 => (x"87",x"cf",x"c1",x"58"),
   794 => (x"97",x"f2",x"d2",x"c1"),
   795 => (x"31",x"c8",x"49",x"bf"),
   796 => (x"97",x"f1",x"d2",x"c1"),
   797 => (x"81",x"72",x"4a",x"bf"),
   798 => (x"59",x"d0",x"db",x"c1"),
   799 => (x"ff",x"c7",x"31",x"c5"),
   800 => (x"c1",x"29",x"c9",x"81"),
   801 => (x"c1",x"59",x"c8",x"db"),
   802 => (x"bf",x"97",x"f7",x"d2"),
   803 => (x"c1",x"32",x"c8",x"4a"),
   804 => (x"bf",x"97",x"f6",x"d2"),
   805 => (x"c1",x"82",x"73",x"4b"),
   806 => (x"c1",x"5a",x"d4",x"db"),
   807 => (x"92",x"bf",x"c8",x"db"),
   808 => (x"bf",x"f4",x"da",x"c1"),
   809 => (x"c4",x"db",x"c1",x"82"),
   810 => (x"fc",x"da",x"c1",x"5a"),
   811 => (x"72",x"78",x"c0",x"48"),
   812 => (x"c1",x"80",x"71",x"48"),
   813 => (x"c1",x"58",x"fc",x"da"),
   814 => (x"87",x"ea",x"f3",x"48"),
   815 => (x"64",x"61",x"65",x"52"),
   816 => (x"20",x"66",x"6f",x"20"),
   817 => (x"20",x"52",x"42",x"4d"),
   818 => (x"6c",x"69",x"61",x"66"),
   819 => (x"00",x"0a",x"64",x"65"),
   820 => (x"70",x"20",x"6f",x"4e"),
   821 => (x"69",x"74",x"72",x"61"),
   822 => (x"6e",x"6f",x"69",x"74"),
   823 => (x"67",x"69",x"73",x"20"),
   824 => (x"75",x"74",x"61",x"6e"),
   825 => (x"66",x"20",x"65",x"72"),
   826 => (x"64",x"6e",x"75",x"6f"),
   827 => (x"42",x"4d",x"00",x"0a"),
   828 => (x"7a",x"69",x"73",x"52"),
   829 => (x"25",x"20",x"3a",x"65"),
   830 => (x"70",x"20",x"2c",x"64"),
   831 => (x"69",x"74",x"72",x"61"),
   832 => (x"6e",x"6f",x"69",x"74"),
   833 => (x"65",x"7a",x"69",x"73"),
   834 => (x"64",x"25",x"20",x"3a"),
   835 => (x"66",x"6f",x"20",x"2c"),
   836 => (x"74",x"65",x"73",x"66"),
   837 => (x"20",x"66",x"6f",x"20"),
   838 => (x"3a",x"67",x"69",x"73"),
   839 => (x"2c",x"64",x"25",x"20"),
   840 => (x"67",x"69",x"73",x"20"),
   841 => (x"25",x"78",x"30",x"20"),
   842 => (x"52",x"00",x"0a",x"78"),
   843 => (x"69",x"64",x"61",x"65"),
   844 => (x"62",x"20",x"67",x"6e"),
   845 => (x"20",x"74",x"6f",x"6f"),
   846 => (x"74",x"63",x"65",x"73"),
   847 => (x"25",x"20",x"72",x"6f"),
   848 => (x"52",x"00",x"0a",x"64"),
   849 => (x"20",x"64",x"61",x"65"),
   850 => (x"74",x"6f",x"6f",x"62"),
   851 => (x"63",x"65",x"73",x"20"),
   852 => (x"20",x"72",x"6f",x"74"),
   853 => (x"6d",x"6f",x"72",x"66"),
   854 => (x"72",x"69",x"66",x"20"),
   855 => (x"70",x"20",x"74",x"73"),
   856 => (x"69",x"74",x"72",x"61"),
   857 => (x"6e",x"6f",x"69",x"74"),
   858 => (x"6e",x"55",x"00",x"0a"),
   859 => (x"70",x"70",x"75",x"73"),
   860 => (x"65",x"74",x"72",x"6f"),
   861 => (x"61",x"70",x"20",x"64"),
   862 => (x"74",x"69",x"74",x"72"),
   863 => (x"20",x"6e",x"6f",x"69"),
   864 => (x"65",x"70",x"79",x"74"),
   865 => (x"46",x"00",x"0d",x"21"),
   866 => (x"32",x"33",x"54",x"41"),
   867 => (x"00",x"20",x"20",x"20"),
   868 => (x"64",x"61",x"65",x"52"),
   869 => (x"20",x"67",x"6e",x"69"),
   870 => (x"0a",x"52",x"42",x"4d"),
   871 => (x"52",x"42",x"4d",x"00"),
   872 => (x"63",x"75",x"73",x"20"),
   873 => (x"73",x"73",x"65",x"63"),
   874 => (x"6c",x"6c",x"75",x"66"),
   875 => (x"65",x"72",x"20",x"79"),
   876 => (x"00",x"0a",x"64",x"61"),
   877 => (x"31",x"54",x"41",x"46"),
   878 => (x"20",x"20",x"20",x"36"),
   879 => (x"54",x"41",x"46",x"00"),
   880 => (x"20",x"20",x"32",x"33"),
   881 => (x"61",x"50",x"00",x"20"),
   882 => (x"74",x"69",x"74",x"72"),
   883 => (x"63",x"6e",x"6f",x"69"),
   884 => (x"74",x"6e",x"75",x"6f"),
   885 => (x"0a",x"64",x"25",x"20"),
   886 => (x"6e",x"75",x"48",x"00"),
   887 => (x"67",x"6e",x"69",x"74"),
   888 => (x"72",x"6f",x"66",x"20"),
   889 => (x"6c",x"69",x"66",x"20"),
   890 => (x"73",x"79",x"73",x"65"),
   891 => (x"0a",x"6d",x"65",x"74"),
   892 => (x"54",x"41",x"46",x"00"),
   893 => (x"20",x"20",x"32",x"33"),
   894 => (x"41",x"46",x"00",x"20"),
   895 => (x"20",x"36",x"31",x"54"),
   896 => (x"43",x"00",x"20",x"20"),
   897 => (x"74",x"73",x"75",x"6c"),
   898 => (x"73",x"20",x"72",x"65"),
   899 => (x"3a",x"65",x"7a",x"69"),
   900 => (x"2c",x"64",x"25",x"20"),
   901 => (x"75",x"6c",x"43",x"20"),
   902 => (x"72",x"65",x"74",x"73"),
   903 => (x"73",x"61",x"6d",x"20"),
   904 => (x"25",x"20",x"2c",x"6b"),
   905 => (x"0e",x"00",x"0a",x"64"),
   906 => (x"0e",x"5c",x"5b",x"5e"),
   907 => (x"bf",x"e8",x"da",x"c1"),
   908 => (x"cc",x"87",x"ce",x"02"),
   909 => (x"b7",x"c7",x"4a",x"66"),
   910 => (x"4b",x"66",x"cc",x"2a"),
   911 => (x"cc",x"9b",x"ff",x"c1"),
   912 => (x"4a",x"66",x"cc",x"87"),
   913 => (x"cc",x"2a",x"b7",x"c8"),
   914 => (x"ff",x"c3",x"4b",x"66"),
   915 => (x"e0",x"d2",x"c1",x"9b"),
   916 => (x"f4",x"da",x"c1",x"1e"),
   917 => (x"81",x"72",x"49",x"bf"),
   918 => (x"cc",x"e3",x"1e",x"71"),
   919 => (x"70",x"86",x"c8",x"87"),
   920 => (x"87",x"c5",x"05",x"98"),
   921 => (x"e8",x"c0",x"48",x"c0"),
   922 => (x"e8",x"da",x"c1",x"87"),
   923 => (x"87",x"d3",x"02",x"bf"),
   924 => (x"b7",x"c4",x"49",x"73"),
   925 => (x"e0",x"d2",x"c1",x"91"),
   926 => (x"cf",x"4c",x"69",x"81"),
   927 => (x"ff",x"ff",x"ff",x"ff"),
   928 => (x"73",x"87",x"cc",x"9c"),
   929 => (x"91",x"b7",x"c2",x"49"),
   930 => (x"81",x"e0",x"d2",x"c1"),
   931 => (x"74",x"4c",x"69",x"9f"),
   932 => (x"87",x"d4",x"ec",x"48"),
   933 => (x"5c",x"5b",x"5e",x"0e"),
   934 => (x"86",x"f4",x"0e",x"5d"),
   935 => (x"48",x"76",x"4b",x"c0"),
   936 => (x"bf",x"fc",x"da",x"c1"),
   937 => (x"c1",x"80",x"c4",x"78"),
   938 => (x"78",x"bf",x"c0",x"db"),
   939 => (x"bf",x"e8",x"da",x"c1"),
   940 => (x"c1",x"87",x"c9",x"02"),
   941 => (x"49",x"bf",x"e0",x"da"),
   942 => (x"87",x"c7",x"31",x"c4"),
   943 => (x"bf",x"c4",x"db",x"c1"),
   944 => (x"cc",x"31",x"c4",x"49"),
   945 => (x"4d",x"c0",x"59",x"a6"),
   946 => (x"c0",x"48",x"66",x"c8"),
   947 => (x"ed",x"c2",x"06",x"a8"),
   948 => (x"cf",x"49",x"75",x"87"),
   949 => (x"87",x"da",x"05",x"99"),
   950 => (x"1e",x"e0",x"d2",x"c1"),
   951 => (x"48",x"49",x"66",x"c8"),
   952 => (x"a6",x"cc",x"80",x"c1"),
   953 => (x"e0",x"1e",x"71",x"58"),
   954 => (x"86",x"c8",x"87",x"ff"),
   955 => (x"4b",x"e0",x"d2",x"c1"),
   956 => (x"e0",x"c0",x"87",x"c3"),
   957 => (x"49",x"6b",x"97",x"83"),
   958 => (x"c1",x"02",x"99",x"71"),
   959 => (x"6b",x"97",x"87",x"f7"),
   960 => (x"a9",x"e5",x"c3",x"49"),
   961 => (x"87",x"ed",x"c1",x"02"),
   962 => (x"81",x"cb",x"49",x"73"),
   963 => (x"d8",x"49",x"69",x"97"),
   964 => (x"e0",x"c1",x"05",x"99"),
   965 => (x"ff",x"1e",x"73",x"87"),
   966 => (x"c4",x"87",x"fb",x"c4"),
   967 => (x"c0",x"1e",x"cb",x"86"),
   968 => (x"73",x"1e",x"66",x"e4"),
   969 => (x"87",x"f4",x"e8",x"1e"),
   970 => (x"98",x"70",x"86",x"cc"),
   971 => (x"87",x"c5",x"c1",x"05"),
   972 => (x"82",x"dc",x"4a",x"73"),
   973 => (x"c4",x"49",x"66",x"dc"),
   974 => (x"73",x"79",x"6a",x"81"),
   975 => (x"dc",x"82",x"da",x"4a"),
   976 => (x"81",x"c8",x"49",x"66"),
   977 => (x"70",x"48",x"6a",x"9f"),
   978 => (x"c1",x"4c",x"71",x"79"),
   979 => (x"02",x"bf",x"e8",x"da"),
   980 => (x"49",x"73",x"87",x"d1"),
   981 => (x"69",x"9f",x"81",x"d4"),
   982 => (x"ff",x"ff",x"c0",x"49"),
   983 => (x"d0",x"4a",x"71",x"99"),
   984 => (x"c0",x"87",x"c2",x"32"),
   985 => (x"6c",x"48",x"72",x"4a"),
   986 => (x"dc",x"7c",x"70",x"80"),
   987 => (x"78",x"c0",x"48",x"66"),
   988 => (x"ff",x"c0",x"48",x"c1"),
   989 => (x"c8",x"85",x"c1",x"87"),
   990 => (x"fd",x"04",x"ad",x"66"),
   991 => (x"da",x"c1",x"87",x"d3"),
   992 => (x"c0",x"02",x"bf",x"e8"),
   993 => (x"1e",x"6e",x"87",x"ec"),
   994 => (x"c4",x"87",x"dc",x"fa"),
   995 => (x"58",x"a6",x"c4",x"86"),
   996 => (x"ff",x"cf",x"49",x"6e"),
   997 => (x"99",x"f8",x"ff",x"ff"),
   998 => (x"87",x"d6",x"02",x"a9"),
   999 => (x"89",x"c2",x"49",x"6e"),
  1000 => (x"bf",x"e0",x"da",x"c1"),
  1001 => (x"f8",x"da",x"c1",x"91"),
  1002 => (x"80",x"71",x"48",x"bf"),
  1003 => (x"fc",x"58",x"a6",x"c8"),
  1004 => (x"48",x"c0",x"87",x"d4"),
  1005 => (x"ed",x"e7",x"8e",x"f4"),
  1006 => (x"5b",x"5e",x"0e",x"87"),
  1007 => (x"bf",x"66",x"c8",x"0e"),
  1008 => (x"c8",x"81",x"c1",x"49"),
  1009 => (x"09",x"79",x"09",x"66"),
  1010 => (x"bf",x"e4",x"da",x"c1"),
  1011 => (x"87",x"d0",x"05",x"99"),
  1012 => (x"c8",x"4b",x"66",x"c8"),
  1013 => (x"f9",x"1e",x"6b",x"83"),
  1014 => (x"86",x"c4",x"87",x"cd"),
  1015 => (x"7b",x"71",x"49",x"70"),
  1016 => (x"c5",x"e7",x"48",x"c1"),
  1017 => (x"0e",x"5e",x"0e",x"87"),
  1018 => (x"bf",x"f8",x"da",x"c1"),
  1019 => (x"4a",x"66",x"c4",x"49"),
  1020 => (x"4a",x"6a",x"82",x"c8"),
  1021 => (x"da",x"c1",x"8a",x"c2"),
  1022 => (x"72",x"92",x"bf",x"e0"),
  1023 => (x"e4",x"da",x"c1",x"81"),
  1024 => (x"66",x"c4",x"4a",x"bf"),
  1025 => (x"81",x"72",x"9a",x"bf"),
  1026 => (x"71",x"1e",x"66",x"c8"),
  1027 => (x"d8",x"dc",x"ff",x"1e"),
  1028 => (x"70",x"86",x"c8",x"87"),
  1029 => (x"87",x"c4",x"05",x"98"),
  1030 => (x"87",x"c2",x"48",x"c0"),
  1031 => (x"cb",x"e6",x"48",x"c1"),
  1032 => (x"5b",x"5e",x"0e",x"87"),
  1033 => (x"66",x"cc",x"0e",x"5c"),
  1034 => (x"d8",x"db",x"c1",x"1e"),
  1035 => (x"87",x"e4",x"f9",x"1e"),
  1036 => (x"98",x"70",x"86",x"c8"),
  1037 => (x"87",x"d2",x"c1",x"02"),
  1038 => (x"bf",x"dc",x"db",x"c1"),
  1039 => (x"81",x"ff",x"c7",x"49"),
  1040 => (x"4c",x"71",x"29",x"c9"),
  1041 => (x"c2",x"c1",x"4b",x"c0"),
  1042 => (x"c0",x"ff",x"1e",x"e0"),
  1043 => (x"86",x"c4",x"87",x"c8"),
  1044 => (x"06",x"ac",x"b7",x"c0"),
  1045 => (x"d0",x"87",x"c4",x"c1"),
  1046 => (x"db",x"c1",x"1e",x"66"),
  1047 => (x"c4",x"fe",x"1e",x"d8"),
  1048 => (x"70",x"86",x"c8",x"87"),
  1049 => (x"87",x"c5",x"05",x"98"),
  1050 => (x"f0",x"c0",x"48",x"c0"),
  1051 => (x"d8",x"db",x"c1",x"87"),
  1052 => (x"87",x"c5",x"fd",x"1e"),
  1053 => (x"66",x"d0",x"86",x"c4"),
  1054 => (x"80",x"c0",x"c8",x"48"),
  1055 => (x"c1",x"58",x"a6",x"d4"),
  1056 => (x"ab",x"b7",x"74",x"83"),
  1057 => (x"87",x"cf",x"ff",x"04"),
  1058 => (x"66",x"cc",x"87",x"d1"),
  1059 => (x"f9",x"c2",x"c1",x"1e"),
  1060 => (x"f2",x"ff",x"fe",x"1e"),
  1061 => (x"c0",x"86",x"c8",x"87"),
  1062 => (x"c1",x"87",x"c2",x"48"),
  1063 => (x"87",x"c8",x"e4",x"48"),
  1064 => (x"6e",x"65",x"70",x"4f"),
  1065 => (x"66",x"20",x"64",x"65"),
  1066 => (x"2c",x"65",x"6c",x"69"),
  1067 => (x"61",x"6f",x"6c",x"20"),
  1068 => (x"67",x"6e",x"69",x"64"),
  1069 => (x"0a",x"2e",x"2e",x"2e"),
  1070 => (x"6e",x"61",x"43",x"00"),
  1071 => (x"6f",x"20",x"74",x"27"),
  1072 => (x"20",x"6e",x"65",x"70"),
  1073 => (x"00",x"0a",x"73",x"25"),
  1074 => (x"c4",x"0e",x"5e",x"0e"),
  1075 => (x"29",x"d8",x"49",x"66"),
  1076 => (x"c4",x"99",x"ff",x"c3"),
  1077 => (x"2a",x"c8",x"4a",x"66"),
  1078 => (x"9a",x"c0",x"fc",x"cf"),
  1079 => (x"66",x"c4",x"b1",x"72"),
  1080 => (x"c0",x"32",x"c8",x"4a"),
  1081 => (x"c0",x"c0",x"f0",x"ff"),
  1082 => (x"c4",x"b1",x"72",x"9a"),
  1083 => (x"32",x"d8",x"4a",x"66"),
  1084 => (x"c0",x"c0",x"c0",x"ff"),
  1085 => (x"b1",x"72",x"9a",x"c0"),
  1086 => (x"87",x"c6",x"48",x"71"),
  1087 => (x"4c",x"26",x"4d",x"26"),
  1088 => (x"4f",x"26",x"4b",x"26"),
  1089 => (x"d0",x"1e",x"73",x"1e"),
  1090 => (x"c0",x"c0",x"c0",x"c0"),
  1091 => (x"fe",x"0f",x"73",x"4b"),
  1092 => (x"26",x"87",x"c4",x"87"),
  1093 => (x"26",x"4c",x"26",x"4d"),
  1094 => (x"1e",x"4f",x"26",x"4b"),
  1095 => (x"c3",x"49",x"66",x"c8"),
  1096 => (x"f7",x"c0",x"99",x"df"),
  1097 => (x"a9",x"b7",x"c0",x"89"),
  1098 => (x"c0",x"87",x"c3",x"03"),
  1099 => (x"66",x"c4",x"81",x"e7"),
  1100 => (x"c8",x"30",x"c4",x"48"),
  1101 => (x"66",x"c4",x"58",x"a6"),
  1102 => (x"c8",x"b0",x"71",x"48"),
  1103 => (x"66",x"c4",x"58",x"a6"),
  1104 => (x"87",x"d5",x"ff",x"48"),
  1105 => (x"5c",x"5b",x"5e",x"0e"),
  1106 => (x"c0",x"c0",x"d0",x"0e"),
  1107 => (x"c1",x"4c",x"c0",x"c0"),
  1108 => (x"48",x"bf",x"e4",x"db"),
  1109 => (x"db",x"c1",x"80",x"c1"),
  1110 => (x"cc",x"97",x"58",x"e8"),
  1111 => (x"c0",x"fe",x"49",x"66"),
  1112 => (x"d3",x"c1",x"b9",x"81"),
  1113 => (x"87",x"db",x"05",x"a9"),
  1114 => (x"48",x"e4",x"db",x"c1"),
  1115 => (x"db",x"c1",x"78",x"c0"),
  1116 => (x"78",x"c0",x"48",x"e8"),
  1117 => (x"48",x"f0",x"db",x"c1"),
  1118 => (x"db",x"c1",x"78",x"c0"),
  1119 => (x"78",x"c0",x"48",x"f4"),
  1120 => (x"c1",x"87",x"fb",x"c6"),
  1121 => (x"48",x"bf",x"e4",x"db"),
  1122 => (x"c0",x"05",x"a8",x"c1"),
  1123 => (x"cc",x"97",x"87",x"f8"),
  1124 => (x"c0",x"fe",x"49",x"66"),
  1125 => (x"1e",x"71",x"b9",x"81"),
  1126 => (x"bf",x"f4",x"db",x"c1"),
  1127 => (x"87",x"fb",x"fd",x"1e"),
  1128 => (x"db",x"c1",x"86",x"c8"),
  1129 => (x"db",x"c1",x"58",x"f8"),
  1130 => (x"c3",x"4a",x"bf",x"f4"),
  1131 => (x"c6",x"06",x"aa",x"b7"),
  1132 => (x"72",x"48",x"ca",x"87"),
  1133 => (x"72",x"4a",x"70",x"88"),
  1134 => (x"71",x"81",x"c1",x"49"),
  1135 => (x"c1",x"30",x"c1",x"48"),
  1136 => (x"c5",x"58",x"f0",x"db"),
  1137 => (x"db",x"c1",x"87",x"f8"),
  1138 => (x"c9",x"48",x"bf",x"f4"),
  1139 => (x"c5",x"01",x"a8",x"b7"),
  1140 => (x"db",x"c1",x"87",x"ec"),
  1141 => (x"c0",x"48",x"bf",x"f4"),
  1142 => (x"c5",x"06",x"a8",x"b7"),
  1143 => (x"db",x"c1",x"87",x"e0"),
  1144 => (x"c3",x"48",x"bf",x"e4"),
  1145 => (x"db",x"01",x"a8",x"b7"),
  1146 => (x"66",x"cc",x"97",x"87"),
  1147 => (x"81",x"c0",x"fe",x"49"),
  1148 => (x"c1",x"1e",x"71",x"b9"),
  1149 => (x"1e",x"bf",x"f0",x"db"),
  1150 => (x"c8",x"87",x"e0",x"fc"),
  1151 => (x"f4",x"db",x"c1",x"86"),
  1152 => (x"87",x"fa",x"c4",x"58"),
  1153 => (x"bf",x"ec",x"db",x"c1"),
  1154 => (x"c1",x"81",x"c3",x"49"),
  1155 => (x"b7",x"bf",x"e4",x"db"),
  1156 => (x"e1",x"c0",x"04",x"a9"),
  1157 => (x"66",x"cc",x"97",x"87"),
  1158 => (x"81",x"c0",x"fe",x"49"),
  1159 => (x"c1",x"1e",x"71",x"b9"),
  1160 => (x"1e",x"bf",x"e8",x"db"),
  1161 => (x"c8",x"87",x"f4",x"fb"),
  1162 => (x"ec",x"db",x"c1",x"86"),
  1163 => (x"f8",x"db",x"c1",x"58"),
  1164 => (x"c4",x"78",x"c1",x"48"),
  1165 => (x"db",x"c1",x"87",x"c8"),
  1166 => (x"c0",x"48",x"bf",x"f4"),
  1167 => (x"c2",x"06",x"a8",x"b7"),
  1168 => (x"db",x"c1",x"87",x"db"),
  1169 => (x"c3",x"48",x"bf",x"f4"),
  1170 => (x"c2",x"01",x"a8",x"b7"),
  1171 => (x"db",x"c1",x"87",x"cf"),
  1172 => (x"c1",x"49",x"bf",x"f0"),
  1173 => (x"db",x"c1",x"81",x"31"),
  1174 => (x"a9",x"b7",x"bf",x"e4"),
  1175 => (x"87",x"df",x"c1",x"04"),
  1176 => (x"49",x"66",x"cc",x"97"),
  1177 => (x"b9",x"81",x"c0",x"fe"),
  1178 => (x"db",x"c1",x"1e",x"71"),
  1179 => (x"fa",x"1e",x"bf",x"fc"),
  1180 => (x"86",x"c8",x"87",x"e9"),
  1181 => (x"58",x"c0",x"dc",x"c1"),
  1182 => (x"bf",x"f8",x"db",x"c1"),
  1183 => (x"c1",x"89",x"c1",x"49"),
  1184 => (x"c0",x"59",x"fc",x"db"),
  1185 => (x"c2",x"03",x"a9",x"b7"),
  1186 => (x"db",x"c1",x"87",x"f4"),
  1187 => (x"c1",x"49",x"bf",x"e8"),
  1188 => (x"bf",x"97",x"fc",x"db"),
  1189 => (x"98",x"ff",x"c3",x"51"),
  1190 => (x"bf",x"e8",x"db",x"c1"),
  1191 => (x"c1",x"81",x"c1",x"49"),
  1192 => (x"c1",x"59",x"ec",x"db"),
  1193 => (x"b7",x"bf",x"c0",x"dc"),
  1194 => (x"c9",x"c0",x"06",x"a9"),
  1195 => (x"c0",x"dc",x"c1",x"87"),
  1196 => (x"e8",x"db",x"c1",x"48"),
  1197 => (x"db",x"c1",x"78",x"bf"),
  1198 => (x"78",x"c1",x"48",x"f8"),
  1199 => (x"c1",x"87",x"ff",x"c1"),
  1200 => (x"05",x"bf",x"f8",x"db"),
  1201 => (x"c1",x"87",x"f7",x"c1"),
  1202 => (x"49",x"bf",x"fc",x"db"),
  1203 => (x"dc",x"c1",x"31",x"c4"),
  1204 => (x"db",x"c1",x"59",x"c0"),
  1205 => (x"97",x"09",x"bf",x"e8"),
  1206 => (x"e1",x"c1",x"09",x"79"),
  1207 => (x"f4",x"db",x"c1",x"87"),
  1208 => (x"b7",x"c7",x"48",x"bf"),
  1209 => (x"d5",x"c1",x"04",x"a8"),
  1210 => (x"fe",x"4b",x"c0",x"87"),
  1211 => (x"78",x"c1",x"48",x"f4"),
  1212 => (x"bf",x"c0",x"dc",x"c1"),
  1213 => (x"c1",x"1e",x"74",x"1e"),
  1214 => (x"fe",x"1e",x"c1",x"cd"),
  1215 => (x"cc",x"87",x"c8",x"f6"),
  1216 => (x"ec",x"db",x"c1",x"86"),
  1217 => (x"e8",x"db",x"c1",x"5c"),
  1218 => (x"dc",x"c1",x"48",x"bf"),
  1219 => (x"a8",x"b7",x"bf",x"c0"),
  1220 => (x"87",x"db",x"c0",x"03"),
  1221 => (x"bf",x"e8",x"db",x"c1"),
  1222 => (x"db",x"c1",x"83",x"bf"),
  1223 => (x"c4",x"49",x"bf",x"e8"),
  1224 => (x"ec",x"db",x"c1",x"81"),
  1225 => (x"c0",x"dc",x"c1",x"59"),
  1226 => (x"04",x"a9",x"b7",x"bf"),
  1227 => (x"73",x"87",x"e5",x"ff"),
  1228 => (x"e0",x"cd",x"c1",x"1e"),
  1229 => (x"ce",x"f5",x"fe",x"1e"),
  1230 => (x"f7",x"86",x"c8",x"87"),
  1231 => (x"d4",x"f7",x"87",x"c6"),
  1232 => (x"65",x"68",x"43",x"87"),
  1233 => (x"75",x"73",x"6b",x"63"),
  1234 => (x"6e",x"69",x"6d",x"6d"),
  1235 => (x"72",x"66",x"20",x"67"),
  1236 => (x"25",x"20",x"6d",x"6f"),
  1237 => (x"6f",x"74",x"20",x"64"),
  1238 => (x"2e",x"64",x"25",x"20"),
  1239 => (x"00",x"20",x"2e",x"2e"),
  1240 => (x"00",x"0a",x"64",x"25"),
  1241 => (x"5c",x"5b",x"5e",x"0e"),
  1242 => (x"d0",x"c1",x"0e",x"5d"),
  1243 => (x"f3",x"fe",x"1e",x"fb"),
  1244 => (x"86",x"c4",x"87",x"e4"),
  1245 => (x"87",x"f1",x"c4",x"ff"),
  1246 => (x"cd",x"02",x"98",x"70"),
  1247 => (x"ed",x"d8",x"ff",x"87"),
  1248 => (x"02",x"98",x"70",x"87"),
  1249 => (x"49",x"c1",x"87",x"c4"),
  1250 => (x"49",x"c0",x"87",x"c2"),
  1251 => (x"d1",x"c1",x"4d",x"71"),
  1252 => (x"f3",x"fe",x"1e",x"d1"),
  1253 => (x"86",x"c4",x"87",x"c0"),
  1254 => (x"48",x"c0",x"dc",x"c1"),
  1255 => (x"ee",x"c0",x"78",x"c0"),
  1256 => (x"d7",x"f2",x"fe",x"1e"),
  1257 => (x"c3",x"86",x"c4",x"87"),
  1258 => (x"4a",x"ff",x"c8",x"f4"),
  1259 => (x"4c",x"bf",x"c0",x"ff"),
  1260 => (x"c0",x"c8",x"49",x"74"),
  1261 => (x"ca",x"c1",x"02",x"99"),
  1262 => (x"c3",x"4b",x"74",x"87"),
  1263 => (x"ab",x"db",x"9b",x"ff"),
  1264 => (x"87",x"f3",x"c0",x"05"),
  1265 => (x"c0",x"02",x"9d",x"75"),
  1266 => (x"c0",x"d0",x"87",x"e3"),
  1267 => (x"1e",x"c0",x"c0",x"c0"),
  1268 => (x"1e",x"df",x"d0",x"c1"),
  1269 => (x"c8",x"87",x"ca",x"f1"),
  1270 => (x"02",x"98",x"70",x"86"),
  1271 => (x"d0",x"c1",x"87",x"cf"),
  1272 => (x"f1",x"fe",x"1e",x"d3"),
  1273 => (x"86",x"c4",x"87",x"f0"),
  1274 => (x"ca",x"87",x"d9",x"f4"),
  1275 => (x"eb",x"d0",x"c1",x"87"),
  1276 => (x"e1",x"f1",x"fe",x"1e"),
  1277 => (x"73",x"86",x"c4",x"87"),
  1278 => (x"87",x"c8",x"f5",x"1e"),
  1279 => (x"f4",x"c3",x"86",x"c4"),
  1280 => (x"72",x"4a",x"c0",x"c9"),
  1281 => (x"71",x"8a",x"c1",x"49"),
  1282 => (x"df",x"fe",x"05",x"99"),
  1283 => (x"87",x"ce",x"fe",x"87"),
  1284 => (x"42",x"87",x"c0",x"f4"),
  1285 => (x"69",x"74",x"6f",x"6f"),
  1286 => (x"2e",x"2e",x"67",x"6e"),
  1287 => (x"42",x"00",x"0a",x"2e"),
  1288 => (x"38",x"54",x"4f",x"4f"),
  1289 => (x"42",x"20",x"32",x"33"),
  1290 => (x"53",x"00",x"4e",x"49"),
  1291 => (x"6f",x"62",x"20",x"44"),
  1292 => (x"66",x"20",x"74",x"6f"),
  1293 => (x"65",x"6c",x"69",x"61"),
  1294 => (x"49",x"00",x"0a",x"64"),
  1295 => (x"69",x"74",x"69",x"6e"),
  1296 => (x"7a",x"69",x"6c",x"61"),
  1297 => (x"20",x"67",x"6e",x"69"),
  1298 => (x"63",x"20",x"44",x"53"),
  1299 => (x"0a",x"64",x"72",x"61"),
  1300 => (x"32",x"53",x"52",x"00"),
  1301 => (x"62",x"20",x"32",x"33"),
  1302 => (x"20",x"74",x"6f",x"6f"),
  1303 => (x"72",x"70",x"20",x"2d"),
  1304 => (x"20",x"73",x"73",x"65"),
  1305 => (x"20",x"43",x"53",x"45"),
  1306 => (x"62",x"20",x"6f",x"74"),
  1307 => (x"20",x"74",x"6f",x"6f"),
  1308 => (x"6d",x"6f",x"72",x"66"),
  1309 => (x"2e",x"44",x"53",x"20"),
  1310 => (x"2e",x"44",x"53",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
