
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"c9",x"01"),
     1 => (x"cf",x"03",x"87",x"cc"),
     2 => (x"87",x"fd",x"00",x"87"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"36",x"27",x"4f",x"00"),
     5 => (x"4f",x"00",x"00",x"00"),
     6 => (x"0e",x"1e",x"18",x"0e"),
     7 => (x"00",x"00",x"44",x"27"),
     8 => (x"48",x"26",x"0f",x"00"),
     9 => (x"08",x"26",x"80",x"ff"),
    10 => (x"c0",x"c0",x"c2",x"4f"),
    11 => (x"05",x"38",x"27",x"4e"),
    12 => (x"00",x"0f",x"00",x"00"),
    13 => (x"f0",x"c1",x"87",x"fd"),
    14 => (x"43",x"27",x"4e",x"c0"),
    15 => (x"0f",x"00",x"00",x"00"),
    16 => (x"4f",x"87",x"fd",x"00"),
    17 => (x"0e",x"1e",x"18",x"0e"),
    18 => (x"80",x"ff",x"48",x"26"),
    19 => (x"1e",x"4f",x"08",x"26"),
    20 => (x"ff",x"1e",x"1e",x"72"),
    21 => (x"48",x"6a",x"4a",x"c0"),
    22 => (x"c4",x"98",x"c0",x"c4"),
    23 => (x"02",x"6e",x"58",x"a6"),
    24 => (x"cc",x"87",x"f3",x"ff"),
    25 => (x"66",x"cc",x"7a",x"66"),
    26 => (x"4a",x"26",x"26",x"48"),
    27 => (x"5e",x"0e",x"4f",x"26"),
    28 => (x"5d",x"5c",x"5b",x"5a"),
    29 => (x"4b",x"66",x"d4",x"0e"),
    30 => (x"4c",x"13",x"4d",x"c0"),
    31 => (x"c0",x"02",x"9c",x"74"),
    32 => (x"4a",x"74",x"87",x"d6"),
    33 => (x"4f",x"27",x"1e",x"72"),
    34 => (x"0f",x"00",x"00",x"00"),
    35 => (x"85",x"c1",x"86",x"c4"),
    36 => (x"9c",x"74",x"4c",x"13"),
    37 => (x"87",x"ea",x"ff",x"05"),
    38 => (x"4d",x"26",x"48",x"75"),
    39 => (x"4b",x"26",x"4c",x"26"),
    40 => (x"4f",x"26",x"4a",x"26"),
    41 => (x"5b",x"5a",x"5e",x"0e"),
    42 => (x"c8",x"0e",x"5d",x"5c"),
    43 => (x"66",x"e0",x"c0",x"8e"),
    44 => (x"4c",x"66",x"dc",x"4d"),
    45 => (x"00",x"16",x"88",x"27"),
    46 => (x"49",x"76",x"4b",x"00"),
    47 => (x"00",x"0e",x"cc",x"27"),
    48 => (x"a6",x"c4",x"79",x"00"),
    49 => (x"c0",x"79",x"c0",x"49"),
    50 => (x"c0",x"03",x"ac",x"b7"),
    51 => (x"ed",x"c0",x"87",x"cd"),
    52 => (x"00",x"4f",x"27",x"1e"),
    53 => (x"c4",x"0f",x"00",x"00"),
    54 => (x"74",x"8c",x"0c",x"86"),
    55 => (x"c6",x"c0",x"05",x"9c"),
    56 => (x"53",x"f0",x"c0",x"87"),
    57 => (x"74",x"87",x"f6",x"c0"),
    58 => (x"f0",x"c0",x"02",x"9c"),
    59 => (x"72",x"49",x"74",x"87"),
    60 => (x"66",x"e8",x"c0",x"1e"),
    61 => (x"04",x"da",x"27",x"4a"),
    62 => (x"26",x"0f",x"00",x"00"),
    63 => (x"72",x"4a",x"71",x"4a"),
    64 => (x"12",x"82",x"6e",x"4a"),
    65 => (x"72",x"49",x"74",x"53"),
    66 => (x"66",x"e8",x"c0",x"1e"),
    67 => (x"04",x"da",x"27",x"4a"),
    68 => (x"26",x"0f",x"00",x"00"),
    69 => (x"74",x"4c",x"70",x"4a"),
    70 => (x"d0",x"ff",x"05",x"9c"),
    71 => (x"16",x"88",x"27",x"87"),
    72 => (x"ab",x"b7",x"00",x"00"),
    73 => (x"87",x"d8",x"c0",x"02"),
    74 => (x"6b",x"97",x"8b",x"c1"),
    75 => (x"48",x"66",x"c4",x"55"),
    76 => (x"a6",x"c8",x"80",x"c1"),
    77 => (x"16",x"88",x"27",x"58"),
    78 => (x"ab",x"b7",x"00",x"00"),
    79 => (x"87",x"e8",x"ff",x"05"),
    80 => (x"66",x"c4",x"55",x"c0"),
    81 => (x"26",x"86",x"c8",x"48"),
    82 => (x"26",x"4c",x"26",x"4d"),
    83 => (x"26",x"4a",x"26",x"4b"),
    84 => (x"5a",x"5e",x"0e",x"4f"),
    85 => (x"0e",x"5d",x"5c",x"5b"),
    86 => (x"76",x"4c",x"c0",x"1e"),
    87 => (x"dc",x"79",x"c0",x"49"),
    88 => (x"66",x"d8",x"4b",x"a6"),
    89 => (x"48",x"66",x"d8",x"4a"),
    90 => (x"a6",x"dc",x"80",x"c1"),
    91 => (x"c1",x"4d",x"12",x"58"),
    92 => (x"c0",x"c0",x"c0",x"c0"),
    93 => (x"b7",x"c0",x"c4",x"95"),
    94 => (x"9d",x"75",x"4d",x"95"),
    95 => (x"87",x"d2",x"c4",x"02"),
    96 => (x"d7",x"c3",x"02",x"6e"),
    97 => (x"c0",x"49",x"76",x"87"),
    98 => (x"c1",x"4a",x"75",x"79"),
    99 => (x"c2",x"02",x"ad",x"e3"),
   100 => (x"e4",x"c1",x"87",x"dd"),
   101 => (x"d8",x"c0",x"02",x"aa"),
   102 => (x"aa",x"ec",x"c1",x"87"),
   103 => (x"87",x"c8",x"c2",x"02"),
   104 => (x"02",x"aa",x"f3",x"c1"),
   105 => (x"c1",x"87",x"e8",x"c1"),
   106 => (x"c0",x"02",x"aa",x"f8"),
   107 => (x"d3",x"c2",x"87",x"f2"),
   108 => (x"27",x"1e",x"ca",x"87"),
   109 => (x"00",x"00",x"16",x"d8"),
   110 => (x"73",x"83",x"c4",x"1e"),
   111 => (x"6a",x"8a",x"c4",x"4a"),
   112 => (x"00",x"a4",x"27",x"1e"),
   113 => (x"cc",x"0f",x"00",x"00"),
   114 => (x"74",x"4a",x"70",x"86"),
   115 => (x"27",x"84",x"72",x"4c"),
   116 => (x"00",x"00",x"16",x"d8"),
   117 => (x"00",x"6e",x"27",x"1e"),
   118 => (x"c4",x"0f",x"00",x"00"),
   119 => (x"87",x"d4",x"c2",x"86"),
   120 => (x"d8",x"27",x"1e",x"d0"),
   121 => (x"1e",x"00",x"00",x"16"),
   122 => (x"4a",x"73",x"83",x"c4"),
   123 => (x"1e",x"6a",x"8a",x"c4"),
   124 => (x"00",x"00",x"a4",x"27"),
   125 => (x"86",x"cc",x"0f",x"00"),
   126 => (x"4c",x"74",x"4a",x"70"),
   127 => (x"d8",x"27",x"84",x"72"),
   128 => (x"1e",x"00",x"00",x"16"),
   129 => (x"00",x"00",x"6e",x"27"),
   130 => (x"86",x"c4",x"0f",x"00"),
   131 => (x"c4",x"87",x"e5",x"c1"),
   132 => (x"c4",x"4a",x"73",x"83"),
   133 => (x"27",x"1e",x"6a",x"8a"),
   134 => (x"00",x"00",x"00",x"6e"),
   135 => (x"70",x"86",x"c4",x"0f"),
   136 => (x"72",x"4c",x"74",x"4a"),
   137 => (x"87",x"cc",x"c1",x"84"),
   138 => (x"79",x"c1",x"49",x"76"),
   139 => (x"c4",x"87",x"c5",x"c1"),
   140 => (x"c4",x"4a",x"73",x"83"),
   141 => (x"27",x"1e",x"6a",x"8a"),
   142 => (x"00",x"00",x"00",x"4f"),
   143 => (x"c1",x"86",x"c4",x"0f"),
   144 => (x"87",x"f0",x"c0",x"84"),
   145 => (x"27",x"1e",x"e5",x"c0"),
   146 => (x"00",x"00",x"00",x"4f"),
   147 => (x"75",x"86",x"c4",x"0f"),
   148 => (x"00",x"4f",x"27",x"1e"),
   149 => (x"c4",x"0f",x"00",x"00"),
   150 => (x"87",x"d8",x"c0",x"86"),
   151 => (x"05",x"ad",x"e5",x"c0"),
   152 => (x"76",x"87",x"c7",x"c0"),
   153 => (x"c0",x"79",x"c1",x"49"),
   154 => (x"1e",x"75",x"87",x"ca"),
   155 => (x"00",x"00",x"4f",x"27"),
   156 => (x"86",x"c4",x"0f",x"00"),
   157 => (x"d8",x"4a",x"66",x"d8"),
   158 => (x"80",x"c1",x"48",x"66"),
   159 => (x"12",x"58",x"a6",x"dc"),
   160 => (x"c0",x"c0",x"c1",x"4d"),
   161 => (x"c4",x"95",x"c0",x"c0"),
   162 => (x"4d",x"95",x"b7",x"c0"),
   163 => (x"fb",x"05",x"9d",x"75"),
   164 => (x"48",x"74",x"87",x"ee"),
   165 => (x"26",x"4d",x"26",x"26"),
   166 => (x"26",x"4b",x"26",x"4c"),
   167 => (x"0e",x"4f",x"26",x"4a"),
   168 => (x"0e",x"5b",x"5a",x"5e"),
   169 => (x"cc",x"4b",x"66",x"d0"),
   170 => (x"66",x"cc",x"7b",x"66"),
   171 => (x"04",x"c6",x"27",x"1e"),
   172 => (x"c4",x"0f",x"00",x"00"),
   173 => (x"72",x"4a",x"70",x"86"),
   174 => (x"c2",x"c0",x"05",x"9a"),
   175 => (x"cc",x"7b",x"c3",x"87"),
   176 => (x"66",x"cc",x"4a",x"66"),
   177 => (x"a9",x"b7",x"c0",x"49"),
   178 => (x"87",x"df",x"c0",x"02"),
   179 => (x"02",x"aa",x"b7",x"c1"),
   180 => (x"c2",x"87",x"dd",x"c0"),
   181 => (x"c0",x"02",x"aa",x"b7"),
   182 => (x"b7",x"c3",x"87",x"ef"),
   183 => (x"ef",x"c0",x"02",x"aa"),
   184 => (x"aa",x"b7",x"c4",x"87"),
   185 => (x"87",x"e6",x"c0",x"02"),
   186 => (x"c0",x"87",x"e5",x"c0"),
   187 => (x"87",x"e0",x"c0",x"7b"),
   188 => (x"00",x"17",x"00",x"27"),
   189 => (x"c1",x"49",x"bf",x"00"),
   190 => (x"06",x"a9",x"b7",x"e4"),
   191 => (x"c0",x"87",x"c5",x"c0"),
   192 => (x"87",x"cc",x"c0",x"7b"),
   193 => (x"c7",x"c0",x"7b",x"c3"),
   194 => (x"c0",x"7b",x"c1",x"87"),
   195 => (x"7b",x"c2",x"87",x"c2"),
   196 => (x"4a",x"26",x"4b",x"26"),
   197 => (x"72",x"1e",x"4f",x"26"),
   198 => (x"4a",x"66",x"c8",x"1e"),
   199 => (x"66",x"cc",x"82",x"c2"),
   200 => (x"d0",x"80",x"72",x"48"),
   201 => (x"79",x"70",x"49",x"66"),
   202 => (x"4f",x"26",x"4a",x"26"),
   203 => (x"5b",x"5a",x"5e",x"0e"),
   204 => (x"dc",x"0e",x"5d",x"5c"),
   205 => (x"85",x"c5",x"4d",x"66"),
   206 => (x"92",x"c4",x"4a",x"75"),
   207 => (x"66",x"d4",x"4a",x"72"),
   208 => (x"66",x"e0",x"c0",x"82"),
   209 => (x"c4",x"4b",x"72",x"7a"),
   210 => (x"c1",x"7b",x"6a",x"83"),
   211 => (x"7a",x"75",x"82",x"f8"),
   212 => (x"4a",x"75",x"4c",x"75"),
   213 => (x"b7",x"72",x"82",x"c1"),
   214 => (x"e1",x"c0",x"01",x"ad"),
   215 => (x"c3",x"4b",x"75",x"87"),
   216 => (x"4b",x"73",x"93",x"c8"),
   217 => (x"74",x"83",x"66",x"d8"),
   218 => (x"72",x"92",x"c4",x"4a"),
   219 => (x"75",x"82",x"73",x"4a"),
   220 => (x"75",x"84",x"c1",x"7a"),
   221 => (x"72",x"82",x"c1",x"4a"),
   222 => (x"ff",x"06",x"ac",x"b7"),
   223 => (x"4c",x"75",x"87",x"df"),
   224 => (x"74",x"94",x"c8",x"c3"),
   225 => (x"84",x"66",x"d8",x"4c"),
   226 => (x"92",x"c4",x"4a",x"75"),
   227 => (x"83",x"72",x"4b",x"74"),
   228 => (x"48",x"6b",x"8b",x"c4"),
   229 => (x"7b",x"70",x"80",x"c1"),
   230 => (x"72",x"4b",x"66",x"d4"),
   231 => (x"e0",x"fe",x"c0",x"83"),
   232 => (x"74",x"4a",x"72",x"84"),
   233 => (x"27",x"7a",x"6b",x"82"),
   234 => (x"00",x"00",x"17",x"00"),
   235 => (x"26",x"79",x"c5",x"49"),
   236 => (x"26",x"4c",x"26",x"4d"),
   237 => (x"26",x"4a",x"26",x"4b"),
   238 => (x"5a",x"5e",x"0e",x"4f"),
   239 => (x"97",x"0e",x"5c",x"5b"),
   240 => (x"74",x"4c",x"66",x"d0"),
   241 => (x"c0",x"c0",x"c1",x"4b"),
   242 => (x"c4",x"93",x"c0",x"c0"),
   243 => (x"4b",x"93",x"b7",x"c0"),
   244 => (x"4a",x"66",x"d4",x"97"),
   245 => (x"c0",x"c0",x"c0",x"c1"),
   246 => (x"c0",x"c4",x"92",x"c0"),
   247 => (x"72",x"4a",x"92",x"b7"),
   248 => (x"c0",x"02",x"ab",x"b7"),
   249 => (x"48",x"c0",x"87",x"c5"),
   250 => (x"27",x"87",x"ca",x"c0"),
   251 => (x"00",x"00",x"17",x"08"),
   252 => (x"c1",x"51",x"74",x"49"),
   253 => (x"26",x"4c",x"26",x"48"),
   254 => (x"26",x"4a",x"26",x"4b"),
   255 => (x"5a",x"5e",x"0e",x"4f"),
   256 => (x"1e",x"0e",x"5c",x"5b"),
   257 => (x"c2",x"4c",x"6e",x"97"),
   258 => (x"4a",x"66",x"d8",x"4b"),
   259 => (x"82",x"73",x"82",x"c1"),
   260 => (x"c1",x"4a",x"6a",x"97"),
   261 => (x"c0",x"c0",x"c0",x"c0"),
   262 => (x"b7",x"c0",x"c4",x"92"),
   263 => (x"1e",x"72",x"4a",x"92"),
   264 => (x"73",x"4a",x"66",x"d8"),
   265 => (x"4a",x"6a",x"97",x"82"),
   266 => (x"c0",x"c0",x"c0",x"c1"),
   267 => (x"c0",x"c4",x"92",x"c0"),
   268 => (x"72",x"4a",x"92",x"b7"),
   269 => (x"03",x"b9",x"27",x"1e"),
   270 => (x"c8",x"0f",x"00",x"00"),
   271 => (x"72",x"4a",x"70",x"86"),
   272 => (x"c5",x"c0",x"05",x"9a"),
   273 => (x"4c",x"c1",x"c1",x"87"),
   274 => (x"b7",x"c2",x"83",x"c1"),
   275 => (x"f8",x"fe",x"06",x"ab"),
   276 => (x"c1",x"4a",x"74",x"87"),
   277 => (x"c0",x"c0",x"c0",x"c0"),
   278 => (x"b7",x"c0",x"c4",x"92"),
   279 => (x"d7",x"c1",x"4a",x"92"),
   280 => (x"c0",x"04",x"aa",x"b7"),
   281 => (x"4a",x"74",x"87",x"d7"),
   282 => (x"c0",x"c0",x"c0",x"c1"),
   283 => (x"c0",x"c4",x"92",x"c0"),
   284 => (x"c1",x"4a",x"92",x"b7"),
   285 => (x"03",x"aa",x"b7",x"da"),
   286 => (x"c7",x"87",x"c2",x"c0"),
   287 => (x"c1",x"4a",x"74",x"4b"),
   288 => (x"c0",x"c0",x"c0",x"c0"),
   289 => (x"b7",x"c0",x"c4",x"92"),
   290 => (x"d2",x"c1",x"4a",x"92"),
   291 => (x"c0",x"05",x"aa",x"b7"),
   292 => (x"48",x"c1",x"87",x"c5"),
   293 => (x"d4",x"87",x"e6",x"c0"),
   294 => (x"66",x"d8",x"4a",x"66"),
   295 => (x"05",x"24",x"27",x"49"),
   296 => (x"70",x"0f",x"00",x"00"),
   297 => (x"aa",x"b7",x"c0",x"4a"),
   298 => (x"87",x"cf",x"c0",x"06"),
   299 => (x"80",x"c7",x"48",x"73"),
   300 => (x"00",x"17",x"04",x"27"),
   301 => (x"48",x"c1",x"58",x"00"),
   302 => (x"c0",x"87",x"c2",x"c0"),
   303 => (x"4c",x"26",x"26",x"48"),
   304 => (x"4a",x"26",x"4b",x"26"),
   305 => (x"c4",x"1e",x"4f",x"26"),
   306 => (x"b7",x"c2",x"49",x"66"),
   307 => (x"c5",x"c0",x"05",x"a9"),
   308 => (x"c0",x"48",x"c1",x"87"),
   309 => (x"48",x"c0",x"87",x"c2"),
   310 => (x"73",x"1e",x"4f",x"26"),
   311 => (x"02",x"9a",x"72",x"1e"),
   312 => (x"48",x"c0",x"87",x"d9"),
   313 => (x"a9",x"72",x"4b",x"c1"),
   314 => (x"83",x"73",x"82",x"01"),
   315 => (x"a9",x"72",x"87",x"f8"),
   316 => (x"80",x"73",x"89",x"03"),
   317 => (x"2b",x"2a",x"c1",x"07"),
   318 => (x"26",x"87",x"f3",x"05"),
   319 => (x"1e",x"4f",x"26",x"4b"),
   320 => (x"4d",x"c0",x"1e",x"75"),
   321 => (x"ff",x"04",x"a1",x"71"),
   322 => (x"bd",x"81",x"c1",x"b9"),
   323 => (x"04",x"a2",x"72",x"07"),
   324 => (x"82",x"c1",x"ba",x"ff"),
   325 => (x"87",x"c2",x"07",x"bd"),
   326 => (x"ff",x"05",x"9d",x"75"),
   327 => (x"07",x"80",x"c1",x"b8"),
   328 => (x"4f",x"26",x"4d",x"25"),
   329 => (x"11",x"48",x"12",x"1e"),
   330 => (x"88",x"87",x"c4",x"02"),
   331 => (x"26",x"87",x"f6",x"02"),
   332 => (x"c8",x"ff",x"1e",x"4f"),
   333 => (x"4f",x"26",x"48",x"bf"),
   334 => (x"5b",x"5a",x"5e",x"0e"),
   335 => (x"d0",x"0e",x"5d",x"5c"),
   336 => (x"4c",x"66",x"c4",x"8e"),
   337 => (x"00",x"16",x"fc",x"27"),
   338 => (x"00",x"27",x"49",x"00"),
   339 => (x"79",x"00",x"00",x"3f"),
   340 => (x"00",x"16",x"f8",x"27"),
   341 => (x"30",x"27",x"49",x"00"),
   342 => (x"79",x"00",x"00",x"3f"),
   343 => (x"00",x"3f",x"30",x"27"),
   344 => (x"00",x"27",x"49",x"00"),
   345 => (x"79",x"00",x"00",x"3f"),
   346 => (x"00",x"3f",x"34",x"27"),
   347 => (x"79",x"c0",x"49",x"00"),
   348 => (x"00",x"3f",x"38",x"27"),
   349 => (x"79",x"c2",x"49",x"00"),
   350 => (x"00",x"3f",x"3c",x"27"),
   351 => (x"e8",x"c0",x"49",x"00"),
   352 => (x"3f",x"40",x"27",x"79"),
   353 => (x"27",x"49",x"00",x"00"),
   354 => (x"00",x"00",x"10",x"56"),
   355 => (x"20",x"1e",x"72",x"48"),
   356 => (x"20",x"81",x"c4",x"79"),
   357 => (x"20",x"81",x"c4",x"79"),
   358 => (x"20",x"81",x"c4",x"79"),
   359 => (x"20",x"81",x"c4",x"79"),
   360 => (x"20",x"81",x"c4",x"79"),
   361 => (x"20",x"81",x"c4",x"79"),
   362 => (x"10",x"81",x"c4",x"79"),
   363 => (x"10",x"51",x"10",x"51"),
   364 => (x"27",x"4a",x"26",x"51"),
   365 => (x"00",x"00",x"3f",x"60"),
   366 => (x"10",x"75",x"27",x"49"),
   367 => (x"72",x"48",x"00",x"00"),
   368 => (x"c4",x"79",x"20",x"1e"),
   369 => (x"c4",x"79",x"20",x"81"),
   370 => (x"c4",x"79",x"20",x"81"),
   371 => (x"c4",x"79",x"20",x"81"),
   372 => (x"c4",x"79",x"20",x"81"),
   373 => (x"c4",x"79",x"20",x"81"),
   374 => (x"c4",x"79",x"20",x"81"),
   375 => (x"10",x"51",x"10",x"81"),
   376 => (x"26",x"51",x"10",x"51"),
   377 => (x"1e",x"34",x"27",x"4a"),
   378 => (x"ca",x"49",x"00",x"00"),
   379 => (x"10",x"94",x"27",x"79"),
   380 => (x"27",x"1e",x"00",x"00"),
   381 => (x"00",x"00",x"01",x"51"),
   382 => (x"27",x"86",x"c4",x"0f"),
   383 => (x"00",x"00",x"10",x"96"),
   384 => (x"01",x"51",x"27",x"1e"),
   385 => (x"c4",x"0f",x"00",x"00"),
   386 => (x"10",x"c6",x"27",x"86"),
   387 => (x"27",x"1e",x"00",x"00"),
   388 => (x"00",x"00",x"01",x"51"),
   389 => (x"27",x"86",x"c4",x"0f"),
   390 => (x"00",x"00",x"16",x"7c"),
   391 => (x"df",x"c0",x"02",x"bf"),
   392 => (x"0e",x"dd",x"27",x"87"),
   393 => (x"27",x"1e",x"00",x"00"),
   394 => (x"00",x"00",x"01",x"51"),
   395 => (x"27",x"86",x"c4",x"0f"),
   396 => (x"00",x"00",x"0f",x"09"),
   397 => (x"01",x"51",x"27",x"1e"),
   398 => (x"c4",x"0f",x"00",x"00"),
   399 => (x"87",x"dc",x"c0",x"86"),
   400 => (x"00",x"0f",x"0b",x"27"),
   401 => (x"51",x"27",x"1e",x"00"),
   402 => (x"0f",x"00",x"00",x"01"),
   403 => (x"3a",x"27",x"86",x"c4"),
   404 => (x"1e",x"00",x"00",x"0f"),
   405 => (x"00",x"01",x"51",x"27"),
   406 => (x"86",x"c4",x"0f",x"00"),
   407 => (x"00",x"16",x"80",x"27"),
   408 => (x"27",x"1e",x"bf",x"00"),
   409 => (x"00",x"00",x"10",x"c8"),
   410 => (x"01",x"51",x"27",x"1e"),
   411 => (x"c8",x"0f",x"00",x"00"),
   412 => (x"05",x"31",x"27",x"86"),
   413 => (x"27",x"0f",x"00",x"00"),
   414 => (x"00",x"00",x"3e",x"ec"),
   415 => (x"27",x"4d",x"c1",x"58"),
   416 => (x"00",x"00",x"16",x"80"),
   417 => (x"b7",x"c0",x"49",x"bf"),
   418 => (x"d5",x"c7",x"06",x"a9"),
   419 => (x"0e",x"b8",x"27",x"87"),
   420 => (x"27",x"0f",x"00",x"00"),
   421 => (x"00",x"00",x"0e",x"77"),
   422 => (x"c2",x"49",x"76",x"0f"),
   423 => (x"27",x"4c",x"c3",x"79"),
   424 => (x"00",x"00",x"3f",x"80"),
   425 => (x"0f",x"5b",x"27",x"49"),
   426 => (x"72",x"48",x"00",x"00"),
   427 => (x"c4",x"79",x"20",x"1e"),
   428 => (x"c4",x"79",x"20",x"81"),
   429 => (x"c4",x"79",x"20",x"81"),
   430 => (x"c4",x"79",x"20",x"81"),
   431 => (x"c4",x"79",x"20",x"81"),
   432 => (x"c4",x"79",x"20",x"81"),
   433 => (x"c4",x"79",x"20",x"81"),
   434 => (x"10",x"51",x"10",x"81"),
   435 => (x"26",x"51",x"10",x"51"),
   436 => (x"49",x"a6",x"c8",x"4a"),
   437 => (x"80",x"27",x"79",x"c1"),
   438 => (x"1e",x"00",x"00",x"3f"),
   439 => (x"00",x"3f",x"60",x"27"),
   440 => (x"fd",x"27",x"1e",x"00"),
   441 => (x"0f",x"00",x"00",x"03"),
   442 => (x"4a",x"70",x"86",x"c8"),
   443 => (x"c0",x"05",x"9a",x"72"),
   444 => (x"4a",x"c1",x"87",x"c5"),
   445 => (x"c0",x"87",x"c2",x"c0"),
   446 => (x"17",x"04",x"27",x"4a"),
   447 => (x"72",x"49",x"00",x"00"),
   448 => (x"74",x"49",x"6e",x"79"),
   449 => (x"c0",x"03",x"a9",x"b7"),
   450 => (x"4a",x"6e",x"87",x"ed"),
   451 => (x"48",x"72",x"92",x"c5"),
   452 => (x"a6",x"d0",x"88",x"74"),
   453 => (x"4a",x"a6",x"cc",x"58"),
   454 => (x"1e",x"74",x"1e",x"72"),
   455 => (x"27",x"1e",x"66",x"c8"),
   456 => (x"00",x"00",x"03",x"16"),
   457 => (x"6e",x"86",x"cc",x"0f"),
   458 => (x"c4",x"80",x"c1",x"48"),
   459 => (x"49",x"6e",x"58",x"a6"),
   460 => (x"04",x"a9",x"b7",x"74"),
   461 => (x"cc",x"87",x"d3",x"ff"),
   462 => (x"66",x"c4",x"1e",x"66"),
   463 => (x"17",x"d8",x"27",x"1e"),
   464 => (x"27",x"1e",x"00",x"00"),
   465 => (x"00",x"00",x"17",x"10"),
   466 => (x"03",x"2c",x"27",x"1e"),
   467 => (x"d0",x"0f",x"00",x"00"),
   468 => (x"16",x"f8",x"27",x"86"),
   469 => (x"1e",x"bf",x"00",x"00"),
   470 => (x"00",x"0d",x"54",x"27"),
   471 => (x"86",x"c4",x"0f",x"00"),
   472 => (x"c1",x"49",x"a6",x"c4"),
   473 => (x"09",x"27",x"51",x"c1"),
   474 => (x"97",x"00",x"00",x"17"),
   475 => (x"c0",x"c1",x"4a",x"bf"),
   476 => (x"92",x"c0",x"c0",x"c0"),
   477 => (x"92",x"b7",x"c0",x"c4"),
   478 => (x"b7",x"c1",x"c1",x"4a"),
   479 => (x"e6",x"c2",x"04",x"aa"),
   480 => (x"1e",x"c3",x"c1",x"87"),
   481 => (x"4a",x"66",x"c8",x"97"),
   482 => (x"c0",x"c0",x"c0",x"c1"),
   483 => (x"c0",x"c4",x"92",x"c0"),
   484 => (x"72",x"4a",x"92",x"b7"),
   485 => (x"03",x"b9",x"27",x"1e"),
   486 => (x"c8",x"0f",x"00",x"00"),
   487 => (x"c8",x"4a",x"70",x"86"),
   488 => (x"b7",x"72",x"49",x"66"),
   489 => (x"cb",x"c1",x"05",x"a9"),
   490 => (x"4a",x"a6",x"c8",x"87"),
   491 => (x"1e",x"c0",x"1e",x"72"),
   492 => (x"00",x"02",x"9f",x"27"),
   493 => (x"86",x"c8",x"0f",x"00"),
   494 => (x"00",x"3f",x"80",x"27"),
   495 => (x"3c",x"27",x"49",x"00"),
   496 => (x"48",x"00",x"00",x"0f"),
   497 => (x"79",x"20",x"1e",x"72"),
   498 => (x"79",x"20",x"81",x"c4"),
   499 => (x"79",x"20",x"81",x"c4"),
   500 => (x"79",x"20",x"81",x"c4"),
   501 => (x"79",x"20",x"81",x"c4"),
   502 => (x"79",x"20",x"81",x"c4"),
   503 => (x"79",x"20",x"81",x"c4"),
   504 => (x"51",x"10",x"81",x"c4"),
   505 => (x"51",x"10",x"51",x"10"),
   506 => (x"4c",x"75",x"4a",x"26"),
   507 => (x"00",x"17",x"00",x"27"),
   508 => (x"79",x"75",x"49",x"00"),
   509 => (x"48",x"66",x"c4",x"97"),
   510 => (x"a6",x"c4",x"80",x"c1"),
   511 => (x"c4",x"97",x"50",x"08"),
   512 => (x"c0",x"c1",x"4b",x"66"),
   513 => (x"93",x"c0",x"c0",x"c0"),
   514 => (x"93",x"b7",x"c0",x"c4"),
   515 => (x"17",x"09",x"27",x"4b"),
   516 => (x"bf",x"97",x"00",x"00"),
   517 => (x"c0",x"c0",x"c1",x"4a"),
   518 => (x"c4",x"92",x"c0",x"c0"),
   519 => (x"4a",x"92",x"b7",x"c0"),
   520 => (x"06",x"ab",x"b7",x"72"),
   521 => (x"6e",x"87",x"da",x"fd"),
   522 => (x"72",x"49",x"74",x"94"),
   523 => (x"4a",x"66",x"d0",x"1e"),
   524 => (x"00",x"04",x"da",x"27"),
   525 => (x"4a",x"26",x"0f",x"00"),
   526 => (x"a6",x"c4",x"48",x"70"),
   527 => (x"cc",x"4a",x"74",x"58"),
   528 => (x"92",x"c7",x"8a",x"66"),
   529 => (x"8c",x"6e",x"4c",x"72"),
   530 => (x"1e",x"72",x"4a",x"76"),
   531 => (x"00",x"0d",x"f3",x"27"),
   532 => (x"86",x"c4",x"0f",x"00"),
   533 => (x"80",x"27",x"85",x"c1"),
   534 => (x"bf",x"00",x"00",x"16"),
   535 => (x"f8",x"06",x"ad",x"b7"),
   536 => (x"31",x"27",x"87",x"eb"),
   537 => (x"0f",x"00",x"00",x"05"),
   538 => (x"00",x"3e",x"f0",x"27"),
   539 => (x"f5",x"27",x"58",x"00"),
   540 => (x"1e",x"00",x"00",x"10"),
   541 => (x"00",x"01",x"51",x"27"),
   542 => (x"86",x"c4",x"0f",x"00"),
   543 => (x"00",x"11",x"05",x"27"),
   544 => (x"51",x"27",x"1e",x"00"),
   545 => (x"0f",x"00",x"00",x"01"),
   546 => (x"07",x"27",x"86",x"c4"),
   547 => (x"1e",x"00",x"00",x"11"),
   548 => (x"00",x"01",x"51",x"27"),
   549 => (x"86",x"c4",x"0f",x"00"),
   550 => (x"00",x"11",x"3d",x"27"),
   551 => (x"51",x"27",x"1e",x"00"),
   552 => (x"0f",x"00",x"00",x"01"),
   553 => (x"00",x"27",x"86",x"c4"),
   554 => (x"bf",x"00",x"00",x"17"),
   555 => (x"11",x"3f",x"27",x"1e"),
   556 => (x"27",x"1e",x"00",x"00"),
   557 => (x"00",x"00",x"01",x"51"),
   558 => (x"c5",x"86",x"c8",x"0f"),
   559 => (x"11",x"58",x"27",x"1e"),
   560 => (x"27",x"1e",x"00",x"00"),
   561 => (x"00",x"00",x"01",x"51"),
   562 => (x"27",x"86",x"c8",x"0f"),
   563 => (x"00",x"00",x"17",x"04"),
   564 => (x"71",x"27",x"1e",x"bf"),
   565 => (x"1e",x"00",x"00",x"11"),
   566 => (x"00",x"01",x"51",x"27"),
   567 => (x"86",x"c8",x"0f",x"00"),
   568 => (x"8a",x"27",x"1e",x"c1"),
   569 => (x"1e",x"00",x"00",x"11"),
   570 => (x"00",x"01",x"51",x"27"),
   571 => (x"86",x"c8",x"0f",x"00"),
   572 => (x"00",x"17",x"08",x"27"),
   573 => (x"4a",x"bf",x"97",x"00"),
   574 => (x"c0",x"c0",x"c0",x"c1"),
   575 => (x"c0",x"c4",x"92",x"c0"),
   576 => (x"72",x"4a",x"92",x"b7"),
   577 => (x"11",x"a3",x"27",x"1e"),
   578 => (x"27",x"1e",x"00",x"00"),
   579 => (x"00",x"00",x"01",x"51"),
   580 => (x"c1",x"86",x"c8",x"0f"),
   581 => (x"bc",x"27",x"1e",x"c1"),
   582 => (x"1e",x"00",x"00",x"11"),
   583 => (x"00",x"01",x"51",x"27"),
   584 => (x"86",x"c8",x"0f",x"00"),
   585 => (x"00",x"17",x"09",x"27"),
   586 => (x"4a",x"bf",x"97",x"00"),
   587 => (x"c0",x"c0",x"c0",x"c1"),
   588 => (x"c0",x"c4",x"92",x"c0"),
   589 => (x"72",x"4a",x"92",x"b7"),
   590 => (x"11",x"d5",x"27",x"1e"),
   591 => (x"27",x"1e",x"00",x"00"),
   592 => (x"00",x"00",x"01",x"51"),
   593 => (x"c1",x"86",x"c8",x"0f"),
   594 => (x"ee",x"27",x"1e",x"c2"),
   595 => (x"1e",x"00",x"00",x"11"),
   596 => (x"00",x"01",x"51",x"27"),
   597 => (x"86",x"c8",x"0f",x"00"),
   598 => (x"00",x"17",x"30",x"27"),
   599 => (x"27",x"1e",x"bf",x"00"),
   600 => (x"00",x"00",x"12",x"07"),
   601 => (x"01",x"51",x"27",x"1e"),
   602 => (x"c8",x"0f",x"00",x"00"),
   603 => (x"27",x"1e",x"c7",x"86"),
   604 => (x"00",x"00",x"12",x"20"),
   605 => (x"01",x"51",x"27",x"1e"),
   606 => (x"c8",x"0f",x"00",x"00"),
   607 => (x"1e",x"34",x"27",x"86"),
   608 => (x"1e",x"bf",x"00",x"00"),
   609 => (x"00",x"12",x"39",x"27"),
   610 => (x"51",x"27",x"1e",x"00"),
   611 => (x"0f",x"00",x"00",x"01"),
   612 => (x"52",x"27",x"86",x"c8"),
   613 => (x"1e",x"00",x"00",x"12"),
   614 => (x"00",x"01",x"51",x"27"),
   615 => (x"86",x"c4",x"0f",x"00"),
   616 => (x"00",x"12",x"7c",x"27"),
   617 => (x"51",x"27",x"1e",x"00"),
   618 => (x"0f",x"00",x"00",x"01"),
   619 => (x"f8",x"27",x"86",x"c4"),
   620 => (x"bf",x"00",x"00",x"16"),
   621 => (x"88",x"27",x"1e",x"bf"),
   622 => (x"1e",x"00",x"00",x"12"),
   623 => (x"00",x"01",x"51",x"27"),
   624 => (x"86",x"c8",x"0f",x"00"),
   625 => (x"00",x"12",x"a1",x"27"),
   626 => (x"51",x"27",x"1e",x"00"),
   627 => (x"0f",x"00",x"00",x"01"),
   628 => (x"f8",x"27",x"86",x"c4"),
   629 => (x"bf",x"00",x"00",x"16"),
   630 => (x"6a",x"82",x"c4",x"4a"),
   631 => (x"12",x"d2",x"27",x"1e"),
   632 => (x"27",x"1e",x"00",x"00"),
   633 => (x"00",x"00",x"01",x"51"),
   634 => (x"c0",x"86",x"c8",x"0f"),
   635 => (x"12",x"eb",x"27",x"1e"),
   636 => (x"27",x"1e",x"00",x"00"),
   637 => (x"00",x"00",x"01",x"51"),
   638 => (x"27",x"86",x"c8",x"0f"),
   639 => (x"00",x"00",x"16",x"f8"),
   640 => (x"82",x"c8",x"4a",x"bf"),
   641 => (x"04",x"27",x"1e",x"6a"),
   642 => (x"1e",x"00",x"00",x"13"),
   643 => (x"00",x"01",x"51",x"27"),
   644 => (x"86",x"c8",x"0f",x"00"),
   645 => (x"1d",x"27",x"1e",x"c2"),
   646 => (x"1e",x"00",x"00",x"13"),
   647 => (x"00",x"01",x"51",x"27"),
   648 => (x"86",x"c8",x"0f",x"00"),
   649 => (x"00",x"16",x"f8",x"27"),
   650 => (x"cc",x"4a",x"bf",x"00"),
   651 => (x"27",x"1e",x"6a",x"82"),
   652 => (x"00",x"00",x"13",x"36"),
   653 => (x"01",x"51",x"27",x"1e"),
   654 => (x"c8",x"0f",x"00",x"00"),
   655 => (x"27",x"1e",x"d1",x"86"),
   656 => (x"00",x"00",x"13",x"4f"),
   657 => (x"01",x"51",x"27",x"1e"),
   658 => (x"c8",x"0f",x"00",x"00"),
   659 => (x"16",x"f8",x"27",x"86"),
   660 => (x"4a",x"bf",x"00",x"00"),
   661 => (x"1e",x"72",x"82",x"d0"),
   662 => (x"00",x"13",x"68",x"27"),
   663 => (x"51",x"27",x"1e",x"00"),
   664 => (x"0f",x"00",x"00",x"01"),
   665 => (x"81",x"27",x"86",x"c8"),
   666 => (x"1e",x"00",x"00",x"13"),
   667 => (x"00",x"01",x"51",x"27"),
   668 => (x"86",x"c4",x"0f",x"00"),
   669 => (x"00",x"13",x"b6",x"27"),
   670 => (x"51",x"27",x"1e",x"00"),
   671 => (x"0f",x"00",x"00",x"01"),
   672 => (x"fc",x"27",x"86",x"c4"),
   673 => (x"bf",x"00",x"00",x"16"),
   674 => (x"c7",x"27",x"1e",x"bf"),
   675 => (x"1e",x"00",x"00",x"13"),
   676 => (x"00",x"01",x"51",x"27"),
   677 => (x"86",x"c8",x"0f",x"00"),
   678 => (x"00",x"13",x"e0",x"27"),
   679 => (x"51",x"27",x"1e",x"00"),
   680 => (x"0f",x"00",x"00",x"01"),
   681 => (x"fc",x"27",x"86",x"c4"),
   682 => (x"bf",x"00",x"00",x"16"),
   683 => (x"6a",x"82",x"c4",x"4a"),
   684 => (x"14",x"20",x"27",x"1e"),
   685 => (x"27",x"1e",x"00",x"00"),
   686 => (x"00",x"00",x"01",x"51"),
   687 => (x"c0",x"86",x"c8",x"0f"),
   688 => (x"14",x"39",x"27",x"1e"),
   689 => (x"27",x"1e",x"00",x"00"),
   690 => (x"00",x"00",x"01",x"51"),
   691 => (x"27",x"86",x"c8",x"0f"),
   692 => (x"00",x"00",x"16",x"fc"),
   693 => (x"82",x"c8",x"4a",x"bf"),
   694 => (x"52",x"27",x"1e",x"6a"),
   695 => (x"1e",x"00",x"00",x"14"),
   696 => (x"00",x"01",x"51",x"27"),
   697 => (x"86",x"c8",x"0f",x"00"),
   698 => (x"6b",x"27",x"1e",x"c1"),
   699 => (x"1e",x"00",x"00",x"14"),
   700 => (x"00",x"01",x"51",x"27"),
   701 => (x"86",x"c8",x"0f",x"00"),
   702 => (x"00",x"16",x"fc",x"27"),
   703 => (x"cc",x"4a",x"bf",x"00"),
   704 => (x"27",x"1e",x"6a",x"82"),
   705 => (x"00",x"00",x"14",x"84"),
   706 => (x"01",x"51",x"27",x"1e"),
   707 => (x"c8",x"0f",x"00",x"00"),
   708 => (x"27",x"1e",x"d2",x"86"),
   709 => (x"00",x"00",x"14",x"9d"),
   710 => (x"01",x"51",x"27",x"1e"),
   711 => (x"c8",x"0f",x"00",x"00"),
   712 => (x"16",x"fc",x"27",x"86"),
   713 => (x"4a",x"bf",x"00",x"00"),
   714 => (x"1e",x"72",x"82",x"d0"),
   715 => (x"00",x"14",x"b6",x"27"),
   716 => (x"51",x"27",x"1e",x"00"),
   717 => (x"0f",x"00",x"00",x"01"),
   718 => (x"cf",x"27",x"86",x"c8"),
   719 => (x"1e",x"00",x"00",x"14"),
   720 => (x"00",x"01",x"51",x"27"),
   721 => (x"86",x"c4",x"0f",x"00"),
   722 => (x"04",x"27",x"1e",x"6e"),
   723 => (x"1e",x"00",x"00",x"15"),
   724 => (x"00",x"01",x"51",x"27"),
   725 => (x"86",x"c8",x"0f",x"00"),
   726 => (x"1d",x"27",x"1e",x"c5"),
   727 => (x"1e",x"00",x"00",x"15"),
   728 => (x"00",x"01",x"51",x"27"),
   729 => (x"86",x"c8",x"0f",x"00"),
   730 => (x"36",x"27",x"1e",x"74"),
   731 => (x"1e",x"00",x"00",x"15"),
   732 => (x"00",x"01",x"51",x"27"),
   733 => (x"86",x"c8",x"0f",x"00"),
   734 => (x"4f",x"27",x"1e",x"cd"),
   735 => (x"1e",x"00",x"00",x"15"),
   736 => (x"00",x"01",x"51",x"27"),
   737 => (x"86",x"c8",x"0f",x"00"),
   738 => (x"27",x"1e",x"66",x"cc"),
   739 => (x"00",x"00",x"15",x"68"),
   740 => (x"01",x"51",x"27",x"1e"),
   741 => (x"c8",x"0f",x"00",x"00"),
   742 => (x"27",x"1e",x"c7",x"86"),
   743 => (x"00",x"00",x"15",x"81"),
   744 => (x"01",x"51",x"27",x"1e"),
   745 => (x"c8",x"0f",x"00",x"00"),
   746 => (x"1e",x"66",x"c8",x"86"),
   747 => (x"00",x"15",x"9a",x"27"),
   748 => (x"51",x"27",x"1e",x"00"),
   749 => (x"0f",x"00",x"00",x"01"),
   750 => (x"1e",x"c1",x"86",x"c8"),
   751 => (x"00",x"15",x"b3",x"27"),
   752 => (x"51",x"27",x"1e",x"00"),
   753 => (x"0f",x"00",x"00",x"01"),
   754 => (x"60",x"27",x"86",x"c8"),
   755 => (x"1e",x"00",x"00",x"3f"),
   756 => (x"00",x"15",x"cc",x"27"),
   757 => (x"51",x"27",x"1e",x"00"),
   758 => (x"0f",x"00",x"00",x"01"),
   759 => (x"e5",x"27",x"86",x"c8"),
   760 => (x"1e",x"00",x"00",x"15"),
   761 => (x"00",x"01",x"51",x"27"),
   762 => (x"86",x"c4",x"0f",x"00"),
   763 => (x"00",x"3f",x"80",x"27"),
   764 => (x"1a",x"27",x"1e",x"00"),
   765 => (x"1e",x"00",x"00",x"16"),
   766 => (x"00",x"01",x"51",x"27"),
   767 => (x"86",x"c8",x"0f",x"00"),
   768 => (x"00",x"16",x"33",x"27"),
   769 => (x"51",x"27",x"1e",x"00"),
   770 => (x"0f",x"00",x"00",x"01"),
   771 => (x"68",x"27",x"86",x"c4"),
   772 => (x"1e",x"00",x"00",x"16"),
   773 => (x"00",x"01",x"51",x"27"),
   774 => (x"86",x"c4",x"0f",x"00"),
   775 => (x"00",x"3e",x"ec",x"27"),
   776 => (x"27",x"4a",x"bf",x"00"),
   777 => (x"00",x"00",x"3e",x"e8"),
   778 => (x"f0",x"27",x"8a",x"bf"),
   779 => (x"49",x"00",x"00",x"3e"),
   780 => (x"1e",x"72",x"79",x"72"),
   781 => (x"00",x"16",x"6a",x"27"),
   782 => (x"51",x"27",x"1e",x"00"),
   783 => (x"0f",x"00",x"00",x"01"),
   784 => (x"f0",x"27",x"86",x"c8"),
   785 => (x"bf",x"00",x"00",x"3e"),
   786 => (x"b7",x"f8",x"c1",x"49"),
   787 => (x"ea",x"c0",x"03",x"a9"),
   788 => (x"0f",x"7a",x"27",x"87"),
   789 => (x"27",x"1e",x"00",x"00"),
   790 => (x"00",x"00",x"01",x"51"),
   791 => (x"27",x"86",x"c4",x"0f"),
   792 => (x"00",x"00",x"0f",x"b0"),
   793 => (x"01",x"51",x"27",x"1e"),
   794 => (x"c4",x"0f",x"00",x"00"),
   795 => (x"0f",x"d0",x"27",x"86"),
   796 => (x"27",x"1e",x"00",x"00"),
   797 => (x"00",x"00",x"01",x"51"),
   798 => (x"27",x"86",x"c4",x"0f"),
   799 => (x"00",x"00",x"3e",x"f0"),
   800 => (x"4b",x"72",x"4a",x"bf"),
   801 => (x"73",x"93",x"e8",x"cf"),
   802 => (x"27",x"1e",x"72",x"49"),
   803 => (x"00",x"00",x"16",x"80"),
   804 => (x"da",x"27",x"4a",x"bf"),
   805 => (x"0f",x"00",x"00",x"04"),
   806 => (x"48",x"70",x"4a",x"26"),
   807 => (x"00",x"3e",x"f8",x"27"),
   808 => (x"80",x"27",x"58",x"00"),
   809 => (x"bf",x"00",x"00",x"16"),
   810 => (x"cf",x"4c",x"73",x"4b"),
   811 => (x"49",x"74",x"94",x"e8"),
   812 => (x"4a",x"72",x"1e",x"72"),
   813 => (x"00",x"04",x"da",x"27"),
   814 => (x"4a",x"26",x"0f",x"00"),
   815 => (x"fc",x"27",x"48",x"70"),
   816 => (x"58",x"00",x"00",x"3e"),
   817 => (x"73",x"93",x"f9",x"c8"),
   818 => (x"72",x"1e",x"72",x"49"),
   819 => (x"04",x"da",x"27",x"4a"),
   820 => (x"26",x"0f",x"00",x"00"),
   821 => (x"27",x"48",x"70",x"4a"),
   822 => (x"00",x"00",x"3f",x"00"),
   823 => (x"0f",x"d2",x"27",x"58"),
   824 => (x"27",x"1e",x"00",x"00"),
   825 => (x"00",x"00",x"01",x"51"),
   826 => (x"27",x"86",x"c4",x"0f"),
   827 => (x"00",x"00",x"3e",x"f4"),
   828 => (x"ff",x"27",x"1e",x"bf"),
   829 => (x"1e",x"00",x"00",x"0f"),
   830 => (x"00",x"01",x"51",x"27"),
   831 => (x"86",x"c8",x"0f",x"00"),
   832 => (x"00",x"10",x"04",x"27"),
   833 => (x"51",x"27",x"1e",x"00"),
   834 => (x"0f",x"00",x"00",x"01"),
   835 => (x"f8",x"27",x"86",x"c4"),
   836 => (x"bf",x"00",x"00",x"3e"),
   837 => (x"10",x"31",x"27",x"1e"),
   838 => (x"27",x"1e",x"00",x"00"),
   839 => (x"00",x"00",x"01",x"51"),
   840 => (x"27",x"86",x"c8",x"0f"),
   841 => (x"00",x"00",x"3e",x"fc"),
   842 => (x"36",x"27",x"1e",x"bf"),
   843 => (x"1e",x"00",x"00",x"10"),
   844 => (x"00",x"01",x"51",x"27"),
   845 => (x"86",x"c8",x"0f",x"00"),
   846 => (x"00",x"10",x"54",x"27"),
   847 => (x"51",x"27",x"1e",x"00"),
   848 => (x"0f",x"00",x"00",x"01"),
   849 => (x"48",x"c0",x"86",x"c4"),
   850 => (x"4d",x"26",x"86",x"d0"),
   851 => (x"4b",x"26",x"4c",x"26"),
   852 => (x"4f",x"26",x"4a",x"26"),
   853 => (x"5b",x"5a",x"5e",x"0e"),
   854 => (x"d4",x"0e",x"5d",x"5c"),
   855 => (x"72",x"4a",x"bf",x"66"),
   856 => (x"16",x"f8",x"27",x"4d"),
   857 => (x"48",x"bf",x"00",x"00"),
   858 => (x"f0",x"c0",x"1e",x"72"),
   859 => (x"7a",x"20",x"49",x"a2"),
   860 => (x"a9",x"72",x"82",x"c4"),
   861 => (x"26",x"87",x"f7",x"05"),
   862 => (x"4c",x"66",x"d4",x"4a"),
   863 => (x"7c",x"c5",x"84",x"cc"),
   864 => (x"83",x"cc",x"4b",x"72"),
   865 => (x"66",x"d4",x"7b",x"6c"),
   866 => (x"1e",x"72",x"7a",x"bf"),
   867 => (x"00",x"0e",x"3f",x"27"),
   868 => (x"86",x"c4",x"0f",x"00"),
   869 => (x"9a",x"6a",x"82",x"c4"),
   870 => (x"87",x"f4",x"c0",x"05"),
   871 => (x"83",x"c8",x"4b",x"75"),
   872 => (x"82",x"cc",x"4a",x"75"),
   873 => (x"1e",x"73",x"7a",x"c6"),
   874 => (x"c8",x"4b",x"66",x"d8"),
   875 => (x"27",x"1e",x"6b",x"83"),
   876 => (x"00",x"00",x"02",x"9f"),
   877 => (x"27",x"86",x"c8",x"0f"),
   878 => (x"00",x"00",x"16",x"f8"),
   879 => (x"72",x"7d",x"bf",x"bf"),
   880 => (x"6a",x"1e",x"ca",x"1e"),
   881 => (x"03",x"16",x"27",x"1e"),
   882 => (x"cc",x"0f",x"00",x"00"),
   883 => (x"87",x"d9",x"c0",x"86"),
   884 => (x"4a",x"bf",x"66",x"d4"),
   885 => (x"48",x"49",x"66",x"d4"),
   886 => (x"f0",x"c0",x"1e",x"72"),
   887 => (x"79",x"20",x"4a",x"a1"),
   888 => (x"aa",x"71",x"81",x"c4"),
   889 => (x"26",x"87",x"f7",x"05"),
   890 => (x"26",x"4d",x"26",x"4a"),
   891 => (x"26",x"4b",x"26",x"4c"),
   892 => (x"0e",x"4f",x"26",x"4a"),
   893 => (x"5c",x"5b",x"5a",x"5e"),
   894 => (x"6e",x"1e",x"0e",x"5d"),
   895 => (x"4c",x"66",x"d8",x"4d"),
   896 => (x"83",x"ca",x"4b",x"6c"),
   897 => (x"00",x"17",x"08",x"27"),
   898 => (x"4a",x"bf",x"97",x"00"),
   899 => (x"c0",x"c0",x"c0",x"c1"),
   900 => (x"c0",x"c4",x"92",x"c0"),
   901 => (x"c1",x"4a",x"92",x"b7"),
   902 => (x"05",x"aa",x"b7",x"c1"),
   903 => (x"c1",x"87",x"cf",x"c0"),
   904 => (x"27",x"48",x"73",x"8b"),
   905 => (x"00",x"00",x"17",x"00"),
   906 => (x"7c",x"70",x"88",x"bf"),
   907 => (x"9d",x"75",x"4d",x"c0"),
   908 => (x"87",x"d0",x"ff",x"05"),
   909 => (x"26",x"4d",x"26",x"26"),
   910 => (x"26",x"4b",x"26",x"4c"),
   911 => (x"1e",x"4f",x"26",x"4a"),
   912 => (x"f8",x"27",x"1e",x"72"),
   913 => (x"bf",x"00",x"00",x"16"),
   914 => (x"87",x"cb",x"c0",x"02"),
   915 => (x"27",x"49",x"66",x"c8"),
   916 => (x"00",x"00",x"16",x"f8"),
   917 => (x"27",x"79",x"bf",x"bf"),
   918 => (x"00",x"00",x"16",x"f8"),
   919 => (x"82",x"cc",x"4a",x"bf"),
   920 => (x"00",x"27",x"1e",x"72"),
   921 => (x"bf",x"00",x"00",x"17"),
   922 => (x"27",x"1e",x"ca",x"1e"),
   923 => (x"00",x"00",x"03",x"16"),
   924 => (x"26",x"86",x"cc",x"0f"),
   925 => (x"1e",x"4f",x"26",x"4a"),
   926 => (x"08",x"27",x"1e",x"72"),
   927 => (x"97",x"00",x"00",x"17"),
   928 => (x"c0",x"c1",x"4a",x"bf"),
   929 => (x"92",x"c0",x"c0",x"c0"),
   930 => (x"92",x"b7",x"c0",x"c4"),
   931 => (x"b7",x"c1",x"c1",x"4a"),
   932 => (x"c5",x"c0",x"02",x"aa"),
   933 => (x"c0",x"4a",x"c0",x"87"),
   934 => (x"4a",x"c1",x"87",x"c2"),
   935 => (x"00",x"17",x"04",x"27"),
   936 => (x"72",x"48",x"bf",x"00"),
   937 => (x"17",x"08",x"27",x"b0"),
   938 => (x"27",x"58",x"00",x"00"),
   939 => (x"00",x"00",x"17",x"09"),
   940 => (x"51",x"c2",x"c1",x"49"),
   941 => (x"4f",x"26",x"4a",x"26"),
   942 => (x"17",x"08",x"27",x"1e"),
   943 => (x"c1",x"49",x"00",x"00"),
   944 => (x"04",x"27",x"51",x"c1"),
   945 => (x"49",x"00",x"00",x"17"),
   946 => (x"4f",x"26",x"79",x"c0"),
   947 => (x"33",x"32",x"31",x"30"),
   948 => (x"37",x"36",x"35",x"34"),
   949 => (x"42",x"41",x"39",x"38"),
   950 => (x"46",x"45",x"44",x"43"),
   951 => (x"6f",x"72",x"50",x"00"),
   952 => (x"6d",x"61",x"72",x"67"),
   953 => (x"6d",x"6f",x"63",x"20"),
   954 => (x"65",x"6c",x"69",x"70"),
   955 => (x"69",x"77",x"20",x"64"),
   956 => (x"27",x"20",x"68",x"74"),
   957 => (x"69",x"67",x"65",x"72"),
   958 => (x"72",x"65",x"74",x"73"),
   959 => (x"74",x"61",x"20",x"27"),
   960 => (x"62",x"69",x"72",x"74"),
   961 => (x"0a",x"65",x"74",x"75"),
   962 => (x"50",x"00",x"0a",x"00"),
   963 => (x"72",x"67",x"6f",x"72"),
   964 => (x"63",x"20",x"6d",x"61"),
   965 => (x"69",x"70",x"6d",x"6f"),
   966 => (x"20",x"64",x"65",x"6c"),
   967 => (x"68",x"74",x"69",x"77"),
   968 => (x"20",x"74",x"75",x"6f"),
   969 => (x"67",x"65",x"72",x"27"),
   970 => (x"65",x"74",x"73",x"69"),
   971 => (x"61",x"20",x"27",x"72"),
   972 => (x"69",x"72",x"74",x"74"),
   973 => (x"65",x"74",x"75",x"62"),
   974 => (x"00",x"0a",x"00",x"0a"),
   975 => (x"59",x"52",x"48",x"44"),
   976 => (x"4e",x"4f",x"54",x"53"),
   977 => (x"52",x"50",x"20",x"45"),
   978 => (x"41",x"52",x"47",x"4f"),
   979 => (x"33",x"20",x"2c",x"4d"),
   980 => (x"20",x"44",x"52",x"27"),
   981 => (x"49",x"52",x"54",x"53"),
   982 => (x"44",x"00",x"47",x"4e"),
   983 => (x"53",x"59",x"52",x"48"),
   984 => (x"45",x"4e",x"4f",x"54"),
   985 => (x"4f",x"52",x"50",x"20"),
   986 => (x"4d",x"41",x"52",x"47"),
   987 => (x"27",x"32",x"20",x"2c"),
   988 => (x"53",x"20",x"44",x"4e"),
   989 => (x"4e",x"49",x"52",x"54"),
   990 => (x"65",x"4d",x"00",x"47"),
   991 => (x"72",x"75",x"73",x"61"),
   992 => (x"74",x"20",x"64",x"65"),
   993 => (x"20",x"65",x"6d",x"69"),
   994 => (x"20",x"6f",x"6f",x"74"),
   995 => (x"6c",x"61",x"6d",x"73"),
   996 => (x"6f",x"74",x"20",x"6c"),
   997 => (x"74",x"62",x"6f",x"20"),
   998 => (x"20",x"6e",x"69",x"61"),
   999 => (x"6e",x"61",x"65",x"6d"),
  1000 => (x"66",x"67",x"6e",x"69"),
  1001 => (x"72",x"20",x"6c",x"75"),
  1002 => (x"6c",x"75",x"73",x"65"),
  1003 => (x"00",x"0a",x"73",x"74"),
  1004 => (x"61",x"65",x"6c",x"50"),
  1005 => (x"69",x"20",x"65",x"73"),
  1006 => (x"65",x"72",x"63",x"6e"),
  1007 => (x"20",x"65",x"73",x"61"),
  1008 => (x"62",x"6d",x"75",x"6e"),
  1009 => (x"6f",x"20",x"72",x"65"),
  1010 => (x"75",x"72",x"20",x"66"),
  1011 => (x"00",x"0a",x"73",x"6e"),
  1012 => (x"69",x"4d",x"00",x"0a"),
  1013 => (x"73",x"6f",x"72",x"63"),
  1014 => (x"6e",x"6f",x"63",x"65"),
  1015 => (x"66",x"20",x"73",x"64"),
  1016 => (x"6f",x"20",x"72",x"6f"),
  1017 => (x"72",x"20",x"65",x"6e"),
  1018 => (x"74",x"20",x"6e",x"75"),
  1019 => (x"75",x"6f",x"72",x"68"),
  1020 => (x"44",x"20",x"68",x"67"),
  1021 => (x"73",x"79",x"72",x"68"),
  1022 => (x"65",x"6e",x"6f",x"74"),
  1023 => (x"25",x"00",x"20",x"3a"),
  1024 => (x"00",x"0a",x"20",x"64"),
  1025 => (x"79",x"72",x"68",x"44"),
  1026 => (x"6e",x"6f",x"74",x"73"),
  1027 => (x"70",x"20",x"73",x"65"),
  1028 => (x"53",x"20",x"72",x"65"),
  1029 => (x"6e",x"6f",x"63",x"65"),
  1030 => (x"20",x"20",x"3a",x"64"),
  1031 => (x"20",x"20",x"20",x"20"),
  1032 => (x"20",x"20",x"20",x"20"),
  1033 => (x"20",x"20",x"20",x"20"),
  1034 => (x"20",x"20",x"20",x"20"),
  1035 => (x"20",x"20",x"20",x"20"),
  1036 => (x"20",x"64",x"25",x"00"),
  1037 => (x"41",x"56",x"00",x"0a"),
  1038 => (x"49",x"4d",x"20",x"58"),
  1039 => (x"72",x"20",x"53",x"50"),
  1040 => (x"6e",x"69",x"74",x"61"),
  1041 => (x"20",x"2a",x"20",x"67"),
  1042 => (x"30",x"30",x"30",x"31"),
  1043 => (x"25",x"20",x"3d",x"20"),
  1044 => (x"00",x"0a",x"20",x"64"),
  1045 => (x"48",x"44",x"00",x"0a"),
  1046 => (x"54",x"53",x"59",x"52"),
  1047 => (x"20",x"45",x"4e",x"4f"),
  1048 => (x"47",x"4f",x"52",x"50"),
  1049 => (x"2c",x"4d",x"41",x"52"),
  1050 => (x"4d",x"4f",x"53",x"20"),
  1051 => (x"54",x"53",x"20",x"45"),
  1052 => (x"47",x"4e",x"49",x"52"),
  1053 => (x"52",x"48",x"44",x"00"),
  1054 => (x"4f",x"54",x"53",x"59"),
  1055 => (x"50",x"20",x"45",x"4e"),
  1056 => (x"52",x"47",x"4f",x"52"),
  1057 => (x"20",x"2c",x"4d",x"41"),
  1058 => (x"54",x"53",x"27",x"31"),
  1059 => (x"52",x"54",x"53",x"20"),
  1060 => (x"00",x"47",x"4e",x"49"),
  1061 => (x"68",x"44",x"00",x"0a"),
  1062 => (x"74",x"73",x"79",x"72"),
  1063 => (x"20",x"65",x"6e",x"6f"),
  1064 => (x"63",x"6e",x"65",x"42"),
  1065 => (x"72",x"61",x"6d",x"68"),
  1066 => (x"56",x"20",x"2c",x"6b"),
  1067 => (x"69",x"73",x"72",x"65"),
  1068 => (x"32",x"20",x"6e",x"6f"),
  1069 => (x"28",x"20",x"31",x"2e"),
  1070 => (x"67",x"6e",x"61",x"4c"),
  1071 => (x"65",x"67",x"61",x"75"),
  1072 => (x"29",x"43",x"20",x"3a"),
  1073 => (x"00",x"0a",x"00",x"0a"),
  1074 => (x"63",x"65",x"78",x"45"),
  1075 => (x"6f",x"69",x"74",x"75"),
  1076 => (x"74",x"73",x"20",x"6e"),
  1077 => (x"73",x"74",x"72",x"61"),
  1078 => (x"64",x"25",x"20",x"2c"),
  1079 => (x"6e",x"75",x"72",x"20"),
  1080 => (x"68",x"74",x"20",x"73"),
  1081 => (x"67",x"75",x"6f",x"72"),
  1082 => (x"68",x"44",x"20",x"68"),
  1083 => (x"74",x"73",x"79",x"72"),
  1084 => (x"0a",x"65",x"6e",x"6f"),
  1085 => (x"65",x"78",x"45",x"00"),
  1086 => (x"69",x"74",x"75",x"63"),
  1087 => (x"65",x"20",x"6e",x"6f"),
  1088 => (x"0a",x"73",x"64",x"6e"),
  1089 => (x"46",x"00",x"0a",x"00"),
  1090 => (x"6c",x"61",x"6e",x"69"),
  1091 => (x"6c",x"61",x"76",x"20"),
  1092 => (x"20",x"73",x"65",x"75"),
  1093 => (x"74",x"20",x"66",x"6f"),
  1094 => (x"76",x"20",x"65",x"68"),
  1095 => (x"61",x"69",x"72",x"61"),
  1096 => (x"73",x"65",x"6c",x"62"),
  1097 => (x"65",x"73",x"75",x"20"),
  1098 => (x"6e",x"69",x"20",x"64"),
  1099 => (x"65",x"68",x"74",x"20"),
  1100 => (x"6e",x"65",x"62",x"20"),
  1101 => (x"61",x"6d",x"68",x"63"),
  1102 => (x"0a",x"3a",x"6b",x"72"),
  1103 => (x"49",x"00",x"0a",x"00"),
  1104 => (x"47",x"5f",x"74",x"6e"),
  1105 => (x"3a",x"62",x"6f",x"6c"),
  1106 => (x"20",x"20",x"20",x"20"),
  1107 => (x"20",x"20",x"20",x"20"),
  1108 => (x"20",x"20",x"20",x"20"),
  1109 => (x"00",x"0a",x"64",x"25"),
  1110 => (x"20",x"20",x"20",x"20"),
  1111 => (x"20",x"20",x"20",x"20"),
  1112 => (x"75",x"6f",x"68",x"73"),
  1113 => (x"62",x"20",x"64",x"6c"),
  1114 => (x"20",x"20",x"3a",x"65"),
  1115 => (x"0a",x"64",x"25",x"20"),
  1116 => (x"6f",x"6f",x"42",x"00"),
  1117 => (x"6c",x"47",x"5f",x"6c"),
  1118 => (x"20",x"3a",x"62",x"6f"),
  1119 => (x"20",x"20",x"20",x"20"),
  1120 => (x"20",x"20",x"20",x"20"),
  1121 => (x"64",x"25",x"20",x"20"),
  1122 => (x"20",x"20",x"00",x"0a"),
  1123 => (x"20",x"20",x"20",x"20"),
  1124 => (x"68",x"73",x"20",x"20"),
  1125 => (x"64",x"6c",x"75",x"6f"),
  1126 => (x"3a",x"65",x"62",x"20"),
  1127 => (x"25",x"20",x"20",x"20"),
  1128 => (x"43",x"00",x"0a",x"64"),
  1129 => (x"5f",x"31",x"5f",x"68"),
  1130 => (x"62",x"6f",x"6c",x"47"),
  1131 => (x"20",x"20",x"20",x"3a"),
  1132 => (x"20",x"20",x"20",x"20"),
  1133 => (x"20",x"20",x"20",x"20"),
  1134 => (x"00",x"0a",x"63",x"25"),
  1135 => (x"20",x"20",x"20",x"20"),
  1136 => (x"20",x"20",x"20",x"20"),
  1137 => (x"75",x"6f",x"68",x"73"),
  1138 => (x"62",x"20",x"64",x"6c"),
  1139 => (x"20",x"20",x"3a",x"65"),
  1140 => (x"0a",x"63",x"25",x"20"),
  1141 => (x"5f",x"68",x"43",x"00"),
  1142 => (x"6c",x"47",x"5f",x"32"),
  1143 => (x"20",x"3a",x"62",x"6f"),
  1144 => (x"20",x"20",x"20",x"20"),
  1145 => (x"20",x"20",x"20",x"20"),
  1146 => (x"63",x"25",x"20",x"20"),
  1147 => (x"20",x"20",x"00",x"0a"),
  1148 => (x"20",x"20",x"20",x"20"),
  1149 => (x"68",x"73",x"20",x"20"),
  1150 => (x"64",x"6c",x"75",x"6f"),
  1151 => (x"3a",x"65",x"62",x"20"),
  1152 => (x"25",x"20",x"20",x"20"),
  1153 => (x"41",x"00",x"0a",x"63"),
  1154 => (x"31",x"5f",x"72",x"72"),
  1155 => (x"6f",x"6c",x"47",x"5f"),
  1156 => (x"5d",x"38",x"5b",x"62"),
  1157 => (x"20",x"20",x"20",x"3a"),
  1158 => (x"20",x"20",x"20",x"20"),
  1159 => (x"00",x"0a",x"64",x"25"),
  1160 => (x"20",x"20",x"20",x"20"),
  1161 => (x"20",x"20",x"20",x"20"),
  1162 => (x"75",x"6f",x"68",x"73"),
  1163 => (x"62",x"20",x"64",x"6c"),
  1164 => (x"20",x"20",x"3a",x"65"),
  1165 => (x"0a",x"64",x"25",x"20"),
  1166 => (x"72",x"72",x"41",x"00"),
  1167 => (x"47",x"5f",x"32",x"5f"),
  1168 => (x"5b",x"62",x"6f",x"6c"),
  1169 => (x"37",x"5b",x"5d",x"38"),
  1170 => (x"20",x"20",x"3a",x"5d"),
  1171 => (x"64",x"25",x"20",x"20"),
  1172 => (x"20",x"20",x"00",x"0a"),
  1173 => (x"20",x"20",x"20",x"20"),
  1174 => (x"68",x"73",x"20",x"20"),
  1175 => (x"64",x"6c",x"75",x"6f"),
  1176 => (x"3a",x"65",x"62",x"20"),
  1177 => (x"4e",x"20",x"20",x"20"),
  1178 => (x"65",x"62",x"6d",x"75"),
  1179 => (x"66",x"4f",x"5f",x"72"),
  1180 => (x"6e",x"75",x"52",x"5f"),
  1181 => (x"20",x"2b",x"20",x"73"),
  1182 => (x"00",x"0a",x"30",x"31"),
  1183 => (x"5f",x"72",x"74",x"50"),
  1184 => (x"62",x"6f",x"6c",x"47"),
  1185 => (x"00",x"0a",x"3e",x"2d"),
  1186 => (x"74",x"50",x"20",x"20"),
  1187 => (x"6f",x"43",x"5f",x"72"),
  1188 => (x"20",x"3a",x"70",x"6d"),
  1189 => (x"20",x"20",x"20",x"20"),
  1190 => (x"20",x"20",x"20",x"20"),
  1191 => (x"0a",x"64",x"25",x"20"),
  1192 => (x"20",x"20",x"20",x"00"),
  1193 => (x"20",x"20",x"20",x"20"),
  1194 => (x"6f",x"68",x"73",x"20"),
  1195 => (x"20",x"64",x"6c",x"75"),
  1196 => (x"20",x"3a",x"65",x"62"),
  1197 => (x"69",x"28",x"20",x"20"),
  1198 => (x"65",x"6c",x"70",x"6d"),
  1199 => (x"74",x"6e",x"65",x"6d"),
  1200 => (x"6f",x"69",x"74",x"61"),
  1201 => (x"65",x"64",x"2d",x"6e"),
  1202 => (x"64",x"6e",x"65",x"70"),
  1203 => (x"29",x"74",x"6e",x"65"),
  1204 => (x"20",x"20",x"00",x"0a"),
  1205 => (x"63",x"73",x"69",x"44"),
  1206 => (x"20",x"20",x"3a",x"72"),
  1207 => (x"20",x"20",x"20",x"20"),
  1208 => (x"20",x"20",x"20",x"20"),
  1209 => (x"25",x"20",x"20",x"20"),
  1210 => (x"20",x"00",x"0a",x"64"),
  1211 => (x"20",x"20",x"20",x"20"),
  1212 => (x"73",x"20",x"20",x"20"),
  1213 => (x"6c",x"75",x"6f",x"68"),
  1214 => (x"65",x"62",x"20",x"64"),
  1215 => (x"20",x"20",x"20",x"3a"),
  1216 => (x"00",x"0a",x"64",x"25"),
  1217 => (x"6e",x"45",x"20",x"20"),
  1218 => (x"43",x"5f",x"6d",x"75"),
  1219 => (x"3a",x"70",x"6d",x"6f"),
  1220 => (x"20",x"20",x"20",x"20"),
  1221 => (x"20",x"20",x"20",x"20"),
  1222 => (x"0a",x"64",x"25",x"20"),
  1223 => (x"20",x"20",x"20",x"00"),
  1224 => (x"20",x"20",x"20",x"20"),
  1225 => (x"6f",x"68",x"73",x"20"),
  1226 => (x"20",x"64",x"6c",x"75"),
  1227 => (x"20",x"3a",x"65",x"62"),
  1228 => (x"64",x"25",x"20",x"20"),
  1229 => (x"20",x"20",x"00",x"0a"),
  1230 => (x"5f",x"74",x"6e",x"49"),
  1231 => (x"70",x"6d",x"6f",x"43"),
  1232 => (x"20",x"20",x"20",x"3a"),
  1233 => (x"20",x"20",x"20",x"20"),
  1234 => (x"25",x"20",x"20",x"20"),
  1235 => (x"20",x"00",x"0a",x"64"),
  1236 => (x"20",x"20",x"20",x"20"),
  1237 => (x"73",x"20",x"20",x"20"),
  1238 => (x"6c",x"75",x"6f",x"68"),
  1239 => (x"65",x"62",x"20",x"64"),
  1240 => (x"20",x"20",x"20",x"3a"),
  1241 => (x"00",x"0a",x"64",x"25"),
  1242 => (x"74",x"53",x"20",x"20"),
  1243 => (x"6f",x"43",x"5f",x"72"),
  1244 => (x"20",x"3a",x"70",x"6d"),
  1245 => (x"20",x"20",x"20",x"20"),
  1246 => (x"20",x"20",x"20",x"20"),
  1247 => (x"0a",x"73",x"25",x"20"),
  1248 => (x"20",x"20",x"20",x"00"),
  1249 => (x"20",x"20",x"20",x"20"),
  1250 => (x"6f",x"68",x"73",x"20"),
  1251 => (x"20",x"64",x"6c",x"75"),
  1252 => (x"20",x"3a",x"65",x"62"),
  1253 => (x"48",x"44",x"20",x"20"),
  1254 => (x"54",x"53",x"59",x"52"),
  1255 => (x"20",x"45",x"4e",x"4f"),
  1256 => (x"47",x"4f",x"52",x"50"),
  1257 => (x"2c",x"4d",x"41",x"52"),
  1258 => (x"4d",x"4f",x"53",x"20"),
  1259 => (x"54",x"53",x"20",x"45"),
  1260 => (x"47",x"4e",x"49",x"52"),
  1261 => (x"65",x"4e",x"00",x"0a"),
  1262 => (x"50",x"5f",x"74",x"78"),
  1263 => (x"47",x"5f",x"72",x"74"),
  1264 => (x"2d",x"62",x"6f",x"6c"),
  1265 => (x"20",x"00",x"0a",x"3e"),
  1266 => (x"72",x"74",x"50",x"20"),
  1267 => (x"6d",x"6f",x"43",x"5f"),
  1268 => (x"20",x"20",x"3a",x"70"),
  1269 => (x"20",x"20",x"20",x"20"),
  1270 => (x"20",x"20",x"20",x"20"),
  1271 => (x"00",x"0a",x"64",x"25"),
  1272 => (x"20",x"20",x"20",x"20"),
  1273 => (x"20",x"20",x"20",x"20"),
  1274 => (x"75",x"6f",x"68",x"73"),
  1275 => (x"62",x"20",x"64",x"6c"),
  1276 => (x"20",x"20",x"3a",x"65"),
  1277 => (x"6d",x"69",x"28",x"20"),
  1278 => (x"6d",x"65",x"6c",x"70"),
  1279 => (x"61",x"74",x"6e",x"65"),
  1280 => (x"6e",x"6f",x"69",x"74"),
  1281 => (x"70",x"65",x"64",x"2d"),
  1282 => (x"65",x"64",x"6e",x"65"),
  1283 => (x"2c",x"29",x"74",x"6e"),
  1284 => (x"6d",x"61",x"73",x"20"),
  1285 => (x"73",x"61",x"20",x"65"),
  1286 => (x"6f",x"62",x"61",x"20"),
  1287 => (x"00",x"0a",x"65",x"76"),
  1288 => (x"69",x"44",x"20",x"20"),
  1289 => (x"3a",x"72",x"63",x"73"),
  1290 => (x"20",x"20",x"20",x"20"),
  1291 => (x"20",x"20",x"20",x"20"),
  1292 => (x"20",x"20",x"20",x"20"),
  1293 => (x"0a",x"64",x"25",x"20"),
  1294 => (x"20",x"20",x"20",x"00"),
  1295 => (x"20",x"20",x"20",x"20"),
  1296 => (x"6f",x"68",x"73",x"20"),
  1297 => (x"20",x"64",x"6c",x"75"),
  1298 => (x"20",x"3a",x"65",x"62"),
  1299 => (x"64",x"25",x"20",x"20"),
  1300 => (x"20",x"20",x"00",x"0a"),
  1301 => (x"6d",x"75",x"6e",x"45"),
  1302 => (x"6d",x"6f",x"43",x"5f"),
  1303 => (x"20",x"20",x"3a",x"70"),
  1304 => (x"20",x"20",x"20",x"20"),
  1305 => (x"25",x"20",x"20",x"20"),
  1306 => (x"20",x"00",x"0a",x"64"),
  1307 => (x"20",x"20",x"20",x"20"),
  1308 => (x"73",x"20",x"20",x"20"),
  1309 => (x"6c",x"75",x"6f",x"68"),
  1310 => (x"65",x"62",x"20",x"64"),
  1311 => (x"20",x"20",x"20",x"3a"),
  1312 => (x"00",x"0a",x"64",x"25"),
  1313 => (x"6e",x"49",x"20",x"20"),
  1314 => (x"6f",x"43",x"5f",x"74"),
  1315 => (x"20",x"3a",x"70",x"6d"),
  1316 => (x"20",x"20",x"20",x"20"),
  1317 => (x"20",x"20",x"20",x"20"),
  1318 => (x"0a",x"64",x"25",x"20"),
  1319 => (x"20",x"20",x"20",x"00"),
  1320 => (x"20",x"20",x"20",x"20"),
  1321 => (x"6f",x"68",x"73",x"20"),
  1322 => (x"20",x"64",x"6c",x"75"),
  1323 => (x"20",x"3a",x"65",x"62"),
  1324 => (x"64",x"25",x"20",x"20"),
  1325 => (x"20",x"20",x"00",x"0a"),
  1326 => (x"5f",x"72",x"74",x"53"),
  1327 => (x"70",x"6d",x"6f",x"43"),
  1328 => (x"20",x"20",x"20",x"3a"),
  1329 => (x"20",x"20",x"20",x"20"),
  1330 => (x"25",x"20",x"20",x"20"),
  1331 => (x"20",x"00",x"0a",x"73"),
  1332 => (x"20",x"20",x"20",x"20"),
  1333 => (x"73",x"20",x"20",x"20"),
  1334 => (x"6c",x"75",x"6f",x"68"),
  1335 => (x"65",x"62",x"20",x"64"),
  1336 => (x"20",x"20",x"20",x"3a"),
  1337 => (x"59",x"52",x"48",x"44"),
  1338 => (x"4e",x"4f",x"54",x"53"),
  1339 => (x"52",x"50",x"20",x"45"),
  1340 => (x"41",x"52",x"47",x"4f"),
  1341 => (x"53",x"20",x"2c",x"4d"),
  1342 => (x"20",x"45",x"4d",x"4f"),
  1343 => (x"49",x"52",x"54",x"53"),
  1344 => (x"00",x"0a",x"47",x"4e"),
  1345 => (x"5f",x"74",x"6e",x"49"),
  1346 => (x"6f",x"4c",x"5f",x"31"),
  1347 => (x"20",x"20",x"3a",x"63"),
  1348 => (x"20",x"20",x"20",x"20"),
  1349 => (x"20",x"20",x"20",x"20"),
  1350 => (x"0a",x"64",x"25",x"20"),
  1351 => (x"20",x"20",x"20",x"00"),
  1352 => (x"20",x"20",x"20",x"20"),
  1353 => (x"6f",x"68",x"73",x"20"),
  1354 => (x"20",x"64",x"6c",x"75"),
  1355 => (x"20",x"3a",x"65",x"62"),
  1356 => (x"64",x"25",x"20",x"20"),
  1357 => (x"6e",x"49",x"00",x"0a"),
  1358 => (x"5f",x"32",x"5f",x"74"),
  1359 => (x"3a",x"63",x"6f",x"4c"),
  1360 => (x"20",x"20",x"20",x"20"),
  1361 => (x"20",x"20",x"20",x"20"),
  1362 => (x"25",x"20",x"20",x"20"),
  1363 => (x"20",x"00",x"0a",x"64"),
  1364 => (x"20",x"20",x"20",x"20"),
  1365 => (x"73",x"20",x"20",x"20"),
  1366 => (x"6c",x"75",x"6f",x"68"),
  1367 => (x"65",x"62",x"20",x"64"),
  1368 => (x"20",x"20",x"20",x"3a"),
  1369 => (x"00",x"0a",x"64",x"25"),
  1370 => (x"5f",x"74",x"6e",x"49"),
  1371 => (x"6f",x"4c",x"5f",x"33"),
  1372 => (x"20",x"20",x"3a",x"63"),
  1373 => (x"20",x"20",x"20",x"20"),
  1374 => (x"20",x"20",x"20",x"20"),
  1375 => (x"0a",x"64",x"25",x"20"),
  1376 => (x"20",x"20",x"20",x"00"),
  1377 => (x"20",x"20",x"20",x"20"),
  1378 => (x"6f",x"68",x"73",x"20"),
  1379 => (x"20",x"64",x"6c",x"75"),
  1380 => (x"20",x"3a",x"65",x"62"),
  1381 => (x"64",x"25",x"20",x"20"),
  1382 => (x"6e",x"45",x"00",x"0a"),
  1383 => (x"4c",x"5f",x"6d",x"75"),
  1384 => (x"20",x"3a",x"63",x"6f"),
  1385 => (x"20",x"20",x"20",x"20"),
  1386 => (x"20",x"20",x"20",x"20"),
  1387 => (x"25",x"20",x"20",x"20"),
  1388 => (x"20",x"00",x"0a",x"64"),
  1389 => (x"20",x"20",x"20",x"20"),
  1390 => (x"73",x"20",x"20",x"20"),
  1391 => (x"6c",x"75",x"6f",x"68"),
  1392 => (x"65",x"62",x"20",x"64"),
  1393 => (x"20",x"20",x"20",x"3a"),
  1394 => (x"00",x"0a",x"64",x"25"),
  1395 => (x"5f",x"72",x"74",x"53"),
  1396 => (x"6f",x"4c",x"5f",x"31"),
  1397 => (x"20",x"20",x"3a",x"63"),
  1398 => (x"20",x"20",x"20",x"20"),
  1399 => (x"20",x"20",x"20",x"20"),
  1400 => (x"0a",x"73",x"25",x"20"),
  1401 => (x"20",x"20",x"20",x"00"),
  1402 => (x"20",x"20",x"20",x"20"),
  1403 => (x"6f",x"68",x"73",x"20"),
  1404 => (x"20",x"64",x"6c",x"75"),
  1405 => (x"20",x"3a",x"65",x"62"),
  1406 => (x"48",x"44",x"20",x"20"),
  1407 => (x"54",x"53",x"59",x"52"),
  1408 => (x"20",x"45",x"4e",x"4f"),
  1409 => (x"47",x"4f",x"52",x"50"),
  1410 => (x"2c",x"4d",x"41",x"52"),
  1411 => (x"53",x"27",x"31",x"20"),
  1412 => (x"54",x"53",x"20",x"54"),
  1413 => (x"47",x"4e",x"49",x"52"),
  1414 => (x"74",x"53",x"00",x"0a"),
  1415 => (x"5f",x"32",x"5f",x"72"),
  1416 => (x"3a",x"63",x"6f",x"4c"),
  1417 => (x"20",x"20",x"20",x"20"),
  1418 => (x"20",x"20",x"20",x"20"),
  1419 => (x"25",x"20",x"20",x"20"),
  1420 => (x"20",x"00",x"0a",x"73"),
  1421 => (x"20",x"20",x"20",x"20"),
  1422 => (x"73",x"20",x"20",x"20"),
  1423 => (x"6c",x"75",x"6f",x"68"),
  1424 => (x"65",x"62",x"20",x"64"),
  1425 => (x"20",x"20",x"20",x"3a"),
  1426 => (x"59",x"52",x"48",x"44"),
  1427 => (x"4e",x"4f",x"54",x"53"),
  1428 => (x"52",x"50",x"20",x"45"),
  1429 => (x"41",x"52",x"47",x"4f"),
  1430 => (x"32",x"20",x"2c",x"4d"),
  1431 => (x"20",x"44",x"4e",x"27"),
  1432 => (x"49",x"52",x"54",x"53"),
  1433 => (x"00",x"0a",x"47",x"4e"),
  1434 => (x"73",x"55",x"00",x"0a"),
  1435 => (x"74",x"20",x"72",x"65"),
  1436 => (x"3a",x"65",x"6d",x"69"),
  1437 => (x"0a",x"64",x"25",x"20"),
  1438 => (x"00",x"00",x"00",x"00"),
  1439 => (x"00",x"00",x"00",x"00"),
  1440 => (x"00",x"00",x"61",x"a8"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
