package Board_Config is
	constant Board_HaveSDRAM : boolean := false;
	constant Board_SDRAM_RowBits : integer := 13;
	constant Board_SDRAM_ColBits : integer := 9;
	constant Board_VGA_Bits : integer := 6;
	constant Board_JTAG_Uart : boolean = false;
end package;

