
package Toplevel_Config is
	constant Toplevel_UseSDRAM : boolean := true;
	constant Toplevel_SDRAMWidth : integer := 32;
	constant Toplevel_UseUART : boolean := true;
	constant Toplevel_UseVGA : boolean := true;
	constant Toplevel_UseAudio : boolean := true;
	constant Toplevel_Frequency :  integer := 120;
end package;
