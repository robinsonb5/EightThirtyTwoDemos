
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"d7",x"01"),
     1 => (x"58",x"0e",x"87",x"da"),
     2 => (x"27",x"0e",x"59",x"5e"),
     3 => (x"00",x"00",x"00",x"41"),
     4 => (x"26",x"49",x"26",x"0f"),
     5 => (x"26",x"80",x"ff",x"48"),
     6 => (x"26",x"27",x"4f",x"08"),
     7 => (x"4f",x"00",x"00",x"00"),
     8 => (x"00",x"00",x"33",x"27"),
     9 => (x"c0",x"c2",x"4f",x"00"),
    10 => (x"00",x"27",x"4e",x"c0"),
    11 => (x"0f",x"00",x"00",x"16"),
    12 => (x"c1",x"87",x"fd",x"00"),
    13 => (x"27",x"4e",x"c0",x"f0"),
    14 => (x"00",x"00",x"00",x"40"),
    15 => (x"87",x"fd",x"00",x"0f"),
    16 => (x"72",x"1e",x"4f",x"4f"),
    17 => (x"c0",x"ff",x"1e",x"1e"),
    18 => (x"c4",x"48",x"6a",x"4a"),
    19 => (x"a6",x"c4",x"98",x"c0"),
    20 => (x"ff",x"02",x"6e",x"58"),
    21 => (x"66",x"cc",x"87",x"f3"),
    22 => (x"48",x"66",x"cc",x"7a"),
    23 => (x"26",x"4a",x"26",x"26"),
    24 => (x"5a",x"5e",x"0e",x"4f"),
    25 => (x"0e",x"5d",x"5c",x"5b"),
    26 => (x"c0",x"4b",x"66",x"d4"),
    27 => (x"74",x"4c",x"13",x"4d"),
    28 => (x"d6",x"c0",x"02",x"9c"),
    29 => (x"72",x"4a",x"74",x"87"),
    30 => (x"00",x"42",x"27",x"1e"),
    31 => (x"c4",x"0f",x"00",x"00"),
    32 => (x"13",x"85",x"c1",x"86"),
    33 => (x"05",x"9c",x"74",x"4c"),
    34 => (x"75",x"87",x"ea",x"ff"),
    35 => (x"26",x"4d",x"26",x"48"),
    36 => (x"26",x"4b",x"26",x"4c"),
    37 => (x"0e",x"4f",x"26",x"4a"),
    38 => (x"5c",x"5b",x"5a",x"5e"),
    39 => (x"8e",x"d0",x"0e",x"5d"),
    40 => (x"a6",x"c4",x"4c",x"c0"),
    41 => (x"c0",x"79",x"c0",x"49"),
    42 => (x"c0",x"4b",x"a6",x"e8"),
    43 => (x"c0",x"4a",x"66",x"e4"),
    44 => (x"c1",x"48",x"66",x"e4"),
    45 => (x"a6",x"e8",x"c0",x"80"),
    46 => (x"c1",x"48",x"12",x"58"),
    47 => (x"c0",x"c0",x"c0",x"c0"),
    48 => (x"b7",x"c0",x"c4",x"90"),
    49 => (x"a6",x"c4",x"48",x"90"),
    50 => (x"c5",x"02",x"6e",x"58"),
    51 => (x"66",x"c4",x"87",x"c2"),
    52 => (x"87",x"fe",x"c3",x"02"),
    53 => (x"c0",x"49",x"a6",x"c4"),
    54 => (x"6e",x"4a",x"6e",x"79"),
    55 => (x"a9",x"f0",x"c0",x"49"),
    56 => (x"87",x"c4",x"c3",x"02"),
    57 => (x"02",x"aa",x"e3",x"c1"),
    58 => (x"c1",x"87",x"c5",x"c3"),
    59 => (x"c0",x"02",x"aa",x"e4"),
    60 => (x"ec",x"c1",x"87",x"e3"),
    61 => (x"ef",x"c2",x"02",x"aa"),
    62 => (x"aa",x"f0",x"c1",x"87"),
    63 => (x"87",x"d5",x"c0",x"02"),
    64 => (x"02",x"aa",x"f3",x"c1"),
    65 => (x"c1",x"87",x"c8",x"c2"),
    66 => (x"c0",x"02",x"aa",x"f5"),
    67 => (x"f8",x"c1",x"87",x"c7"),
    68 => (x"f0",x"c2",x"05",x"aa"),
    69 => (x"73",x"83",x"c4",x"87"),
    70 => (x"76",x"8a",x"c4",x"4a"),
    71 => (x"6e",x"79",x"6a",x"49"),
    72 => (x"87",x"db",x"c1",x"02"),
    73 => (x"c0",x"49",x"a6",x"c8"),
    74 => (x"49",x"a6",x"cc",x"79"),
    75 => (x"4a",x"6e",x"79",x"c0"),
    76 => (x"72",x"2a",x"b7",x"dc"),
    77 => (x"6e",x"9d",x"cf",x"4d"),
    78 => (x"c4",x"30",x"c4",x"48"),
    79 => (x"9d",x"75",x"58",x"a6"),
    80 => (x"87",x"c5",x"c0",x"02"),
    81 => (x"c1",x"49",x"a6",x"c8"),
    82 => (x"06",x"ad",x"c9",x"79"),
    83 => (x"c0",x"87",x"c6",x"c0"),
    84 => (x"c3",x"c0",x"85",x"f7"),
    85 => (x"85",x"f0",x"c0",x"87"),
    86 => (x"c0",x"02",x"66",x"c8"),
    87 => (x"1e",x"75",x"87",x"cc"),
    88 => (x"00",x"00",x"42",x"27"),
    89 => (x"86",x"c4",x"0f",x"00"),
    90 => (x"66",x"cc",x"84",x"c1"),
    91 => (x"d0",x"80",x"c1",x"48"),
    92 => (x"66",x"cc",x"58",x"a6"),
    93 => (x"a9",x"b7",x"c8",x"49"),
    94 => (x"87",x"f2",x"fe",x"04"),
    95 => (x"c0",x"87",x"ee",x"c1"),
    96 => (x"42",x"27",x"1e",x"f0"),
    97 => (x"0f",x"00",x"00",x"00"),
    98 => (x"84",x"c1",x"86",x"c4"),
    99 => (x"c4",x"87",x"de",x"c1"),
   100 => (x"c4",x"4a",x"73",x"83"),
   101 => (x"27",x"1e",x"6a",x"8a"),
   102 => (x"00",x"00",x"00",x"61"),
   103 => (x"70",x"86",x"c4",x"0f"),
   104 => (x"72",x"4c",x"74",x"4a"),
   105 => (x"87",x"c5",x"c1",x"84"),
   106 => (x"c1",x"49",x"a6",x"c4"),
   107 => (x"87",x"fd",x"c0",x"79"),
   108 => (x"4a",x"73",x"83",x"c4"),
   109 => (x"1e",x"6a",x"8a",x"c4"),
   110 => (x"00",x"00",x"42",x"27"),
   111 => (x"86",x"c4",x"0f",x"00"),
   112 => (x"e8",x"c0",x"84",x"c1"),
   113 => (x"27",x"1e",x"6e",x"87"),
   114 => (x"00",x"00",x"00",x"42"),
   115 => (x"c0",x"86",x"c4",x"0f"),
   116 => (x"49",x"6e",x"87",x"db"),
   117 => (x"05",x"a9",x"e5",x"c0"),
   118 => (x"c4",x"87",x"c8",x"c0"),
   119 => (x"79",x"c1",x"49",x"a6"),
   120 => (x"6e",x"87",x"ca",x"c0"),
   121 => (x"00",x"42",x"27",x"1e"),
   122 => (x"c4",x"0f",x"00",x"00"),
   123 => (x"66",x"e4",x"c0",x"86"),
   124 => (x"66",x"e4",x"c0",x"4a"),
   125 => (x"c0",x"80",x"c1",x"48"),
   126 => (x"12",x"58",x"a6",x"e8"),
   127 => (x"c0",x"c0",x"c1",x"48"),
   128 => (x"c4",x"90",x"c0",x"c0"),
   129 => (x"48",x"90",x"b7",x"c0"),
   130 => (x"6e",x"58",x"a6",x"c4"),
   131 => (x"87",x"fe",x"fa",x"05"),
   132 => (x"86",x"d0",x"48",x"74"),
   133 => (x"4c",x"26",x"4d",x"26"),
   134 => (x"4a",x"26",x"4b",x"26"),
   135 => (x"00",x"00",x"4f",x"26"),
   136 => (x"75",x"1e",x"00",x"00"),
   137 => (x"4d",x"d4",x"ff",x"1e"),
   138 => (x"7d",x"49",x"ff",x"c3"),
   139 => (x"38",x"c8",x"48",x"6d"),
   140 => (x"b0",x"6d",x"7d",x"71"),
   141 => (x"7d",x"71",x"38",x"c8"),
   142 => (x"38",x"c8",x"b0",x"6d"),
   143 => (x"b0",x"6d",x"7d",x"71"),
   144 => (x"4d",x"26",x"38",x"c8"),
   145 => (x"75",x"1e",x"4f",x"26"),
   146 => (x"4d",x"d4",x"ff",x"1e"),
   147 => (x"7d",x"49",x"ff",x"c3"),
   148 => (x"30",x"c8",x"48",x"6d"),
   149 => (x"b0",x"6d",x"7d",x"71"),
   150 => (x"7d",x"71",x"30",x"c8"),
   151 => (x"30",x"c8",x"b0",x"6d"),
   152 => (x"b0",x"6d",x"7d",x"71"),
   153 => (x"4f",x"26",x"4d",x"26"),
   154 => (x"ff",x"1e",x"75",x"1e"),
   155 => (x"66",x"cc",x"4d",x"d4"),
   156 => (x"48",x"66",x"c8",x"49"),
   157 => (x"67",x"e6",x"fe",x"7d"),
   158 => (x"07",x"31",x"c9",x"02"),
   159 => (x"7d",x"09",x"39",x"d8"),
   160 => (x"7d",x"09",x"39",x"09"),
   161 => (x"7d",x"09",x"39",x"09"),
   162 => (x"7d",x"09",x"39",x"09"),
   163 => (x"7d",x"70",x"38",x"d0"),
   164 => (x"49",x"c0",x"f1",x"c9"),
   165 => (x"6d",x"48",x"ff",x"c3"),
   166 => (x"c7",x"05",x"a8",x"08"),
   167 => (x"c1",x"7d",x"08",x"87"),
   168 => (x"87",x"f3",x"05",x"89"),
   169 => (x"4f",x"26",x"4d",x"26"),
   170 => (x"49",x"d4",x"ff",x"1e"),
   171 => (x"ff",x"48",x"c8",x"c3"),
   172 => (x"fa",x"05",x"80",x"79"),
   173 => (x"0e",x"4f",x"26",x"87"),
   174 => (x"5c",x"5b",x"5a",x"5e"),
   175 => (x"ff",x"c0",x"0e",x"5d"),
   176 => (x"4d",x"f7",x"c1",x"f0"),
   177 => (x"c0",x"c0",x"c0",x"c1"),
   178 => (x"27",x"4b",x"c0",x"c0"),
   179 => (x"00",x"00",x"02",x"a8"),
   180 => (x"df",x"f8",x"c4",x"0f"),
   181 => (x"75",x"1e",x"c0",x"4c"),
   182 => (x"02",x"68",x"27",x"1e"),
   183 => (x"c8",x"0f",x"00",x"00"),
   184 => (x"c1",x"4a",x"70",x"86"),
   185 => (x"c0",x"05",x"aa",x"b7"),
   186 => (x"d4",x"ff",x"87",x"ef"),
   187 => (x"79",x"ff",x"c3",x"49"),
   188 => (x"e1",x"c0",x"1e",x"73"),
   189 => (x"1e",x"e9",x"c1",x"f0"),
   190 => (x"00",x"02",x"68",x"27"),
   191 => (x"86",x"c8",x"0f",x"00"),
   192 => (x"9a",x"72",x"4a",x"70"),
   193 => (x"87",x"cb",x"c0",x"05"),
   194 => (x"c3",x"49",x"d4",x"ff"),
   195 => (x"48",x"c1",x"79",x"ff"),
   196 => (x"27",x"87",x"d0",x"c0"),
   197 => (x"00",x"00",x"02",x"a8"),
   198 => (x"74",x"8c",x"c1",x"0f"),
   199 => (x"f4",x"fe",x"05",x"9c"),
   200 => (x"26",x"48",x"c0",x"87"),
   201 => (x"26",x"4c",x"26",x"4d"),
   202 => (x"26",x"4a",x"26",x"4b"),
   203 => (x"5a",x"5e",x"0e",x"4f"),
   204 => (x"c0",x"0e",x"5c",x"5b"),
   205 => (x"c1",x"c1",x"f0",x"ff"),
   206 => (x"49",x"d4",x"ff",x"4c"),
   207 => (x"27",x"79",x"ff",x"c3"),
   208 => (x"00",x"00",x"17",x"51"),
   209 => (x"00",x"61",x"27",x"1e"),
   210 => (x"c4",x"0f",x"00",x"00"),
   211 => (x"c0",x"4b",x"d3",x"86"),
   212 => (x"27",x"1e",x"74",x"1e"),
   213 => (x"00",x"00",x"02",x"68"),
   214 => (x"70",x"86",x"c8",x"0f"),
   215 => (x"05",x"9a",x"72",x"4a"),
   216 => (x"ff",x"87",x"cb",x"c0"),
   217 => (x"ff",x"c3",x"49",x"d4"),
   218 => (x"c0",x"48",x"c1",x"79"),
   219 => (x"a8",x"27",x"87",x"d0"),
   220 => (x"0f",x"00",x"00",x"02"),
   221 => (x"9b",x"73",x"8b",x"c1"),
   222 => (x"87",x"d3",x"ff",x"05"),
   223 => (x"4c",x"26",x"48",x"c0"),
   224 => (x"4a",x"26",x"4b",x"26"),
   225 => (x"5e",x"0e",x"4f",x"26"),
   226 => (x"5d",x"5c",x"5b",x"5a"),
   227 => (x"ff",x"c3",x"1e",x"0e"),
   228 => (x"4c",x"d4",x"ff",x"4d"),
   229 => (x"00",x"02",x"a8",x"27"),
   230 => (x"ea",x"c6",x"0f",x"00"),
   231 => (x"f0",x"e1",x"c0",x"1e"),
   232 => (x"27",x"1e",x"c8",x"c1"),
   233 => (x"00",x"00",x"02",x"68"),
   234 => (x"70",x"86",x"c8",x"0f"),
   235 => (x"27",x"1e",x"72",x"4a"),
   236 => (x"00",x"00",x"04",x"e5"),
   237 => (x"00",x"97",x"27",x"1e"),
   238 => (x"c8",x"0f",x"00",x"00"),
   239 => (x"aa",x"b7",x"c1",x"86"),
   240 => (x"87",x"cb",x"c0",x"02"),
   241 => (x"00",x"03",x"2d",x"27"),
   242 => (x"48",x"c0",x"0f",x"00"),
   243 => (x"27",x"87",x"c9",x"c3"),
   244 => (x"00",x"00",x"02",x"46"),
   245 => (x"cf",x"4a",x"70",x"0f"),
   246 => (x"c6",x"9a",x"ff",x"ff"),
   247 => (x"02",x"aa",x"b7",x"ea"),
   248 => (x"27",x"87",x"cb",x"c0"),
   249 => (x"00",x"00",x"03",x"2d"),
   250 => (x"c2",x"48",x"c0",x"0f"),
   251 => (x"7c",x"75",x"87",x"ea"),
   252 => (x"f1",x"c0",x"49",x"76"),
   253 => (x"02",x"b7",x"27",x"79"),
   254 => (x"70",x"0f",x"00",x"00"),
   255 => (x"02",x"9a",x"72",x"4a"),
   256 => (x"c0",x"87",x"eb",x"c1"),
   257 => (x"f0",x"ff",x"c0",x"1e"),
   258 => (x"27",x"1e",x"fa",x"c1"),
   259 => (x"00",x"00",x"02",x"68"),
   260 => (x"70",x"86",x"c8",x"0f"),
   261 => (x"05",x"9b",x"73",x"4b"),
   262 => (x"73",x"87",x"c3",x"c1"),
   263 => (x"04",x"a3",x"27",x"1e"),
   264 => (x"27",x"1e",x"00",x"00"),
   265 => (x"00",x"00",x"00",x"97"),
   266 => (x"75",x"86",x"c8",x"0f"),
   267 => (x"75",x"4b",x"6c",x"7c"),
   268 => (x"27",x"1e",x"73",x"9b"),
   269 => (x"00",x"00",x"04",x"af"),
   270 => (x"00",x"97",x"27",x"1e"),
   271 => (x"c8",x"0f",x"00",x"00"),
   272 => (x"75",x"7c",x"75",x"86"),
   273 => (x"75",x"7c",x"75",x"7c"),
   274 => (x"c1",x"4a",x"73",x"7c"),
   275 => (x"9a",x"72",x"9a",x"c0"),
   276 => (x"87",x"c5",x"c0",x"02"),
   277 => (x"ff",x"c0",x"48",x"c1"),
   278 => (x"c0",x"48",x"c0",x"87"),
   279 => (x"1e",x"73",x"87",x"fa"),
   280 => (x"00",x"04",x"bd",x"27"),
   281 => (x"97",x"27",x"1e",x"00"),
   282 => (x"0f",x"00",x"00",x"00"),
   283 => (x"49",x"6e",x"86",x"c8"),
   284 => (x"05",x"a9",x"b7",x"c2"),
   285 => (x"27",x"87",x"d3",x"c0"),
   286 => (x"00",x"00",x"04",x"c9"),
   287 => (x"00",x"97",x"27",x"1e"),
   288 => (x"c4",x"0f",x"00",x"00"),
   289 => (x"c0",x"48",x"c0",x"86"),
   290 => (x"48",x"6e",x"87",x"ce"),
   291 => (x"a6",x"c4",x"88",x"c1"),
   292 => (x"fd",x"05",x"6e",x"58"),
   293 => (x"48",x"c0",x"87",x"df"),
   294 => (x"26",x"4d",x"26",x"26"),
   295 => (x"26",x"4b",x"26",x"4c"),
   296 => (x"43",x"4f",x"26",x"4a"),
   297 => (x"38",x"35",x"44",x"4d"),
   298 => (x"0a",x"64",x"25",x"20"),
   299 => (x"43",x"00",x"20",x"20"),
   300 => (x"38",x"35",x"44",x"4d"),
   301 => (x"25",x"20",x"32",x"5f"),
   302 => (x"20",x"20",x"0a",x"64"),
   303 => (x"44",x"4d",x"43",x"00"),
   304 => (x"25",x"20",x"38",x"35"),
   305 => (x"20",x"20",x"0a",x"64"),
   306 => (x"48",x"44",x"53",x"00"),
   307 => (x"6e",x"49",x"20",x"43"),
   308 => (x"61",x"69",x"74",x"69"),
   309 => (x"61",x"7a",x"69",x"6c"),
   310 => (x"6e",x"6f",x"69",x"74"),
   311 => (x"72",x"72",x"65",x"20"),
   312 => (x"0a",x"21",x"72",x"6f"),
   313 => (x"64",x"6d",x"63",x"00"),
   314 => (x"44",x"4d",x"43",x"5f"),
   315 => (x"65",x"72",x"20",x"38"),
   316 => (x"6e",x"6f",x"70",x"73"),
   317 => (x"20",x"3a",x"65",x"73"),
   318 => (x"00",x"0a",x"64",x"25"),
   319 => (x"5b",x"5a",x"5e",x"0e"),
   320 => (x"1e",x"0e",x"5d",x"5c"),
   321 => (x"c8",x"4c",x"d0",x"ff"),
   322 => (x"27",x"4b",x"c0",x"c0"),
   323 => (x"00",x"00",x"02",x"1e"),
   324 => (x"27",x"79",x"c1",x"49"),
   325 => (x"00",x"00",x"06",x"19"),
   326 => (x"00",x"61",x"27",x"1e"),
   327 => (x"c4",x"0f",x"00",x"00"),
   328 => (x"6c",x"4d",x"c7",x"86"),
   329 => (x"c4",x"98",x"73",x"48"),
   330 => (x"02",x"6e",x"58",x"a6"),
   331 => (x"6c",x"87",x"cc",x"c0"),
   332 => (x"c4",x"98",x"73",x"48"),
   333 => (x"05",x"6e",x"58",x"a6"),
   334 => (x"c0",x"87",x"f4",x"ff"),
   335 => (x"02",x"a8",x"27",x"7c"),
   336 => (x"6c",x"0f",x"00",x"00"),
   337 => (x"c4",x"98",x"73",x"48"),
   338 => (x"02",x"6e",x"58",x"a6"),
   339 => (x"6c",x"87",x"cc",x"c0"),
   340 => (x"c4",x"98",x"73",x"48"),
   341 => (x"05",x"6e",x"58",x"a6"),
   342 => (x"c1",x"87",x"f4",x"ff"),
   343 => (x"c0",x"1e",x"c0",x"7c"),
   344 => (x"c0",x"c1",x"d0",x"e5"),
   345 => (x"02",x"68",x"27",x"1e"),
   346 => (x"c8",x"0f",x"00",x"00"),
   347 => (x"c1",x"4a",x"70",x"86"),
   348 => (x"c0",x"05",x"aa",x"b7"),
   349 => (x"4d",x"c1",x"87",x"c2"),
   350 => (x"05",x"ad",x"b7",x"c2"),
   351 => (x"27",x"87",x"d3",x"c0"),
   352 => (x"00",x"00",x"06",x"14"),
   353 => (x"00",x"61",x"27",x"1e"),
   354 => (x"c4",x"0f",x"00",x"00"),
   355 => (x"c1",x"48",x"c0",x"86"),
   356 => (x"8d",x"c1",x"87",x"f7"),
   357 => (x"fe",x"05",x"9d",x"75"),
   358 => (x"86",x"27",x"87",x"c9"),
   359 => (x"0f",x"00",x"00",x"03"),
   360 => (x"00",x"02",x"22",x"27"),
   361 => (x"1e",x"27",x"58",x"00"),
   362 => (x"bf",x"00",x"00",x"02"),
   363 => (x"87",x"d0",x"c0",x"05"),
   364 => (x"ff",x"c0",x"1e",x"c1"),
   365 => (x"1e",x"d0",x"c1",x"f0"),
   366 => (x"00",x"02",x"68",x"27"),
   367 => (x"86",x"c8",x"0f",x"00"),
   368 => (x"c3",x"49",x"d4",x"ff"),
   369 => (x"af",x"27",x"79",x"ff"),
   370 => (x"0f",x"00",x"00",x"08"),
   371 => (x"00",x"18",x"f0",x"27"),
   372 => (x"ec",x"27",x"58",x"00"),
   373 => (x"bf",x"00",x"00",x"18"),
   374 => (x"06",x"1d",x"27",x"1e"),
   375 => (x"27",x"1e",x"00",x"00"),
   376 => (x"00",x"00",x"00",x"97"),
   377 => (x"6c",x"86",x"c8",x"0f"),
   378 => (x"c4",x"98",x"73",x"48"),
   379 => (x"02",x"6e",x"58",x"a6"),
   380 => (x"6c",x"87",x"cc",x"c0"),
   381 => (x"c4",x"98",x"73",x"48"),
   382 => (x"05",x"6e",x"58",x"a6"),
   383 => (x"c0",x"87",x"f4",x"ff"),
   384 => (x"49",x"d4",x"ff",x"7c"),
   385 => (x"c1",x"79",x"ff",x"c3"),
   386 => (x"4d",x"26",x"26",x"48"),
   387 => (x"4b",x"26",x"4c",x"26"),
   388 => (x"4f",x"26",x"4a",x"26"),
   389 => (x"52",x"52",x"45",x"49"),
   390 => (x"49",x"50",x"53",x"00"),
   391 => (x"20",x"44",x"53",x"00"),
   392 => (x"64",x"72",x"61",x"63"),
   393 => (x"7a",x"69",x"73",x"20"),
   394 => (x"73",x"69",x"20",x"65"),
   395 => (x"0a",x"64",x"25",x"20"),
   396 => (x"5a",x"5e",x"0e",x"00"),
   397 => (x"0e",x"5d",x"5c",x"5b"),
   398 => (x"4d",x"ff",x"c3",x"1e"),
   399 => (x"75",x"4c",x"d4",x"ff"),
   400 => (x"bf",x"d0",x"ff",x"7c"),
   401 => (x"c0",x"c0",x"c8",x"48"),
   402 => (x"58",x"a6",x"c4",x"98"),
   403 => (x"d2",x"c0",x"02",x"6e"),
   404 => (x"c0",x"c0",x"c8",x"87"),
   405 => (x"bf",x"d0",x"ff",x"4a"),
   406 => (x"c4",x"98",x"72",x"48"),
   407 => (x"05",x"6e",x"58",x"a6"),
   408 => (x"ff",x"87",x"f2",x"ff"),
   409 => (x"c1",x"c4",x"49",x"d0"),
   410 => (x"d8",x"7c",x"75",x"79"),
   411 => (x"ff",x"c0",x"1e",x"66"),
   412 => (x"1e",x"d8",x"c1",x"f0"),
   413 => (x"00",x"02",x"68",x"27"),
   414 => (x"86",x"c8",x"0f",x"00"),
   415 => (x"9a",x"72",x"4a",x"70"),
   416 => (x"87",x"d3",x"c0",x"02"),
   417 => (x"00",x"07",x"39",x"27"),
   418 => (x"61",x"27",x"1e",x"00"),
   419 => (x"0f",x"00",x"00",x"00"),
   420 => (x"48",x"c1",x"86",x"c4"),
   421 => (x"75",x"87",x"d7",x"c2"),
   422 => (x"7c",x"fe",x"c3",x"7c"),
   423 => (x"79",x"c0",x"49",x"76"),
   424 => (x"4a",x"bf",x"66",x"dc"),
   425 => (x"b7",x"d8",x"4b",x"72"),
   426 => (x"75",x"48",x"73",x"2b"),
   427 => (x"72",x"7c",x"70",x"98"),
   428 => (x"2b",x"b7",x"d0",x"4b"),
   429 => (x"98",x"75",x"48",x"73"),
   430 => (x"4b",x"72",x"7c",x"70"),
   431 => (x"73",x"2b",x"b7",x"c8"),
   432 => (x"70",x"98",x"75",x"48"),
   433 => (x"75",x"48",x"72",x"7c"),
   434 => (x"dc",x"7c",x"70",x"98"),
   435 => (x"80",x"c4",x"48",x"66"),
   436 => (x"58",x"a6",x"e0",x"c0"),
   437 => (x"80",x"c1",x"48",x"6e"),
   438 => (x"6e",x"58",x"a6",x"c4"),
   439 => (x"b7",x"c0",x"c2",x"49"),
   440 => (x"fb",x"fe",x"04",x"a9"),
   441 => (x"75",x"7c",x"75",x"87"),
   442 => (x"d8",x"7c",x"75",x"7c"),
   443 => (x"75",x"4b",x"e0",x"da"),
   444 => (x"75",x"4a",x"6c",x"7c"),
   445 => (x"05",x"9a",x"72",x"9a"),
   446 => (x"c1",x"87",x"c8",x"c0"),
   447 => (x"05",x"9b",x"73",x"8b"),
   448 => (x"75",x"87",x"ec",x"ff"),
   449 => (x"bf",x"d0",x"ff",x"7c"),
   450 => (x"c0",x"c0",x"c8",x"48"),
   451 => (x"58",x"a6",x"c4",x"98"),
   452 => (x"d2",x"c0",x"02",x"6e"),
   453 => (x"c0",x"c0",x"c8",x"87"),
   454 => (x"bf",x"d0",x"ff",x"4a"),
   455 => (x"c4",x"98",x"72",x"48"),
   456 => (x"05",x"6e",x"58",x"a6"),
   457 => (x"ff",x"87",x"f2",x"ff"),
   458 => (x"79",x"c0",x"49",x"d0"),
   459 => (x"26",x"26",x"48",x"c0"),
   460 => (x"26",x"4c",x"26",x"4d"),
   461 => (x"26",x"4a",x"26",x"4b"),
   462 => (x"69",x"72",x"57",x"4f"),
   463 => (x"66",x"20",x"65",x"74"),
   464 => (x"65",x"6c",x"69",x"61"),
   465 => (x"0e",x"00",x"0a",x"64"),
   466 => (x"5c",x"5b",x"5a",x"5e"),
   467 => (x"d8",x"1e",x"0e",x"5d"),
   468 => (x"66",x"dc",x"4c",x"66"),
   469 => (x"c0",x"49",x"76",x"4b"),
   470 => (x"cd",x"ee",x"c5",x"79"),
   471 => (x"d4",x"ff",x"4d",x"df"),
   472 => (x"79",x"ff",x"c3",x"49"),
   473 => (x"4a",x"bf",x"d4",x"ff"),
   474 => (x"c3",x"9a",x"ff",x"c3"),
   475 => (x"05",x"aa",x"b7",x"fe"),
   476 => (x"27",x"87",x"e5",x"c1"),
   477 => (x"00",x"00",x"18",x"e8"),
   478 => (x"c4",x"79",x"c0",x"49"),
   479 => (x"c0",x"04",x"ab",x"b7"),
   480 => (x"22",x"27",x"87",x"e4"),
   481 => (x"0f",x"00",x"00",x"02"),
   482 => (x"7c",x"72",x"4a",x"70"),
   483 => (x"e8",x"27",x"84",x"c4"),
   484 => (x"bf",x"00",x"00",x"18"),
   485 => (x"27",x"80",x"72",x"48"),
   486 => (x"00",x"00",x"18",x"ec"),
   487 => (x"c4",x"8b",x"c4",x"58"),
   488 => (x"ff",x"03",x"ab",x"b7"),
   489 => (x"b7",x"c0",x"87",x"dc"),
   490 => (x"e5",x"c0",x"06",x"ab"),
   491 => (x"4d",x"d4",x"ff",x"87"),
   492 => (x"6d",x"7d",x"ff",x"c3"),
   493 => (x"7c",x"97",x"72",x"4a"),
   494 => (x"e8",x"27",x"84",x"c1"),
   495 => (x"bf",x"00",x"00",x"18"),
   496 => (x"27",x"80",x"72",x"48"),
   497 => (x"00",x"00",x"18",x"ec"),
   498 => (x"c0",x"8b",x"c1",x"58"),
   499 => (x"ff",x"01",x"ab",x"b7"),
   500 => (x"4d",x"c1",x"87",x"de"),
   501 => (x"79",x"c1",x"49",x"76"),
   502 => (x"9d",x"75",x"8d",x"c1"),
   503 => (x"87",x"fe",x"fd",x"05"),
   504 => (x"c3",x"49",x"d4",x"ff"),
   505 => (x"48",x"6e",x"79",x"ff"),
   506 => (x"26",x"4d",x"26",x"26"),
   507 => (x"26",x"4b",x"26",x"4c"),
   508 => (x"0e",x"4f",x"26",x"4a"),
   509 => (x"5c",x"5b",x"5a",x"5e"),
   510 => (x"ff",x"1e",x"0e",x"5d"),
   511 => (x"c0",x"c8",x"4b",x"d0"),
   512 => (x"4c",x"c0",x"4a",x"c0"),
   513 => (x"c3",x"49",x"d4",x"ff"),
   514 => (x"48",x"6b",x"79",x"ff"),
   515 => (x"a6",x"c4",x"98",x"72"),
   516 => (x"c0",x"02",x"6e",x"58"),
   517 => (x"48",x"6b",x"87",x"cc"),
   518 => (x"a6",x"c4",x"98",x"72"),
   519 => (x"ff",x"05",x"6e",x"58"),
   520 => (x"c1",x"c4",x"87",x"f4"),
   521 => (x"49",x"d4",x"ff",x"7b"),
   522 => (x"d8",x"79",x"ff",x"c3"),
   523 => (x"ff",x"c0",x"1e",x"66"),
   524 => (x"1e",x"d1",x"c1",x"f0"),
   525 => (x"00",x"02",x"68",x"27"),
   526 => (x"86",x"c8",x"0f",x"00"),
   527 => (x"9d",x"75",x"4d",x"70"),
   528 => (x"87",x"d6",x"c0",x"02"),
   529 => (x"66",x"dc",x"1e",x"75"),
   530 => (x"08",x"8f",x"27",x"1e"),
   531 => (x"27",x"1e",x"00",x"00"),
   532 => (x"00",x"00",x"00",x"97"),
   533 => (x"c0",x"86",x"cc",x"0f"),
   534 => (x"c0",x"c8",x"87",x"e8"),
   535 => (x"66",x"e0",x"c0",x"1e"),
   536 => (x"87",x"e3",x"fb",x"1e"),
   537 => (x"4c",x"70",x"86",x"c8"),
   538 => (x"98",x"72",x"48",x"6b"),
   539 => (x"6e",x"58",x"a6",x"c4"),
   540 => (x"87",x"cc",x"c0",x"02"),
   541 => (x"98",x"72",x"48",x"6b"),
   542 => (x"6e",x"58",x"a6",x"c4"),
   543 => (x"87",x"f4",x"ff",x"05"),
   544 => (x"48",x"74",x"7b",x"c0"),
   545 => (x"26",x"4d",x"26",x"26"),
   546 => (x"26",x"4b",x"26",x"4c"),
   547 => (x"52",x"4f",x"26",x"4a"),
   548 => (x"20",x"64",x"61",x"65"),
   549 => (x"6d",x"6d",x"6f",x"63"),
   550 => (x"20",x"64",x"6e",x"61"),
   551 => (x"6c",x"69",x"61",x"66"),
   552 => (x"61",x"20",x"64",x"65"),
   553 => (x"64",x"25",x"20",x"74"),
   554 => (x"64",x"25",x"28",x"20"),
   555 => (x"0e",x"00",x"0a",x"29"),
   556 => (x"5c",x"5b",x"5a",x"5e"),
   557 => (x"c0",x"1e",x"0e",x"5d"),
   558 => (x"f0",x"ff",x"c0",x"1e"),
   559 => (x"27",x"1e",x"c9",x"c1"),
   560 => (x"00",x"00",x"02",x"68"),
   561 => (x"d2",x"86",x"c8",x"0f"),
   562 => (x"18",x"f8",x"27",x"1e"),
   563 => (x"f9",x"1e",x"00",x"00"),
   564 => (x"86",x"c8",x"87",x"f5"),
   565 => (x"85",x"c1",x"4d",x"c0"),
   566 => (x"04",x"ad",x"b7",x"d2"),
   567 => (x"27",x"87",x"f7",x"ff"),
   568 => (x"00",x"00",x"18",x"f8"),
   569 => (x"c3",x"4a",x"bf",x"97"),
   570 => (x"c0",x"c1",x"9a",x"c0"),
   571 => (x"c0",x"05",x"aa",x"b7"),
   572 => (x"ff",x"27",x"87",x"f2"),
   573 => (x"97",x"00",x"00",x"18"),
   574 => (x"32",x"d0",x"4a",x"bf"),
   575 => (x"00",x"19",x"00",x"27"),
   576 => (x"4b",x"bf",x"97",x"00"),
   577 => (x"4a",x"72",x"33",x"c8"),
   578 => (x"01",x"27",x"b2",x"73"),
   579 => (x"97",x"00",x"00",x"19"),
   580 => (x"4a",x"72",x"4b",x"bf"),
   581 => (x"ff",x"cf",x"b2",x"73"),
   582 => (x"72",x"9a",x"ff",x"ff"),
   583 => (x"ca",x"85",x"c1",x"4d"),
   584 => (x"87",x"cb",x"c3",x"35"),
   585 => (x"00",x"19",x"01",x"27"),
   586 => (x"4a",x"bf",x"97",x"00"),
   587 => (x"9a",x"c6",x"32",x"c1"),
   588 => (x"00",x"19",x"02",x"27"),
   589 => (x"4b",x"bf",x"97",x"00"),
   590 => (x"72",x"2b",x"b7",x"c7"),
   591 => (x"27",x"b2",x"73",x"4a"),
   592 => (x"00",x"00",x"18",x"fd"),
   593 => (x"73",x"4b",x"bf",x"97"),
   594 => (x"c4",x"98",x"cf",x"48"),
   595 => (x"fe",x"27",x"58",x"a6"),
   596 => (x"97",x"00",x"00",x"18"),
   597 => (x"9b",x"c3",x"4b",x"bf"),
   598 => (x"ff",x"27",x"33",x"ca"),
   599 => (x"97",x"00",x"00",x"18"),
   600 => (x"34",x"c2",x"4c",x"bf"),
   601 => (x"b3",x"74",x"4b",x"73"),
   602 => (x"00",x"19",x"00",x"27"),
   603 => (x"4c",x"bf",x"97",x"00"),
   604 => (x"c6",x"9c",x"c0",x"c3"),
   605 => (x"4b",x"73",x"2c",x"b7"),
   606 => (x"1e",x"73",x"b3",x"74"),
   607 => (x"72",x"1e",x"66",x"c4"),
   608 => (x"09",x"fc",x"27",x"1e"),
   609 => (x"27",x"1e",x"00",x"00"),
   610 => (x"00",x"00",x"00",x"97"),
   611 => (x"c2",x"86",x"d0",x"0f"),
   612 => (x"72",x"48",x"c1",x"82"),
   613 => (x"72",x"4a",x"70",x"30"),
   614 => (x"0a",x"29",x"27",x"1e"),
   615 => (x"27",x"1e",x"00",x"00"),
   616 => (x"00",x"00",x"00",x"97"),
   617 => (x"c1",x"86",x"c8",x"0f"),
   618 => (x"c4",x"30",x"6e",x"48"),
   619 => (x"83",x"c1",x"58",x"a6"),
   620 => (x"95",x"72",x"4d",x"73"),
   621 => (x"1e",x"75",x"1e",x"6e"),
   622 => (x"00",x"0a",x"32",x"27"),
   623 => (x"97",x"27",x"1e",x"00"),
   624 => (x"0f",x"00",x"00",x"00"),
   625 => (x"49",x"6e",x"86",x"cc"),
   626 => (x"a9",x"b7",x"c0",x"c8"),
   627 => (x"87",x"cf",x"c0",x"06"),
   628 => (x"35",x"c1",x"4a",x"6e"),
   629 => (x"c8",x"2a",x"b7",x"c1"),
   630 => (x"01",x"aa",x"b7",x"c0"),
   631 => (x"75",x"87",x"f3",x"ff"),
   632 => (x"0a",x"48",x"27",x"1e"),
   633 => (x"27",x"1e",x"00",x"00"),
   634 => (x"00",x"00",x"00",x"97"),
   635 => (x"75",x"86",x"c8",x"0f"),
   636 => (x"4d",x"26",x"26",x"48"),
   637 => (x"4b",x"26",x"4c",x"26"),
   638 => (x"4f",x"26",x"4a",x"26"),
   639 => (x"69",x"73",x"5f",x"63"),
   640 => (x"6d",x"5f",x"65",x"7a"),
   641 => (x"3a",x"74",x"6c",x"75"),
   642 => (x"2c",x"64",x"25",x"20"),
   643 => (x"61",x"65",x"72",x"20"),
   644 => (x"6c",x"62",x"5f",x"64"),
   645 => (x"6e",x"65",x"6c",x"5f"),
   646 => (x"64",x"25",x"20",x"3a"),
   647 => (x"73",x"63",x"20",x"2c"),
   648 => (x"3a",x"65",x"7a",x"69"),
   649 => (x"0a",x"64",x"25",x"20"),
   650 => (x"6c",x"75",x"4d",x"00"),
   651 => (x"64",x"25",x"20",x"74"),
   652 => (x"64",x"25",x"00",x"0a"),
   653 => (x"6f",x"6c",x"62",x"20"),
   654 => (x"20",x"73",x"6b",x"63"),
   655 => (x"73",x"20",x"66",x"6f"),
   656 => (x"20",x"65",x"7a",x"69"),
   657 => (x"00",x"0a",x"64",x"25"),
   658 => (x"62",x"20",x"64",x"25"),
   659 => (x"6b",x"63",x"6f",x"6c"),
   660 => (x"66",x"6f",x"20",x"73"),
   661 => (x"32",x"31",x"35",x"20"),
   662 => (x"74",x"79",x"62",x"20"),
   663 => (x"00",x"0a",x"73",x"65"),
   664 => (x"5b",x"5a",x"5e",x"0e"),
   665 => (x"d4",x"0e",x"5d",x"5c"),
   666 => (x"4c",x"c0",x"4d",x"66"),
   667 => (x"c0",x"49",x"66",x"dc"),
   668 => (x"c0",x"06",x"a9",x"b7"),
   669 => (x"4b",x"15",x"87",x"fb"),
   670 => (x"c0",x"c0",x"c0",x"c1"),
   671 => (x"c0",x"c4",x"93",x"c0"),
   672 => (x"d8",x"4b",x"93",x"b7"),
   673 => (x"4a",x"bf",x"97",x"66"),
   674 => (x"c0",x"c0",x"c0",x"c1"),
   675 => (x"c0",x"c4",x"92",x"c0"),
   676 => (x"d8",x"4a",x"92",x"b7"),
   677 => (x"80",x"c1",x"48",x"66"),
   678 => (x"72",x"58",x"a6",x"dc"),
   679 => (x"c0",x"02",x"ab",x"b7"),
   680 => (x"48",x"c1",x"87",x"c5"),
   681 => (x"c1",x"87",x"cc",x"c0"),
   682 => (x"b7",x"66",x"dc",x"84"),
   683 => (x"c5",x"ff",x"04",x"ac"),
   684 => (x"26",x"48",x"c0",x"87"),
   685 => (x"26",x"4c",x"26",x"4d"),
   686 => (x"26",x"4a",x"26",x"4b"),
   687 => (x"5a",x"5e",x"0e",x"4f"),
   688 => (x"0e",x"5d",x"5c",x"5b"),
   689 => (x"00",x"1b",x"18",x"27"),
   690 => (x"79",x"c0",x"49",x"00"),
   691 => (x"00",x"18",x"29",x"27"),
   692 => (x"61",x"27",x"1e",x"00"),
   693 => (x"0f",x"00",x"00",x"00"),
   694 => (x"10",x"27",x"86",x"c4"),
   695 => (x"1e",x"00",x"00",x"19"),
   696 => (x"f3",x"27",x"1e",x"c0"),
   697 => (x"0f",x"00",x"00",x"07"),
   698 => (x"4a",x"70",x"86",x"c8"),
   699 => (x"c0",x"05",x"9a",x"72"),
   700 => (x"55",x"27",x"87",x"d3"),
   701 => (x"1e",x"00",x"00",x"17"),
   702 => (x"00",x"00",x"61",x"27"),
   703 => (x"86",x"c4",x"0f",x"00"),
   704 => (x"d8",x"cf",x"48",x"c0"),
   705 => (x"18",x"36",x"27",x"87"),
   706 => (x"27",x"1e",x"00",x"00"),
   707 => (x"00",x"00",x"00",x"61"),
   708 => (x"c0",x"86",x"c4",x"0f"),
   709 => (x"1b",x"44",x"27",x"4c"),
   710 => (x"c1",x"49",x"00",x"00"),
   711 => (x"27",x"1e",x"c8",x"79"),
   712 => (x"00",x"00",x"18",x"4d"),
   713 => (x"19",x"46",x"27",x"1e"),
   714 => (x"27",x"1e",x"00",x"00"),
   715 => (x"00",x"00",x"0a",x"60"),
   716 => (x"70",x"86",x"cc",x"0f"),
   717 => (x"05",x"9a",x"72",x"4a"),
   718 => (x"27",x"87",x"c8",x"c0"),
   719 => (x"00",x"00",x"1b",x"44"),
   720 => (x"c8",x"79",x"c0",x"49"),
   721 => (x"18",x"56",x"27",x"1e"),
   722 => (x"27",x"1e",x"00",x"00"),
   723 => (x"00",x"00",x"19",x"62"),
   724 => (x"0a",x"60",x"27",x"1e"),
   725 => (x"cc",x"0f",x"00",x"00"),
   726 => (x"72",x"4a",x"70",x"86"),
   727 => (x"c8",x"c0",x"05",x"9a"),
   728 => (x"1b",x"44",x"27",x"87"),
   729 => (x"c0",x"49",x"00",x"00"),
   730 => (x"1b",x"44",x"27",x"79"),
   731 => (x"1e",x"bf",x"00",x"00"),
   732 => (x"00",x"18",x"5f",x"27"),
   733 => (x"97",x"27",x"1e",x"00"),
   734 => (x"0f",x"00",x"00",x"00"),
   735 => (x"44",x"27",x"86",x"c8"),
   736 => (x"bf",x"00",x"00",x"1b"),
   737 => (x"87",x"c0",x"c3",x"02"),
   738 => (x"00",x"19",x"10",x"27"),
   739 => (x"ce",x"27",x"4d",x"00"),
   740 => (x"4b",x"00",x"00",x"1a"),
   741 => (x"00",x"1b",x"0e",x"27"),
   742 => (x"4a",x"bf",x"9f",x"00"),
   743 => (x"0e",x"27",x"1e",x"72"),
   744 => (x"4a",x"00",x"00",x"1b"),
   745 => (x"00",x"19",x"10",x"27"),
   746 => (x"1e",x"72",x"8a",x"00"),
   747 => (x"c0",x"c8",x"1e",x"d0"),
   748 => (x"17",x"87",x"27",x"1e"),
   749 => (x"27",x"1e",x"00",x"00"),
   750 => (x"00",x"00",x"00",x"97"),
   751 => (x"73",x"86",x"d4",x"0f"),
   752 => (x"6a",x"82",x"c8",x"4a"),
   753 => (x"1b",x"0e",x"27",x"4c"),
   754 => (x"bf",x"9f",x"00",x"00"),
   755 => (x"ea",x"d6",x"c5",x"4a"),
   756 => (x"c0",x"05",x"aa",x"b7"),
   757 => (x"4a",x"73",x"87",x"d3"),
   758 => (x"1e",x"6a",x"82",x"c8"),
   759 => (x"00",x"12",x"48",x"27"),
   760 => (x"86",x"c4",x"0f",x"00"),
   761 => (x"e4",x"c0",x"4c",x"70"),
   762 => (x"c7",x"4a",x"75",x"87"),
   763 => (x"6a",x"9f",x"82",x"fe"),
   764 => (x"d5",x"e9",x"ca",x"4a"),
   765 => (x"c0",x"02",x"aa",x"b7"),
   766 => (x"69",x"27",x"87",x"d3"),
   767 => (x"1e",x"00",x"00",x"17"),
   768 => (x"00",x"00",x"61",x"27"),
   769 => (x"86",x"c4",x"0f",x"00"),
   770 => (x"d0",x"cb",x"48",x"c0"),
   771 => (x"27",x"1e",x"74",x"87"),
   772 => (x"00",x"00",x"17",x"c4"),
   773 => (x"00",x"97",x"27",x"1e"),
   774 => (x"c8",x"0f",x"00",x"00"),
   775 => (x"19",x"10",x"27",x"86"),
   776 => (x"74",x"1e",x"00",x"00"),
   777 => (x"07",x"f3",x"27",x"1e"),
   778 => (x"c8",x"0f",x"00",x"00"),
   779 => (x"72",x"4a",x"70",x"86"),
   780 => (x"c5",x"c0",x"05",x"9a"),
   781 => (x"ca",x"48",x"c0",x"87"),
   782 => (x"dc",x"27",x"87",x"e3"),
   783 => (x"1e",x"00",x"00",x"17"),
   784 => (x"00",x"00",x"61",x"27"),
   785 => (x"86",x"c4",x"0f",x"00"),
   786 => (x"00",x"18",x"72",x"27"),
   787 => (x"97",x"27",x"1e",x"00"),
   788 => (x"0f",x"00",x"00",x"00"),
   789 => (x"1e",x"c8",x"86",x"c4"),
   790 => (x"00",x"18",x"8a",x"27"),
   791 => (x"62",x"27",x"1e",x"00"),
   792 => (x"1e",x"00",x"00",x"19"),
   793 => (x"00",x"0a",x"60",x"27"),
   794 => (x"86",x"cc",x"0f",x"00"),
   795 => (x"9a",x"72",x"4a",x"70"),
   796 => (x"87",x"cb",x"c0",x"05"),
   797 => (x"00",x"1b",x"18",x"27"),
   798 => (x"79",x"c1",x"49",x"00"),
   799 => (x"c8",x"87",x"f1",x"c0"),
   800 => (x"18",x"93",x"27",x"1e"),
   801 => (x"27",x"1e",x"00",x"00"),
   802 => (x"00",x"00",x"19",x"46"),
   803 => (x"0a",x"60",x"27",x"1e"),
   804 => (x"cc",x"0f",x"00",x"00"),
   805 => (x"72",x"4a",x"70",x"86"),
   806 => (x"d3",x"c0",x"02",x"9a"),
   807 => (x"18",x"03",x"27",x"87"),
   808 => (x"27",x"1e",x"00",x"00"),
   809 => (x"00",x"00",x"00",x"97"),
   810 => (x"c0",x"86",x"c4",x"0f"),
   811 => (x"87",x"ed",x"c8",x"48"),
   812 => (x"00",x"1b",x"0e",x"27"),
   813 => (x"4a",x"bf",x"97",x"00"),
   814 => (x"aa",x"b7",x"d5",x"c1"),
   815 => (x"87",x"d0",x"c0",x"05"),
   816 => (x"00",x"1b",x"0f",x"27"),
   817 => (x"4a",x"bf",x"97",x"00"),
   818 => (x"aa",x"b7",x"ea",x"c2"),
   819 => (x"87",x"c5",x"c0",x"02"),
   820 => (x"c8",x"c8",x"48",x"c0"),
   821 => (x"19",x"10",x"27",x"87"),
   822 => (x"bf",x"97",x"00",x"00"),
   823 => (x"b7",x"e9",x"c3",x"4a"),
   824 => (x"d5",x"c0",x"02",x"aa"),
   825 => (x"19",x"10",x"27",x"87"),
   826 => (x"bf",x"97",x"00",x"00"),
   827 => (x"b7",x"eb",x"c3",x"4a"),
   828 => (x"c5",x"c0",x"02",x"aa"),
   829 => (x"c7",x"48",x"c0",x"87"),
   830 => (x"1b",x"27",x"87",x"e3"),
   831 => (x"97",x"00",x"00",x"19"),
   832 => (x"9a",x"72",x"4a",x"bf"),
   833 => (x"87",x"cf",x"c0",x"05"),
   834 => (x"00",x"19",x"1c",x"27"),
   835 => (x"4a",x"bf",x"97",x"00"),
   836 => (x"02",x"aa",x"b7",x"c2"),
   837 => (x"c0",x"87",x"c5",x"c0"),
   838 => (x"87",x"c1",x"c7",x"48"),
   839 => (x"00",x"19",x"1d",x"27"),
   840 => (x"48",x"bf",x"97",x"00"),
   841 => (x"00",x"1b",x"14",x"27"),
   842 => (x"10",x"27",x"58",x"00"),
   843 => (x"bf",x"00",x"00",x"1b"),
   844 => (x"c1",x"4b",x"72",x"4a"),
   845 => (x"1b",x"14",x"27",x"8b"),
   846 => (x"73",x"49",x"00",x"00"),
   847 => (x"72",x"1e",x"73",x"79"),
   848 => (x"18",x"9c",x"27",x"1e"),
   849 => (x"27",x"1e",x"00",x"00"),
   850 => (x"00",x"00",x"00",x"97"),
   851 => (x"27",x"86",x"cc",x"0f"),
   852 => (x"00",x"00",x"19",x"1e"),
   853 => (x"74",x"4a",x"bf",x"97"),
   854 => (x"19",x"1f",x"27",x"82"),
   855 => (x"bf",x"97",x"00",x"00"),
   856 => (x"73",x"33",x"c8",x"4b"),
   857 => (x"27",x"80",x"72",x"48"),
   858 => (x"00",x"00",x"1b",x"28"),
   859 => (x"19",x"20",x"27",x"58"),
   860 => (x"bf",x"97",x"00",x"00"),
   861 => (x"1b",x"3c",x"27",x"48"),
   862 => (x"27",x"58",x"00",x"00"),
   863 => (x"00",x"00",x"1b",x"18"),
   864 => (x"df",x"c3",x"02",x"bf"),
   865 => (x"27",x"1e",x"c8",x"87"),
   866 => (x"00",x"00",x"18",x"20"),
   867 => (x"19",x"62",x"27",x"1e"),
   868 => (x"27",x"1e",x"00",x"00"),
   869 => (x"00",x"00",x"0a",x"60"),
   870 => (x"70",x"86",x"cc",x"0f"),
   871 => (x"02",x"9a",x"72",x"4a"),
   872 => (x"c0",x"87",x"c5",x"c0"),
   873 => (x"87",x"f5",x"c4",x"48"),
   874 => (x"00",x"1b",x"10",x"27"),
   875 => (x"73",x"4b",x"bf",x"00"),
   876 => (x"27",x"30",x"c4",x"48"),
   877 => (x"00",x"00",x"1b",x"40"),
   878 => (x"1b",x"34",x"27",x"58"),
   879 => (x"73",x"49",x"00",x"00"),
   880 => (x"19",x"35",x"27",x"79"),
   881 => (x"bf",x"97",x"00",x"00"),
   882 => (x"27",x"32",x"c8",x"4a"),
   883 => (x"00",x"00",x"19",x"34"),
   884 => (x"72",x"4c",x"bf",x"97"),
   885 => (x"27",x"82",x"74",x"4a"),
   886 => (x"00",x"00",x"19",x"36"),
   887 => (x"d0",x"4c",x"bf",x"97"),
   888 => (x"74",x"4a",x"72",x"34"),
   889 => (x"19",x"37",x"27",x"82"),
   890 => (x"bf",x"97",x"00",x"00"),
   891 => (x"72",x"34",x"d8",x"4c"),
   892 => (x"27",x"82",x"74",x"4a"),
   893 => (x"00",x"00",x"1b",x"40"),
   894 => (x"72",x"79",x"72",x"49"),
   895 => (x"1b",x"38",x"27",x"4a"),
   896 => (x"92",x"bf",x"00",x"00"),
   897 => (x"24",x"27",x"4a",x"72"),
   898 => (x"bf",x"00",x"00",x"1b"),
   899 => (x"1b",x"28",x"27",x"82"),
   900 => (x"72",x"49",x"00",x"00"),
   901 => (x"19",x"3d",x"27",x"79"),
   902 => (x"bf",x"97",x"00",x"00"),
   903 => (x"27",x"34",x"c8",x"4c"),
   904 => (x"00",x"00",x"19",x"3c"),
   905 => (x"74",x"4d",x"bf",x"97"),
   906 => (x"27",x"84",x"75",x"4c"),
   907 => (x"00",x"00",x"19",x"3e"),
   908 => (x"d0",x"4d",x"bf",x"97"),
   909 => (x"75",x"4c",x"74",x"35"),
   910 => (x"19",x"3f",x"27",x"84"),
   911 => (x"bf",x"97",x"00",x"00"),
   912 => (x"d8",x"9d",x"cf",x"4d"),
   913 => (x"75",x"4c",x"74",x"35"),
   914 => (x"1b",x"2c",x"27",x"84"),
   915 => (x"74",x"49",x"00",x"00"),
   916 => (x"73",x"8c",x"c2",x"79"),
   917 => (x"73",x"93",x"74",x"4b"),
   918 => (x"27",x"80",x"72",x"48"),
   919 => (x"00",x"00",x"1b",x"34"),
   920 => (x"87",x"f7",x"c1",x"58"),
   921 => (x"00",x"19",x"22",x"27"),
   922 => (x"4a",x"bf",x"97",x"00"),
   923 => (x"21",x"27",x"32",x"c8"),
   924 => (x"97",x"00",x"00",x"19"),
   925 => (x"4a",x"72",x"4b",x"bf"),
   926 => (x"3c",x"27",x"82",x"73"),
   927 => (x"49",x"00",x"00",x"1b"),
   928 => (x"32",x"c5",x"79",x"72"),
   929 => (x"c9",x"82",x"ff",x"c7"),
   930 => (x"1b",x"34",x"27",x"2a"),
   931 => (x"72",x"49",x"00",x"00"),
   932 => (x"19",x"27",x"27",x"79"),
   933 => (x"bf",x"97",x"00",x"00"),
   934 => (x"27",x"33",x"c8",x"4b"),
   935 => (x"00",x"00",x"19",x"26"),
   936 => (x"73",x"4c",x"bf",x"97"),
   937 => (x"27",x"83",x"74",x"4b"),
   938 => (x"00",x"00",x"1b",x"40"),
   939 => (x"73",x"79",x"73",x"49"),
   940 => (x"1b",x"38",x"27",x"4b"),
   941 => (x"93",x"bf",x"00",x"00"),
   942 => (x"24",x"27",x"4b",x"73"),
   943 => (x"bf",x"00",x"00",x"1b"),
   944 => (x"1b",x"30",x"27",x"83"),
   945 => (x"73",x"49",x"00",x"00"),
   946 => (x"1b",x"2c",x"27",x"79"),
   947 => (x"c0",x"49",x"00",x"00"),
   948 => (x"72",x"48",x"73",x"79"),
   949 => (x"1b",x"2c",x"27",x"80"),
   950 => (x"c1",x"58",x"00",x"00"),
   951 => (x"26",x"4d",x"26",x"48"),
   952 => (x"26",x"4b",x"26",x"4c"),
   953 => (x"0e",x"4f",x"26",x"4a"),
   954 => (x"5c",x"5b",x"5a",x"5e"),
   955 => (x"18",x"27",x"0e",x"5d"),
   956 => (x"bf",x"00",x"00",x"1b"),
   957 => (x"87",x"cf",x"c0",x"02"),
   958 => (x"c7",x"4c",x"66",x"d4"),
   959 => (x"66",x"d4",x"2c",x"b7"),
   960 => (x"9b",x"ff",x"c1",x"4b"),
   961 => (x"d4",x"87",x"cc",x"c0"),
   962 => (x"b7",x"c8",x"4c",x"66"),
   963 => (x"4b",x"66",x"d4",x"2c"),
   964 => (x"27",x"9b",x"ff",x"c3"),
   965 => (x"00",x"00",x"19",x"10"),
   966 => (x"1b",x"24",x"27",x"1e"),
   967 => (x"4a",x"bf",x"00",x"00"),
   968 => (x"1e",x"72",x"82",x"74"),
   969 => (x"00",x"07",x"f3",x"27"),
   970 => (x"86",x"c8",x"0f",x"00"),
   971 => (x"9a",x"72",x"4a",x"70"),
   972 => (x"87",x"c5",x"c0",x"05"),
   973 => (x"f2",x"c0",x"48",x"c0"),
   974 => (x"1b",x"18",x"27",x"87"),
   975 => (x"02",x"bf",x"00",x"00"),
   976 => (x"73",x"87",x"d7",x"c0"),
   977 => (x"72",x"92",x"c4",x"4a"),
   978 => (x"19",x"10",x"27",x"4a"),
   979 => (x"6a",x"82",x"00",x"00"),
   980 => (x"ff",x"ff",x"cf",x"4d"),
   981 => (x"c0",x"9d",x"ff",x"ff"),
   982 => (x"4a",x"73",x"87",x"cf"),
   983 => (x"4a",x"72",x"92",x"c2"),
   984 => (x"00",x"19",x"10",x"27"),
   985 => (x"6a",x"9f",x"82",x"00"),
   986 => (x"26",x"48",x"75",x"4d"),
   987 => (x"26",x"4c",x"26",x"4d"),
   988 => (x"26",x"4a",x"26",x"4b"),
   989 => (x"5a",x"5e",x"0e",x"4f"),
   990 => (x"0e",x"5d",x"5c",x"5b"),
   991 => (x"ff",x"cf",x"8e",x"cc"),
   992 => (x"4d",x"f8",x"ff",x"ff"),
   993 => (x"49",x"76",x"4c",x"c0"),
   994 => (x"00",x"1b",x"2c",x"27"),
   995 => (x"c4",x"79",x"bf",x"00"),
   996 => (x"30",x"27",x"49",x"a6"),
   997 => (x"bf",x"00",x"00",x"1b"),
   998 => (x"1b",x"18",x"27",x"79"),
   999 => (x"02",x"bf",x"00",x"00"),
  1000 => (x"27",x"87",x"cc",x"c0"),
  1001 => (x"00",x"00",x"1b",x"10"),
  1002 => (x"32",x"c4",x"4a",x"bf"),
  1003 => (x"27",x"87",x"c9",x"c0"),
  1004 => (x"00",x"00",x"1b",x"34"),
  1005 => (x"32",x"c4",x"4a",x"bf"),
  1006 => (x"72",x"49",x"a6",x"c8"),
  1007 => (x"c8",x"4b",x"c0",x"79"),
  1008 => (x"a9",x"c0",x"49",x"66"),
  1009 => (x"87",x"d0",x"c3",x"06"),
  1010 => (x"9a",x"cf",x"4a",x"73"),
  1011 => (x"c0",x"05",x"9a",x"72"),
  1012 => (x"10",x"27",x"87",x"e4"),
  1013 => (x"1e",x"00",x"00",x"19"),
  1014 => (x"c8",x"4a",x"66",x"c8"),
  1015 => (x"80",x"c1",x"48",x"66"),
  1016 => (x"72",x"58",x"a6",x"cc"),
  1017 => (x"07",x"f3",x"27",x"1e"),
  1018 => (x"c8",x"0f",x"00",x"00"),
  1019 => (x"19",x"10",x"27",x"86"),
  1020 => (x"c0",x"4c",x"00",x"00"),
  1021 => (x"e0",x"c0",x"87",x"c3"),
  1022 => (x"4a",x"6c",x"97",x"84"),
  1023 => (x"c2",x"02",x"9a",x"72"),
  1024 => (x"6c",x"97",x"87",x"cd"),
  1025 => (x"b7",x"e5",x"c3",x"4a"),
  1026 => (x"c2",x"c2",x"02",x"aa"),
  1027 => (x"cb",x"4a",x"74",x"87"),
  1028 => (x"4a",x"6a",x"97",x"82"),
  1029 => (x"9a",x"72",x"9a",x"d8"),
  1030 => (x"87",x"f3",x"c1",x"05"),
  1031 => (x"61",x"27",x"1e",x"74"),
  1032 => (x"0f",x"00",x"00",x"00"),
  1033 => (x"1e",x"cb",x"86",x"c4"),
  1034 => (x"1e",x"66",x"e8",x"c0"),
  1035 => (x"60",x"27",x"1e",x"74"),
  1036 => (x"0f",x"00",x"00",x"0a"),
  1037 => (x"4a",x"70",x"86",x"cc"),
  1038 => (x"c1",x"05",x"9a",x"72"),
  1039 => (x"4b",x"74",x"87",x"d1"),
  1040 => (x"e0",x"c0",x"83",x"dc"),
  1041 => (x"82",x"c4",x"4a",x"66"),
  1042 => (x"4b",x"74",x"7a",x"6b"),
  1043 => (x"e0",x"c0",x"83",x"da"),
  1044 => (x"82",x"c8",x"4a",x"66"),
  1045 => (x"70",x"48",x"6b",x"9f"),
  1046 => (x"27",x"4d",x"72",x"7a"),
  1047 => (x"00",x"00",x"1b",x"18"),
  1048 => (x"d5",x"c0",x"02",x"bf"),
  1049 => (x"d4",x"4a",x"74",x"87"),
  1050 => (x"4a",x"6a",x"9f",x"82"),
  1051 => (x"9a",x"ff",x"ff",x"c0"),
  1052 => (x"30",x"d0",x"48",x"72"),
  1053 => (x"c0",x"58",x"a6",x"c4"),
  1054 => (x"49",x"76",x"87",x"c4"),
  1055 => (x"48",x"6e",x"79",x"c0"),
  1056 => (x"7d",x"70",x"80",x"6d"),
  1057 => (x"49",x"66",x"e0",x"c0"),
  1058 => (x"48",x"c1",x"79",x"c0"),
  1059 => (x"c1",x"87",x"ce",x"c1"),
  1060 => (x"ab",x"66",x"c8",x"83"),
  1061 => (x"87",x"f0",x"fc",x"04"),
  1062 => (x"ff",x"ff",x"ff",x"cf"),
  1063 => (x"18",x"27",x"4d",x"f8"),
  1064 => (x"bf",x"00",x"00",x"1b"),
  1065 => (x"87",x"f3",x"c0",x"02"),
  1066 => (x"e7",x"27",x"1e",x"6e"),
  1067 => (x"0f",x"00",x"00",x"0e"),
  1068 => (x"a6",x"c4",x"86",x"c4"),
  1069 => (x"75",x"4a",x"6e",x"58"),
  1070 => (x"02",x"aa",x"75",x"9a"),
  1071 => (x"6e",x"87",x"dc",x"c0"),
  1072 => (x"72",x"8a",x"c2",x"4a"),
  1073 => (x"1b",x"10",x"27",x"4a"),
  1074 => (x"92",x"bf",x"00",x"00"),
  1075 => (x"00",x"1b",x"28",x"27"),
  1076 => (x"72",x"48",x"bf",x"00"),
  1077 => (x"58",x"a6",x"c8",x"80"),
  1078 => (x"c0",x"87",x"e2",x"fb"),
  1079 => (x"ff",x"ff",x"cf",x"48"),
  1080 => (x"cc",x"4d",x"f8",x"ff"),
  1081 => (x"26",x"4d",x"26",x"86"),
  1082 => (x"26",x"4b",x"26",x"4c"),
  1083 => (x"0e",x"4f",x"26",x"4a"),
  1084 => (x"0e",x"5b",x"5a",x"5e"),
  1085 => (x"4a",x"bf",x"66",x"cc"),
  1086 => (x"66",x"cc",x"82",x"c1"),
  1087 => (x"72",x"79",x"72",x"49"),
  1088 => (x"1b",x"14",x"27",x"4a"),
  1089 => (x"9a",x"bf",x"00",x"00"),
  1090 => (x"c0",x"05",x"9a",x"72"),
  1091 => (x"66",x"cc",x"87",x"d3"),
  1092 => (x"6a",x"82",x"c8",x"4a"),
  1093 => (x"0e",x"e7",x"27",x"1e"),
  1094 => (x"c4",x"0f",x"00",x"00"),
  1095 => (x"73",x"4b",x"70",x"86"),
  1096 => (x"26",x"48",x"c1",x"7a"),
  1097 => (x"26",x"4a",x"26",x"4b"),
  1098 => (x"5a",x"5e",x"0e",x"4f"),
  1099 => (x"28",x"27",x"0e",x"5b"),
  1100 => (x"bf",x"00",x"00",x"1b"),
  1101 => (x"4b",x"66",x"cc",x"4a"),
  1102 => (x"4b",x"6b",x"83",x"c8"),
  1103 => (x"4b",x"73",x"8b",x"c2"),
  1104 => (x"00",x"1b",x"10",x"27"),
  1105 => (x"72",x"93",x"bf",x"00"),
  1106 => (x"27",x"82",x"73",x"4a"),
  1107 => (x"00",x"00",x"1b",x"14"),
  1108 => (x"66",x"cc",x"4b",x"bf"),
  1109 => (x"4a",x"72",x"9b",x"bf"),
  1110 => (x"66",x"d0",x"82",x"73"),
  1111 => (x"27",x"1e",x"72",x"1e"),
  1112 => (x"00",x"00",x"07",x"f3"),
  1113 => (x"70",x"86",x"c8",x"0f"),
  1114 => (x"05",x"9a",x"72",x"4a"),
  1115 => (x"c0",x"87",x"c5",x"c0"),
  1116 => (x"87",x"c2",x"c0",x"48"),
  1117 => (x"4b",x"26",x"48",x"c1"),
  1118 => (x"4f",x"26",x"4a",x"26"),
  1119 => (x"5b",x"5a",x"5e",x"0e"),
  1120 => (x"d8",x"0e",x"5d",x"5c"),
  1121 => (x"66",x"d4",x"4c",x"66"),
  1122 => (x"1b",x"48",x"27",x"1e"),
  1123 => (x"27",x"1e",x"00",x"00"),
  1124 => (x"00",x"00",x"0f",x"75"),
  1125 => (x"70",x"86",x"c8",x"0f"),
  1126 => (x"02",x"9a",x"72",x"4a"),
  1127 => (x"27",x"87",x"df",x"c1"),
  1128 => (x"00",x"00",x"1b",x"4c"),
  1129 => (x"ff",x"c7",x"4a",x"bf"),
  1130 => (x"72",x"2a",x"c9",x"82"),
  1131 => (x"27",x"4b",x"c0",x"4d"),
  1132 => (x"00",x"00",x"12",x"20"),
  1133 => (x"00",x"61",x"27",x"1e"),
  1134 => (x"c4",x"0f",x"00",x"00"),
  1135 => (x"ad",x"b7",x"c0",x"86"),
  1136 => (x"87",x"d0",x"c1",x"06"),
  1137 => (x"48",x"27",x"1e",x"74"),
  1138 => (x"1e",x"00",x"00",x"1b"),
  1139 => (x"00",x"11",x"29",x"27"),
  1140 => (x"86",x"c8",x"0f",x"00"),
  1141 => (x"9a",x"72",x"4a",x"70"),
  1142 => (x"87",x"c5",x"c0",x"05"),
  1143 => (x"f5",x"c0",x"48",x"c0"),
  1144 => (x"1b",x"48",x"27",x"87"),
  1145 => (x"27",x"1e",x"00",x"00"),
  1146 => (x"00",x"00",x"10",x"ef"),
  1147 => (x"c8",x"86",x"c4",x"0f"),
  1148 => (x"83",x"c1",x"84",x"c0"),
  1149 => (x"04",x"ab",x"b7",x"75"),
  1150 => (x"c0",x"87",x"c9",x"ff"),
  1151 => (x"66",x"d4",x"87",x"d6"),
  1152 => (x"12",x"39",x"27",x"1e"),
  1153 => (x"27",x"1e",x"00",x"00"),
  1154 => (x"00",x"00",x"00",x"97"),
  1155 => (x"c0",x"86",x"c8",x"0f"),
  1156 => (x"87",x"c2",x"c0",x"48"),
  1157 => (x"4d",x"26",x"48",x"c1"),
  1158 => (x"4b",x"26",x"4c",x"26"),
  1159 => (x"4f",x"26",x"4a",x"26"),
  1160 => (x"6e",x"65",x"70",x"4f"),
  1161 => (x"66",x"20",x"64",x"65"),
  1162 => (x"2c",x"65",x"6c",x"69"),
  1163 => (x"61",x"6f",x"6c",x"20"),
  1164 => (x"67",x"6e",x"69",x"64"),
  1165 => (x"0a",x"2e",x"2e",x"2e"),
  1166 => (x"6e",x"61",x"43",x"00"),
  1167 => (x"6f",x"20",x"74",x"27"),
  1168 => (x"20",x"6e",x"65",x"70"),
  1169 => (x"00",x"0a",x"73",x"25"),
  1170 => (x"5b",x"5a",x"5e",x"0e"),
  1171 => (x"4a",x"66",x"cc",x"0e"),
  1172 => (x"ff",x"c3",x"2a",x"d8"),
  1173 => (x"4b",x"66",x"cc",x"9a"),
  1174 => (x"fc",x"cf",x"2b",x"c8"),
  1175 => (x"4a",x"72",x"9b",x"c0"),
  1176 => (x"66",x"cc",x"b2",x"73"),
  1177 => (x"c0",x"33",x"c8",x"4b"),
  1178 => (x"c0",x"c0",x"f0",x"ff"),
  1179 => (x"73",x"4a",x"72",x"9b"),
  1180 => (x"4b",x"66",x"cc",x"b2"),
  1181 => (x"c0",x"ff",x"33",x"d8"),
  1182 => (x"9b",x"c0",x"c0",x"c0"),
  1183 => (x"b2",x"73",x"4a",x"72"),
  1184 => (x"4b",x"26",x"48",x"72"),
  1185 => (x"4f",x"26",x"4a",x"26"),
  1186 => (x"5b",x"5a",x"5e",x"0e"),
  1187 => (x"4b",x"66",x"cc",x"0e"),
  1188 => (x"ff",x"c3",x"2b",x"c8"),
  1189 => (x"66",x"cc",x"4b",x"9b"),
  1190 => (x"cf",x"32",x"c8",x"4a"),
  1191 => (x"72",x"9a",x"c0",x"fc"),
  1192 => (x"4a",x"b2",x"73",x"4a"),
  1193 => (x"4b",x"26",x"48",x"72"),
  1194 => (x"4f",x"26",x"4a",x"26"),
  1195 => (x"5b",x"5a",x"5e",x"0e"),
  1196 => (x"4a",x"66",x"cc",x"0e"),
  1197 => (x"ff",x"cf",x"2a",x"d0"),
  1198 => (x"cc",x"4a",x"9a",x"ff"),
  1199 => (x"33",x"d0",x"4b",x"66"),
  1200 => (x"9b",x"c0",x"c0",x"f0"),
  1201 => (x"b2",x"73",x"4a",x"72"),
  1202 => (x"4b",x"26",x"48",x"72"),
  1203 => (x"4f",x"26",x"4a",x"26"),
  1204 => (x"d0",x"1e",x"72",x"1e"),
  1205 => (x"c0",x"c0",x"c0",x"c0"),
  1206 => (x"ff",x"0f",x"72",x"4a"),
  1207 => (x"4a",x"26",x"87",x"fd"),
  1208 => (x"72",x"1e",x"4f",x"26"),
  1209 => (x"4a",x"66",x"cc",x"1e"),
  1210 => (x"c0",x"9a",x"df",x"c3"),
  1211 => (x"b7",x"c0",x"8a",x"f7"),
  1212 => (x"c3",x"c0",x"03",x"aa"),
  1213 => (x"82",x"e7",x"c0",x"87"),
  1214 => (x"c4",x"48",x"66",x"c8"),
  1215 => (x"58",x"a6",x"cc",x"30"),
  1216 => (x"72",x"48",x"66",x"c8"),
  1217 => (x"58",x"a6",x"cc",x"b0"),
  1218 => (x"26",x"48",x"66",x"c8"),
  1219 => (x"0e",x"4f",x"26",x"4a"),
  1220 => (x"5c",x"5b",x"5a",x"5e"),
  1221 => (x"c0",x"d0",x"0e",x"5d"),
  1222 => (x"4d",x"c0",x"c0",x"c0"),
  1223 => (x"00",x"1b",x"54",x"27"),
  1224 => (x"c1",x"48",x"bf",x"00"),
  1225 => (x"1b",x"58",x"27",x"80"),
  1226 => (x"97",x"58",x"00",x"00"),
  1227 => (x"c1",x"4a",x"66",x"d4"),
  1228 => (x"c0",x"c0",x"c0",x"c0"),
  1229 => (x"b7",x"c0",x"c4",x"92"),
  1230 => (x"d3",x"c1",x"4a",x"92"),
  1231 => (x"c0",x"05",x"aa",x"b7"),
  1232 => (x"54",x"27",x"87",x"e9"),
  1233 => (x"49",x"00",x"00",x"1b"),
  1234 => (x"58",x"27",x"79",x"c0"),
  1235 => (x"49",x"00",x"00",x"1b"),
  1236 => (x"60",x"27",x"79",x"c0"),
  1237 => (x"49",x"00",x"00",x"1b"),
  1238 => (x"64",x"27",x"79",x"c0"),
  1239 => (x"49",x"00",x"00",x"1b"),
  1240 => (x"c0",x"ff",x"79",x"c0"),
  1241 => (x"79",x"d3",x"c1",x"49"),
  1242 => (x"27",x"87",x"cb",x"ca"),
  1243 => (x"00",x"00",x"1b",x"54"),
  1244 => (x"b7",x"c1",x"49",x"bf"),
  1245 => (x"db",x"c1",x"05",x"a9"),
  1246 => (x"49",x"c0",x"ff",x"87"),
  1247 => (x"97",x"79",x"f4",x"c1"),
  1248 => (x"c1",x"4a",x"66",x"d4"),
  1249 => (x"c0",x"c0",x"c0",x"c0"),
  1250 => (x"b7",x"c0",x"c4",x"92"),
  1251 => (x"1e",x"72",x"4a",x"92"),
  1252 => (x"00",x"1b",x"64",x"27"),
  1253 => (x"27",x"1e",x"bf",x"00"),
  1254 => (x"00",x"00",x"12",x"e2"),
  1255 => (x"27",x"86",x"c8",x"0f"),
  1256 => (x"00",x"00",x"1b",x"68"),
  1257 => (x"1b",x"64",x"27",x"58"),
  1258 => (x"4c",x"bf",x"00",x"00"),
  1259 => (x"06",x"ac",x"b7",x"c3"),
  1260 => (x"ca",x"87",x"c6",x"c0"),
  1261 => (x"70",x"88",x"74",x"48"),
  1262 => (x"c1",x"4a",x"74",x"4c"),
  1263 => (x"c1",x"48",x"72",x"82"),
  1264 => (x"1b",x"60",x"27",x"30"),
  1265 => (x"74",x"58",x"00",x"00"),
  1266 => (x"80",x"f0",x"c0",x"48"),
  1267 => (x"70",x"49",x"c0",x"ff"),
  1268 => (x"87",x"e2",x"c8",x"79"),
  1269 => (x"00",x"1b",x"64",x"27"),
  1270 => (x"c9",x"49",x"bf",x"00"),
  1271 => (x"c8",x"01",x"a9",x"b7"),
  1272 => (x"64",x"27",x"87",x"d4"),
  1273 => (x"bf",x"00",x"00",x"1b"),
  1274 => (x"a9",x"b7",x"c0",x"49"),
  1275 => (x"87",x"c6",x"c8",x"06"),
  1276 => (x"00",x"1b",x"64",x"27"),
  1277 => (x"c0",x"48",x"bf",x"00"),
  1278 => (x"c0",x"ff",x"80",x"f0"),
  1279 => (x"27",x"79",x"70",x"49"),
  1280 => (x"00",x"00",x"1b",x"54"),
  1281 => (x"b7",x"c3",x"49",x"bf"),
  1282 => (x"e9",x"c0",x"01",x"a9"),
  1283 => (x"66",x"d4",x"97",x"87"),
  1284 => (x"c0",x"c0",x"c1",x"4a"),
  1285 => (x"c4",x"92",x"c0",x"c0"),
  1286 => (x"4a",x"92",x"b7",x"c0"),
  1287 => (x"60",x"27",x"1e",x"72"),
  1288 => (x"bf",x"00",x"00",x"1b"),
  1289 => (x"12",x"e2",x"27",x"1e"),
  1290 => (x"c8",x"0f",x"00",x"00"),
  1291 => (x"1b",x"64",x"27",x"86"),
  1292 => (x"c7",x"58",x"00",x"00"),
  1293 => (x"5c",x"27",x"87",x"c0"),
  1294 => (x"bf",x"00",x"00",x"1b"),
  1295 => (x"27",x"82",x"c3",x"4a"),
  1296 => (x"00",x"00",x"1b",x"54"),
  1297 => (x"b7",x"72",x"49",x"bf"),
  1298 => (x"f1",x"c0",x"01",x"a9"),
  1299 => (x"66",x"d4",x"97",x"87"),
  1300 => (x"c0",x"c0",x"c1",x"4a"),
  1301 => (x"c4",x"92",x"c0",x"c0"),
  1302 => (x"4a",x"92",x"b7",x"c0"),
  1303 => (x"58",x"27",x"1e",x"72"),
  1304 => (x"bf",x"00",x"00",x"1b"),
  1305 => (x"12",x"e2",x"27",x"1e"),
  1306 => (x"c8",x"0f",x"00",x"00"),
  1307 => (x"1b",x"5c",x"27",x"86"),
  1308 => (x"27",x"58",x"00",x"00"),
  1309 => (x"00",x"00",x"1b",x"68"),
  1310 => (x"c5",x"79",x"c1",x"49"),
  1311 => (x"64",x"27",x"87",x"f8"),
  1312 => (x"bf",x"00",x"00",x"1b"),
  1313 => (x"a9",x"b7",x"c0",x"49"),
  1314 => (x"87",x"d0",x"c3",x"06"),
  1315 => (x"00",x"1b",x"64",x"27"),
  1316 => (x"c3",x"49",x"bf",x"00"),
  1317 => (x"c3",x"01",x"a9",x"b7"),
  1318 => (x"60",x"27",x"87",x"c2"),
  1319 => (x"bf",x"00",x"00",x"1b"),
  1320 => (x"c1",x"32",x"c1",x"4a"),
  1321 => (x"1b",x"54",x"27",x"82"),
  1322 => (x"49",x"bf",x"00",x"00"),
  1323 => (x"01",x"a9",x"b7",x"72"),
  1324 => (x"97",x"87",x"c2",x"c2"),
  1325 => (x"c1",x"4a",x"66",x"d4"),
  1326 => (x"c0",x"c0",x"c0",x"c0"),
  1327 => (x"b7",x"c0",x"c4",x"92"),
  1328 => (x"1e",x"72",x"4a",x"92"),
  1329 => (x"00",x"1b",x"6c",x"27"),
  1330 => (x"27",x"1e",x"bf",x"00"),
  1331 => (x"00",x"00",x"12",x"e2"),
  1332 => (x"27",x"86",x"c8",x"0f"),
  1333 => (x"00",x"00",x"1b",x"70"),
  1334 => (x"1b",x"68",x"27",x"58"),
  1335 => (x"4a",x"bf",x"00",x"00"),
  1336 => (x"68",x"27",x"8a",x"c1"),
  1337 => (x"49",x"00",x"00",x"1b"),
  1338 => (x"b7",x"c0",x"79",x"72"),
  1339 => (x"c5",x"c4",x"03",x"aa"),
  1340 => (x"1b",x"58",x"27",x"87"),
  1341 => (x"4a",x"bf",x"00",x"00"),
  1342 => (x"00",x"1b",x"6c",x"27"),
  1343 => (x"52",x"bf",x"97",x"00"),
  1344 => (x"00",x"1b",x"58",x"27"),
  1345 => (x"c1",x"4a",x"bf",x"00"),
  1346 => (x"1b",x"58",x"27",x"82"),
  1347 => (x"72",x"49",x"00",x"00"),
  1348 => (x"1b",x"70",x"27",x"79"),
  1349 => (x"b7",x"bf",x"00",x"00"),
  1350 => (x"cd",x"c0",x"06",x"aa"),
  1351 => (x"1b",x"70",x"27",x"87"),
  1352 => (x"27",x"49",x"00",x"00"),
  1353 => (x"00",x"00",x"1b",x"58"),
  1354 => (x"68",x"27",x"79",x"bf"),
  1355 => (x"49",x"00",x"00",x"1b"),
  1356 => (x"c1",x"c3",x"79",x"c1"),
  1357 => (x"1b",x"68",x"27",x"87"),
  1358 => (x"05",x"bf",x"00",x"00"),
  1359 => (x"27",x"87",x"f7",x"c2"),
  1360 => (x"00",x"00",x"1b",x"6c"),
  1361 => (x"33",x"c4",x"4b",x"bf"),
  1362 => (x"00",x"1b",x"6c",x"27"),
  1363 => (x"79",x"73",x"49",x"00"),
  1364 => (x"00",x"1b",x"58",x"27"),
  1365 => (x"73",x"4a",x"bf",x"00"),
  1366 => (x"87",x"da",x"c2",x"52"),
  1367 => (x"00",x"1b",x"64",x"27"),
  1368 => (x"c7",x"49",x"bf",x"00"),
  1369 => (x"c1",x"04",x"a9",x"b7"),
  1370 => (x"4b",x"c0",x"87",x"fd"),
  1371 => (x"c1",x"49",x"f4",x"fe"),
  1372 => (x"1b",x"70",x"27",x"79"),
  1373 => (x"1e",x"bf",x"00",x"00"),
  1374 => (x"c0",x"27",x"1e",x"75"),
  1375 => (x"1e",x"00",x"00",x"18"),
  1376 => (x"00",x"00",x"97",x"27"),
  1377 => (x"86",x"cc",x"0f",x"00"),
  1378 => (x"00",x"1b",x"58",x"27"),
  1379 => (x"79",x"75",x"49",x"00"),
  1380 => (x"00",x"1b",x"58",x"27"),
  1381 => (x"27",x"49",x"bf",x"00"),
  1382 => (x"00",x"00",x"1b",x"70"),
  1383 => (x"03",x"a9",x"b7",x"bf"),
  1384 => (x"27",x"87",x"e5",x"c0"),
  1385 => (x"00",x"00",x"1b",x"58"),
  1386 => (x"27",x"83",x"bf",x"bf"),
  1387 => (x"00",x"00",x"1b",x"58"),
  1388 => (x"82",x"c4",x"4a",x"bf"),
  1389 => (x"00",x"1b",x"58",x"27"),
  1390 => (x"79",x"72",x"49",x"00"),
  1391 => (x"00",x"1b",x"70",x"27"),
  1392 => (x"aa",x"b7",x"bf",x"00"),
  1393 => (x"87",x"db",x"ff",x"04"),
  1394 => (x"df",x"27",x"1e",x"73"),
  1395 => (x"1e",x"00",x"00",x"18"),
  1396 => (x"00",x"00",x"97",x"27"),
  1397 => (x"86",x"c8",x"0f",x"00"),
  1398 => (x"c1",x"49",x"c0",x"ff"),
  1399 => (x"d0",x"27",x"79",x"c2"),
  1400 => (x"0f",x"00",x"00",x"12"),
  1401 => (x"27",x"87",x"cf",x"c0"),
  1402 => (x"00",x"00",x"1b",x"64"),
  1403 => (x"f0",x"c0",x"48",x"bf"),
  1404 => (x"49",x"c0",x"ff",x"80"),
  1405 => (x"4d",x"26",x"79",x"70"),
  1406 => (x"4b",x"26",x"4c",x"26"),
  1407 => (x"4f",x"26",x"4a",x"26"),
  1408 => (x"5b",x"5a",x"5e",x"0e"),
  1409 => (x"1e",x"0e",x"5d",x"5c"),
  1410 => (x"00",x"17",x"13",x"27"),
  1411 => (x"61",x"27",x"1e",x"00"),
  1412 => (x"0f",x"00",x"00",x"00"),
  1413 => (x"fc",x"27",x"86",x"c4"),
  1414 => (x"0f",x"00",x"00",x"04"),
  1415 => (x"9a",x"72",x"4a",x"70"),
  1416 => (x"87",x"d3",x"c0",x"02"),
  1417 => (x"00",x"0a",x"bd",x"27"),
  1418 => (x"4a",x"70",x"0f",x"00"),
  1419 => (x"c0",x"02",x"9a",x"72"),
  1420 => (x"4a",x"c1",x"87",x"c5"),
  1421 => (x"c0",x"87",x"c2",x"c0"),
  1422 => (x"72",x"49",x"76",x"4a"),
  1423 => (x"17",x"29",x"27",x"79"),
  1424 => (x"27",x"1e",x"00",x"00"),
  1425 => (x"00",x"00",x"00",x"61"),
  1426 => (x"27",x"86",x"c4",x"0f"),
  1427 => (x"00",x"00",x"1b",x"70"),
  1428 => (x"c0",x"79",x"c0",x"49"),
  1429 => (x"42",x"27",x"1e",x"ee"),
  1430 => (x"0f",x"00",x"00",x"00"),
  1431 => (x"f4",x"c3",x"86",x"c4"),
  1432 => (x"ff",x"4b",x"ff",x"c8"),
  1433 => (x"74",x"4c",x"bf",x"c0"),
  1434 => (x"9a",x"c0",x"c8",x"4a"),
  1435 => (x"c1",x"02",x"9a",x"72"),
  1436 => (x"4d",x"74",x"87",x"e1"),
  1437 => (x"db",x"9d",x"ff",x"c3"),
  1438 => (x"c1",x"05",x"ad",x"b7"),
  1439 => (x"02",x"6e",x"87",x"c6"),
  1440 => (x"d0",x"87",x"f3",x"c0"),
  1441 => (x"c0",x"c0",x"c0",x"c0"),
  1442 => (x"16",x"f7",x"27",x"1e"),
  1443 => (x"27",x"1e",x"00",x"00"),
  1444 => (x"00",x"00",x"11",x"7c"),
  1445 => (x"70",x"86",x"c8",x"0f"),
  1446 => (x"02",x"9a",x"72",x"4a"),
  1447 => (x"27",x"87",x"d7",x"c0"),
  1448 => (x"00",x"00",x"16",x"eb"),
  1449 => (x"00",x"61",x"27",x"1e"),
  1450 => (x"c4",x"0f",x"00",x"00"),
  1451 => (x"12",x"d0",x"27",x"86"),
  1452 => (x"c0",x"0f",x"00",x"00"),
  1453 => (x"03",x"27",x"87",x"ce"),
  1454 => (x"1e",x"00",x"00",x"17"),
  1455 => (x"00",x"00",x"61",x"27"),
  1456 => (x"86",x"c4",x"0f",x"00"),
  1457 => (x"0f",x"27",x"1e",x"75"),
  1458 => (x"0f",x"00",x"00",x"13"),
  1459 => (x"f4",x"c3",x"86",x"c4"),
  1460 => (x"73",x"4b",x"c0",x"c9"),
  1461 => (x"72",x"8b",x"c1",x"4a"),
  1462 => (x"c6",x"fe",x"05",x"9a"),
  1463 => (x"87",x"f3",x"fd",x"87"),
  1464 => (x"26",x"4d",x"26",x"26"),
  1465 => (x"26",x"4b",x"26",x"4c"),
  1466 => (x"42",x"4f",x"26",x"4a"),
  1467 => (x"69",x"74",x"6f",x"6f"),
  1468 => (x"2e",x"2e",x"67",x"6e"),
  1469 => (x"42",x"00",x"0a",x"2e"),
  1470 => (x"38",x"54",x"4f",x"4f"),
  1471 => (x"42",x"20",x"32",x"33"),
  1472 => (x"53",x"00",x"4e",x"49"),
  1473 => (x"6f",x"62",x"20",x"44"),
  1474 => (x"66",x"20",x"74",x"6f"),
  1475 => (x"65",x"6c",x"69",x"61"),
  1476 => (x"49",x"00",x"0a",x"64"),
  1477 => (x"69",x"74",x"69",x"6e"),
  1478 => (x"7a",x"69",x"6c",x"61"),
  1479 => (x"20",x"67",x"6e",x"69"),
  1480 => (x"63",x"20",x"44",x"53"),
  1481 => (x"0a",x"64",x"72",x"61"),
  1482 => (x"32",x"53",x"52",x"00"),
  1483 => (x"62",x"20",x"32",x"33"),
  1484 => (x"20",x"74",x"6f",x"6f"),
  1485 => (x"72",x"70",x"20",x"2d"),
  1486 => (x"20",x"73",x"73",x"65"),
  1487 => (x"20",x"43",x"53",x"45"),
  1488 => (x"62",x"20",x"6f",x"74"),
  1489 => (x"20",x"74",x"6f",x"6f"),
  1490 => (x"6d",x"6f",x"72",x"66"),
  1491 => (x"2e",x"44",x"53",x"20"),
  1492 => (x"44",x"4d",x"43",x"00"),
  1493 => (x"61",x"65",x"52",x"00"),
  1494 => (x"66",x"6f",x"20",x"64"),
  1495 => (x"52",x"42",x"4d",x"20"),
  1496 => (x"69",x"61",x"66",x"20"),
  1497 => (x"0a",x"64",x"65",x"6c"),
  1498 => (x"20",x"6f",x"4e",x"00"),
  1499 => (x"74",x"72",x"61",x"70"),
  1500 => (x"6f",x"69",x"74",x"69"),
  1501 => (x"69",x"73",x"20",x"6e"),
  1502 => (x"74",x"61",x"6e",x"67"),
  1503 => (x"20",x"65",x"72",x"75"),
  1504 => (x"6e",x"75",x"6f",x"66"),
  1505 => (x"4d",x"00",x"0a",x"64"),
  1506 => (x"69",x"73",x"52",x"42"),
  1507 => (x"20",x"3a",x"65",x"7a"),
  1508 => (x"20",x"2c",x"64",x"25"),
  1509 => (x"74",x"72",x"61",x"70"),
  1510 => (x"6f",x"69",x"74",x"69"),
  1511 => (x"7a",x"69",x"73",x"6e"),
  1512 => (x"25",x"20",x"3a",x"65"),
  1513 => (x"6f",x"20",x"2c",x"64"),
  1514 => (x"65",x"73",x"66",x"66"),
  1515 => (x"66",x"6f",x"20",x"74"),
  1516 => (x"67",x"69",x"73",x"20"),
  1517 => (x"64",x"25",x"20",x"3a"),
  1518 => (x"69",x"73",x"20",x"2c"),
  1519 => (x"78",x"30",x"20",x"67"),
  1520 => (x"00",x"0a",x"78",x"25"),
  1521 => (x"64",x"61",x"65",x"52"),
  1522 => (x"20",x"67",x"6e",x"69"),
  1523 => (x"74",x"6f",x"6f",x"62"),
  1524 => (x"63",x"65",x"73",x"20"),
  1525 => (x"20",x"72",x"6f",x"74"),
  1526 => (x"00",x"0a",x"64",x"25"),
  1527 => (x"64",x"61",x"65",x"52"),
  1528 => (x"6f",x"6f",x"62",x"20"),
  1529 => (x"65",x"73",x"20",x"74"),
  1530 => (x"72",x"6f",x"74",x"63"),
  1531 => (x"6f",x"72",x"66",x"20"),
  1532 => (x"69",x"66",x"20",x"6d"),
  1533 => (x"20",x"74",x"73",x"72"),
  1534 => (x"74",x"72",x"61",x"70"),
  1535 => (x"6f",x"69",x"74",x"69"),
  1536 => (x"55",x"00",x"0a",x"6e"),
  1537 => (x"70",x"75",x"73",x"6e"),
  1538 => (x"74",x"72",x"6f",x"70"),
  1539 => (x"70",x"20",x"64",x"65"),
  1540 => (x"69",x"74",x"72",x"61"),
  1541 => (x"6e",x"6f",x"69",x"74"),
  1542 => (x"70",x"79",x"74",x"20"),
  1543 => (x"00",x"0d",x"21",x"65"),
  1544 => (x"33",x"54",x"41",x"46"),
  1545 => (x"20",x"20",x"20",x"32"),
  1546 => (x"61",x"65",x"52",x"00"),
  1547 => (x"67",x"6e",x"69",x"64"),
  1548 => (x"52",x"42",x"4d",x"20"),
  1549 => (x"42",x"4d",x"00",x"0a"),
  1550 => (x"75",x"73",x"20",x"52"),
  1551 => (x"73",x"65",x"63",x"63"),
  1552 => (x"6c",x"75",x"66",x"73"),
  1553 => (x"72",x"20",x"79",x"6c"),
  1554 => (x"0a",x"64",x"61",x"65"),
  1555 => (x"54",x"41",x"46",x"00"),
  1556 => (x"20",x"20",x"36",x"31"),
  1557 => (x"41",x"46",x"00",x"20"),
  1558 => (x"20",x"32",x"33",x"54"),
  1559 => (x"50",x"00",x"20",x"20"),
  1560 => (x"69",x"74",x"72",x"61"),
  1561 => (x"6e",x"6f",x"69",x"74"),
  1562 => (x"6e",x"75",x"6f",x"63"),
  1563 => (x"64",x"25",x"20",x"74"),
  1564 => (x"75",x"48",x"00",x"0a"),
  1565 => (x"6e",x"69",x"74",x"6e"),
  1566 => (x"6f",x"66",x"20",x"67"),
  1567 => (x"69",x"66",x"20",x"72"),
  1568 => (x"79",x"73",x"65",x"6c"),
  1569 => (x"6d",x"65",x"74",x"73"),
  1570 => (x"41",x"46",x"00",x"0a"),
  1571 => (x"20",x"32",x"33",x"54"),
  1572 => (x"46",x"00",x"20",x"20"),
  1573 => (x"36",x"31",x"54",x"41"),
  1574 => (x"00",x"20",x"20",x"20"),
  1575 => (x"73",x"75",x"6c",x"43"),
  1576 => (x"20",x"72",x"65",x"74"),
  1577 => (x"65",x"7a",x"69",x"73"),
  1578 => (x"64",x"25",x"20",x"3a"),
  1579 => (x"6c",x"43",x"20",x"2c"),
  1580 => (x"65",x"74",x"73",x"75"),
  1581 => (x"61",x"6d",x"20",x"72"),
  1582 => (x"20",x"2c",x"6b",x"73"),
  1583 => (x"00",x"0a",x"64",x"25"),
  1584 => (x"63",x"65",x"68",x"43"),
  1585 => (x"6d",x"75",x"73",x"6b"),
  1586 => (x"67",x"6e",x"69",x"6d"),
  1587 => (x"6f",x"72",x"66",x"20"),
  1588 => (x"64",x"25",x"20",x"6d"),
  1589 => (x"20",x"6f",x"74",x"20"),
  1590 => (x"2e",x"2e",x"64",x"25"),
  1591 => (x"25",x"00",x"20",x"2e"),
  1592 => (x"25",x"00",x"0a",x"64"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
