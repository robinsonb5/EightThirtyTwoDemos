
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"2c",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"29"),
    10 => (x"87",x"fd",x"00",x"4f"),
    11 => (x"f8",x"f1",x"c3",x"4f"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"f8",x"f1",x"c3"),
    14 => (x"48",x"c0",x"cf",x"c1"),
    15 => (x"03",x"89",x"d0",x"89"),
    16 => (x"40",x"40",x"40",x"c0"),
    17 => (x"d0",x"87",x"f6",x"40"),
    18 => (x"50",x"c0",x"05",x"81"),
    19 => (x"f9",x"05",x"89",x"c1"),
    20 => (x"c0",x"cf",x"c1",x"87"),
    21 => (x"c0",x"cf",x"c1",x"4d"),
    22 => (x"02",x"ad",x"74",x"4c"),
    23 => (x"0f",x"24",x"87",x"c4"),
    24 => (x"e3",x"cd",x"87",x"f7"),
    25 => (x"c0",x"cf",x"c1",x"87"),
    26 => (x"c0",x"cf",x"c1",x"4d"),
    27 => (x"02",x"ad",x"74",x"4c"),
    28 => (x"8c",x"c4",x"87",x"c6"),
    29 => (x"87",x"f5",x"0f",x"6c"),
    30 => (x"0e",x"87",x"fd",x"00"),
    31 => (x"5d",x"5c",x"5b",x"5e"),
    32 => (x"71",x"86",x"fc",x"0e"),
    33 => (x"66",x"e0",x"c0",x"4a"),
    34 => (x"c0",x"cf",x"c1",x"4c"),
    35 => (x"72",x"7e",x"c0",x"4b"),
    36 => (x"87",x"ce",x"05",x"9a"),
    37 => (x"4b",x"c1",x"cf",x"c1"),
    38 => (x"48",x"c0",x"cf",x"c1"),
    39 => (x"c1",x"50",x"f0",x"c0"),
    40 => (x"9a",x"72",x"87",x"cd"),
    41 => (x"87",x"e4",x"c0",x"02"),
    42 => (x"72",x"4d",x"66",x"d4"),
    43 => (x"75",x"49",x"72",x"1e"),
    44 => (x"87",x"ef",x"ca",x"4a"),
    45 => (x"e0",x"c4",x"4a",x"26"),
    46 => (x"72",x"53",x"11",x"81"),
    47 => (x"ca",x"4a",x"75",x"49"),
    48 => (x"4a",x"70",x"87",x"e1"),
    49 => (x"9a",x"72",x"8c",x"c1"),
    50 => (x"87",x"df",x"ff",x"05"),
    51 => (x"06",x"ac",x"b7",x"c0"),
    52 => (x"e4",x"c0",x"87",x"dd"),
    53 => (x"87",x"c5",x"02",x"66"),
    54 => (x"c3",x"4a",x"f0",x"c0"),
    55 => (x"4a",x"e0",x"c0",x"87"),
    56 => (x"7a",x"97",x"0a",x"73"),
    57 => (x"8c",x"83",x"c1",x"0a"),
    58 => (x"01",x"ac",x"b7",x"c0"),
    59 => (x"c1",x"87",x"e3",x"ff"),
    60 => (x"02",x"ab",x"c0",x"cf"),
    61 => (x"66",x"d8",x"87",x"de"),
    62 => (x"1e",x"66",x"dc",x"4c"),
    63 => (x"6b",x"97",x"8b",x"c1"),
    64 => (x"c4",x"0f",x"74",x"49"),
    65 => (x"c1",x"48",x"6e",x"86"),
    66 => (x"58",x"a6",x"c4",x"80"),
    67 => (x"ab",x"c0",x"cf",x"c1"),
    68 => (x"87",x"e5",x"ff",x"05"),
    69 => (x"8e",x"fc",x"48",x"6e"),
    70 => (x"4c",x"26",x"4d",x"26"),
    71 => (x"4f",x"26",x"4b",x"26"),
    72 => (x"33",x"32",x"31",x"30"),
    73 => (x"37",x"36",x"35",x"34"),
    74 => (x"42",x"41",x"39",x"38"),
    75 => (x"46",x"45",x"44",x"43"),
    76 => (x"5b",x"5e",x"0e",x"00"),
    77 => (x"71",x"0e",x"5d",x"5c"),
    78 => (x"13",x"4d",x"ff",x"4b"),
    79 => (x"d7",x"02",x"9c",x"4c"),
    80 => (x"d4",x"85",x"c1",x"87"),
    81 => (x"49",x"74",x"1e",x"66"),
    82 => (x"c4",x"0f",x"66",x"d4"),
    83 => (x"05",x"a8",x"74",x"86"),
    84 => (x"4c",x"13",x"87",x"c6"),
    85 => (x"87",x"e9",x"05",x"9c"),
    86 => (x"4d",x"26",x"48",x"75"),
    87 => (x"4b",x"26",x"4c",x"26"),
    88 => (x"5e",x"0e",x"4f",x"26"),
    89 => (x"0e",x"5d",x"5c",x"5b"),
    90 => (x"a6",x"c4",x"86",x"e8"),
    91 => (x"66",x"e8",x"c0",x"59"),
    92 => (x"c8",x"4c",x"c0",x"4d"),
    93 => (x"78",x"c0",x"48",x"a6"),
    94 => (x"4b",x"bf",x"97",x"6e"),
    95 => (x"80",x"c1",x"48",x"6e"),
    96 => (x"73",x"58",x"a6",x"c4"),
    97 => (x"ce",x"c6",x"02",x"9b"),
    98 => (x"02",x"66",x"c8",x"87"),
    99 => (x"cc",x"87",x"d6",x"c5"),
   100 => (x"78",x"c0",x"48",x"a6"),
   101 => (x"78",x"c0",x"80",x"fc"),
   102 => (x"e0",x"c0",x"4a",x"73"),
   103 => (x"c2",x"c3",x"02",x"8a"),
   104 => (x"02",x"8a",x"c3",x"87"),
   105 => (x"c2",x"87",x"fc",x"c2"),
   106 => (x"e4",x"c2",x"02",x"8a"),
   107 => (x"c2",x"02",x"8a",x"87"),
   108 => (x"8a",x"c4",x"87",x"f1"),
   109 => (x"87",x"eb",x"c2",x"02"),
   110 => (x"c2",x"02",x"8a",x"c2"),
   111 => (x"8a",x"c3",x"87",x"e5"),
   112 => (x"87",x"e7",x"c2",x"02"),
   113 => (x"c0",x"02",x"8a",x"d4"),
   114 => (x"02",x"8a",x"87",x"f4"),
   115 => (x"ca",x"87",x"ff",x"c0"),
   116 => (x"f1",x"c0",x"02",x"8a"),
   117 => (x"02",x"8a",x"c1",x"87"),
   118 => (x"8a",x"87",x"df",x"c1"),
   119 => (x"c8",x"87",x"df",x"02"),
   120 => (x"cd",x"c1",x"02",x"8a"),
   121 => (x"02",x"8a",x"c4",x"87"),
   122 => (x"c3",x"87",x"e3",x"c0"),
   123 => (x"e5",x"c0",x"02",x"8a"),
   124 => (x"02",x"8a",x"c2",x"87"),
   125 => (x"8a",x"c3",x"87",x"c8"),
   126 => (x"c1",x"87",x"d3",x"02"),
   127 => (x"a6",x"cc",x"87",x"f9"),
   128 => (x"c2",x"78",x"ca",x"48"),
   129 => (x"a6",x"cc",x"87",x"d1"),
   130 => (x"c2",x"78",x"c2",x"48"),
   131 => (x"a6",x"cc",x"87",x"c9"),
   132 => (x"c2",x"78",x"d0",x"48"),
   133 => (x"f0",x"c0",x"87",x"c1"),
   134 => (x"f0",x"c0",x"1e",x"66"),
   135 => (x"85",x"c4",x"1e",x"66"),
   136 => (x"8a",x"c4",x"4a",x"75"),
   137 => (x"c8",x"fc",x"49",x"6a"),
   138 => (x"70",x"86",x"c8",x"87"),
   139 => (x"c1",x"4c",x"a4",x"49"),
   140 => (x"a6",x"c8",x"87",x"e5"),
   141 => (x"c1",x"78",x"c1",x"48"),
   142 => (x"f0",x"c0",x"87",x"dd"),
   143 => (x"85",x"c4",x"1e",x"66"),
   144 => (x"8a",x"c4",x"4a",x"75"),
   145 => (x"f0",x"c0",x"49",x"6a"),
   146 => (x"86",x"c4",x"0f",x"66"),
   147 => (x"c6",x"c1",x"84",x"c1"),
   148 => (x"66",x"f0",x"c0",x"87"),
   149 => (x"49",x"e5",x"c0",x"1e"),
   150 => (x"0f",x"66",x"f0",x"c0"),
   151 => (x"84",x"c1",x"86",x"c4"),
   152 => (x"c8",x"87",x"f4",x"c0"),
   153 => (x"78",x"c1",x"48",x"a6"),
   154 => (x"d0",x"87",x"ec",x"c0"),
   155 => (x"78",x"c1",x"48",x"a6"),
   156 => (x"78",x"c1",x"80",x"f8"),
   157 => (x"c0",x"87",x"e0",x"c0"),
   158 => (x"da",x"06",x"ab",x"f0"),
   159 => (x"ab",x"f9",x"c0",x"87"),
   160 => (x"d4",x"87",x"d4",x"03"),
   161 => (x"91",x"ca",x"49",x"66"),
   162 => (x"f0",x"c0",x"4a",x"73"),
   163 => (x"48",x"a6",x"d4",x"8a"),
   164 => (x"f4",x"78",x"a1",x"72"),
   165 => (x"cc",x"78",x"c1",x"80"),
   166 => (x"e9",x"c1",x"02",x"66"),
   167 => (x"75",x"85",x"c4",x"87"),
   168 => (x"a6",x"89",x"c4",x"49"),
   169 => (x"c1",x"78",x"69",x"48"),
   170 => (x"d8",x"05",x"ab",x"e4"),
   171 => (x"48",x"66",x"c4",x"87"),
   172 => (x"03",x"a8",x"b7",x"c0"),
   173 => (x"ed",x"c0",x"87",x"cf"),
   174 => (x"87",x"fa",x"c1",x"49"),
   175 => (x"c0",x"48",x"66",x"c4"),
   176 => (x"a6",x"c8",x"88",x"08"),
   177 => (x"1e",x"66",x"d0",x"58"),
   178 => (x"c0",x"1e",x"66",x"d8"),
   179 => (x"c0",x"1e",x"66",x"f8"),
   180 => (x"dc",x"1e",x"66",x"f8"),
   181 => (x"66",x"d8",x"1e",x"66"),
   182 => (x"87",x"df",x"f6",x"49"),
   183 => (x"49",x"70",x"86",x"d4"),
   184 => (x"e1",x"c0",x"4c",x"a4"),
   185 => (x"ab",x"e5",x"c0",x"87"),
   186 => (x"d0",x"87",x"cf",x"05"),
   187 => (x"78",x"c0",x"48",x"a6"),
   188 => (x"78",x"c0",x"80",x"c4"),
   189 => (x"78",x"c1",x"80",x"f4"),
   190 => (x"f0",x"c0",x"87",x"cc"),
   191 => (x"49",x"73",x"1e",x"66"),
   192 => (x"0f",x"66",x"f0",x"c0"),
   193 => (x"97",x"6e",x"86",x"c4"),
   194 => (x"48",x"6e",x"4b",x"bf"),
   195 => (x"a6",x"c4",x"80",x"c1"),
   196 => (x"05",x"9b",x"73",x"58"),
   197 => (x"74",x"87",x"f2",x"f9"),
   198 => (x"26",x"8e",x"e8",x"48"),
   199 => (x"26",x"4c",x"26",x"4d"),
   200 => (x"1e",x"4f",x"26",x"4b"),
   201 => (x"f6",x"cc",x"1e",x"c0"),
   202 => (x"1e",x"a6",x"d0",x"1e"),
   203 => (x"f8",x"49",x"66",x"d0"),
   204 => (x"8e",x"f4",x"87",x"f0"),
   205 => (x"fc",x"1e",x"4f",x"26"),
   206 => (x"ff",x"4a",x"71",x"86"),
   207 => (x"48",x"69",x"49",x"c0"),
   208 => (x"c4",x"98",x"c0",x"c4"),
   209 => (x"98",x"70",x"58",x"a6"),
   210 => (x"72",x"87",x"f3",x"02"),
   211 => (x"8e",x"fc",x"48",x"79"),
   212 => (x"72",x"1e",x"4f",x"26"),
   213 => (x"11",x"48",x"12",x"1e"),
   214 => (x"88",x"87",x"c4",x"02"),
   215 => (x"26",x"87",x"f6",x"02"),
   216 => (x"1e",x"4f",x"26",x"4a"),
   217 => (x"9a",x"72",x"1e",x"73"),
   218 => (x"87",x"e7",x"c0",x"02"),
   219 => (x"4b",x"c1",x"48",x"c0"),
   220 => (x"d1",x"06",x"a9",x"72"),
   221 => (x"06",x"82",x"72",x"87"),
   222 => (x"83",x"73",x"87",x"c9"),
   223 => (x"f4",x"01",x"a9",x"72"),
   224 => (x"c1",x"87",x"c3",x"87"),
   225 => (x"a9",x"72",x"3a",x"b2"),
   226 => (x"80",x"73",x"89",x"03"),
   227 => (x"2b",x"2a",x"c1",x"07"),
   228 => (x"26",x"87",x"f3",x"05"),
   229 => (x"1e",x"4f",x"26",x"4b"),
   230 => (x"4d",x"c4",x"1e",x"75"),
   231 => (x"04",x"a1",x"b7",x"71"),
   232 => (x"81",x"c1",x"b9",x"ff"),
   233 => (x"72",x"07",x"bd",x"c3"),
   234 => (x"ff",x"04",x"a2",x"b7"),
   235 => (x"c1",x"82",x"c1",x"ba"),
   236 => (x"ee",x"fe",x"07",x"bd"),
   237 => (x"04",x"2d",x"c1",x"87"),
   238 => (x"80",x"c1",x"b8",x"ff"),
   239 => (x"ff",x"04",x"2d",x"07"),
   240 => (x"07",x"81",x"c1",x"b9"),
   241 => (x"4f",x"26",x"4d",x"26"),
   242 => (x"5c",x"5b",x"5e",x"0e"),
   243 => (x"dc",x"ff",x"0e",x"5d"),
   244 => (x"d4",x"cf",x"c1",x"86"),
   245 => (x"d8",x"ef",x"c3",x"48"),
   246 => (x"d0",x"cf",x"c1",x"78"),
   247 => (x"c8",x"f0",x"c3",x"48"),
   248 => (x"ef",x"c3",x"48",x"78"),
   249 => (x"f0",x"c3",x"78",x"d8"),
   250 => (x"78",x"c0",x"48",x"cc"),
   251 => (x"78",x"c2",x"80",x"c4"),
   252 => (x"e8",x"c0",x"80",x"c4"),
   253 => (x"c0",x"1e",x"71",x"78"),
   254 => (x"c3",x"48",x"c0",x"ee"),
   255 => (x"20",x"49",x"d8",x"f0"),
   256 => (x"20",x"41",x"20",x"41"),
   257 => (x"20",x"41",x"20",x"41"),
   258 => (x"20",x"41",x"20",x"41"),
   259 => (x"10",x"51",x"10",x"41"),
   260 => (x"26",x"51",x"10",x"51"),
   261 => (x"ee",x"c0",x"1e",x"49"),
   262 => (x"f0",x"c3",x"48",x"e0"),
   263 => (x"41",x"20",x"49",x"f8"),
   264 => (x"41",x"20",x"41",x"20"),
   265 => (x"41",x"20",x"41",x"20"),
   266 => (x"41",x"20",x"41",x"20"),
   267 => (x"51",x"10",x"51",x"10"),
   268 => (x"49",x"26",x"51",x"10"),
   269 => (x"48",x"cc",x"ec",x"c1"),
   270 => (x"ef",x"c0",x"78",x"ca"),
   271 => (x"e2",x"fb",x"1e",x"c0"),
   272 => (x"c4",x"ef",x"c0",x"87"),
   273 => (x"87",x"db",x"fb",x"1e"),
   274 => (x"1e",x"f4",x"ef",x"c0"),
   275 => (x"cc",x"87",x"d4",x"fb"),
   276 => (x"e4",x"e7",x"c0",x"86"),
   277 => (x"87",x"d2",x"02",x"bf"),
   278 => (x"1e",x"ec",x"e7",x"c0"),
   279 => (x"c0",x"87",x"c4",x"fb"),
   280 => (x"fa",x"1e",x"d8",x"e8"),
   281 => (x"86",x"c8",x"87",x"fd"),
   282 => (x"e8",x"c0",x"87",x"d0"),
   283 => (x"f2",x"fa",x"1e",x"dc"),
   284 => (x"cc",x"e9",x"c0",x"87"),
   285 => (x"87",x"eb",x"fa",x"1e"),
   286 => (x"e7",x"c0",x"86",x"c8"),
   287 => (x"c0",x"1e",x"bf",x"e8"),
   288 => (x"fa",x"1e",x"f8",x"ef"),
   289 => (x"86",x"c8",x"87",x"dd"),
   290 => (x"48",x"c0",x"ef",x"c3"),
   291 => (x"78",x"bf",x"c8",x"ff"),
   292 => (x"c1",x"48",x"a6",x"c4"),
   293 => (x"e8",x"e7",x"c0",x"78"),
   294 => (x"b7",x"c0",x"48",x"bf"),
   295 => (x"ea",x"c8",x"06",x"a8"),
   296 => (x"48",x"a6",x"c8",x"87"),
   297 => (x"d0",x"58",x"a6",x"d0"),
   298 => (x"a6",x"d8",x"48",x"a6"),
   299 => (x"48",x"a6",x"d8",x"58"),
   300 => (x"c1",x"58",x"a6",x"c4"),
   301 => (x"c1",x"48",x"e0",x"cf"),
   302 => (x"cf",x"c1",x"50",x"c1"),
   303 => (x"78",x"c0",x"48",x"dc"),
   304 => (x"97",x"e0",x"cf",x"c1"),
   305 => (x"c1",x"c1",x"49",x"bf"),
   306 => (x"c8",x"c0",x"02",x"a9"),
   307 => (x"48",x"a6",x"dc",x"87"),
   308 => (x"c5",x"c0",x"78",x"c0"),
   309 => (x"48",x"a6",x"dc",x"87"),
   310 => (x"cf",x"c1",x"78",x"c1"),
   311 => (x"dc",x"48",x"bf",x"dc"),
   312 => (x"cf",x"c1",x"b0",x"66"),
   313 => (x"cf",x"c1",x"58",x"e0"),
   314 => (x"c2",x"c1",x"48",x"e4"),
   315 => (x"48",x"a6",x"d8",x"50"),
   316 => (x"80",x"c8",x"78",x"c2"),
   317 => (x"e9",x"c0",x"78",x"c3"),
   318 => (x"f1",x"c3",x"48",x"f0"),
   319 => (x"41",x"20",x"49",x"d8"),
   320 => (x"41",x"20",x"41",x"20"),
   321 => (x"41",x"20",x"41",x"20"),
   322 => (x"41",x"20",x"41",x"20"),
   323 => (x"51",x"10",x"51",x"10"),
   324 => (x"a6",x"d0",x"51",x"10"),
   325 => (x"c3",x"78",x"c1",x"48"),
   326 => (x"c3",x"1e",x"d8",x"f1"),
   327 => (x"c0",x"49",x"f8",x"f0"),
   328 => (x"c4",x"87",x"e7",x"f8"),
   329 => (x"05",x"98",x"70",x"86"),
   330 => (x"dc",x"87",x"c8",x"c0"),
   331 => (x"78",x"c1",x"48",x"a6"),
   332 => (x"dc",x"87",x"c5",x"c0"),
   333 => (x"78",x"c0",x"48",x"a6"),
   334 => (x"48",x"dc",x"cf",x"c1"),
   335 => (x"d8",x"78",x"66",x"dc"),
   336 => (x"b7",x"c3",x"48",x"66"),
   337 => (x"ea",x"c0",x"03",x"a8"),
   338 => (x"49",x"66",x"d8",x"87"),
   339 => (x"48",x"71",x"91",x"c5"),
   340 => (x"a6",x"cc",x"88",x"c3"),
   341 => (x"1e",x"66",x"cc",x"58"),
   342 => (x"e0",x"c0",x"1e",x"c3"),
   343 => (x"f4",x"c0",x"49",x"66"),
   344 => (x"86",x"c8",x"87",x"f2"),
   345 => (x"c1",x"48",x"66",x"d8"),
   346 => (x"58",x"a6",x"dc",x"80"),
   347 => (x"04",x"a8",x"b7",x"c3"),
   348 => (x"c8",x"87",x"d6",x"ff"),
   349 => (x"66",x"dc",x"1e",x"66"),
   350 => (x"f0",x"d2",x"c1",x"1e"),
   351 => (x"e8",x"cf",x"c1",x"1e"),
   352 => (x"e0",x"f4",x"c0",x"49"),
   353 => (x"c1",x"86",x"cc",x"87"),
   354 => (x"4c",x"bf",x"d0",x"cf"),
   355 => (x"bf",x"d0",x"cf",x"c1"),
   356 => (x"1e",x"72",x"4b",x"bf"),
   357 => (x"bf",x"d0",x"cf",x"c1"),
   358 => (x"c0",x"49",x"73",x"48"),
   359 => (x"20",x"4a",x"a1",x"f0"),
   360 => (x"05",x"aa",x"71",x"41"),
   361 => (x"26",x"87",x"f8",x"ff"),
   362 => (x"49",x"a4",x"cc",x"4a"),
   363 => (x"a3",x"cc",x"79",x"c5"),
   364 => (x"6c",x"7d",x"69",x"4d"),
   365 => (x"cf",x"49",x"73",x"7b"),
   366 => (x"a3",x"c4",x"87",x"ff"),
   367 => (x"c0",x"05",x"69",x"49"),
   368 => (x"a3",x"c8",x"87",x"e5"),
   369 => (x"71",x"7d",x"c6",x"49"),
   370 => (x"4a",x"a4",x"c8",x"1e"),
   371 => (x"f1",x"c0",x"49",x"6a"),
   372 => (x"cf",x"c1",x"87",x"e5"),
   373 => (x"7b",x"bf",x"bf",x"d0"),
   374 => (x"1e",x"ca",x"1e",x"75"),
   375 => (x"f2",x"c0",x"49",x"6d"),
   376 => (x"86",x"cc",x"87",x"f2"),
   377 => (x"6c",x"87",x"d9",x"c0"),
   378 => (x"1e",x"72",x"1e",x"49"),
   379 => (x"49",x"74",x"48",x"71"),
   380 => (x"4a",x"a1",x"f0",x"c0"),
   381 => (x"aa",x"71",x"41",x"20"),
   382 => (x"87",x"f8",x"ff",x"05"),
   383 => (x"49",x"26",x"4a",x"26"),
   384 => (x"c1",x"48",x"a6",x"dc"),
   385 => (x"cf",x"c1",x"50",x"c1"),
   386 => (x"49",x"bf",x"97",x"e4"),
   387 => (x"a9",x"b7",x"c1",x"c1"),
   388 => (x"87",x"db",x"c1",x"04"),
   389 => (x"4b",x"66",x"97",x"dc"),
   390 => (x"73",x"1e",x"c3",x"c1"),
   391 => (x"c7",x"f4",x"c0",x"49"),
   392 => (x"d0",x"86",x"c4",x"87"),
   393 => (x"c0",x"05",x"a8",x"66"),
   394 => (x"66",x"d4",x"87",x"f5"),
   395 => (x"c0",x"49",x"c0",x"1e"),
   396 => (x"c4",x"87",x"c4",x"f0"),
   397 => (x"d0",x"e9",x"c0",x"86"),
   398 => (x"d8",x"f1",x"c3",x"48"),
   399 => (x"20",x"41",x"20",x"49"),
   400 => (x"20",x"41",x"20",x"41"),
   401 => (x"20",x"41",x"20",x"41"),
   402 => (x"10",x"41",x"20",x"41"),
   403 => (x"10",x"51",x"10",x"51"),
   404 => (x"a6",x"e0",x"c0",x"51"),
   405 => (x"78",x"66",x"c4",x"48"),
   406 => (x"48",x"d8",x"cf",x"c1"),
   407 => (x"c1",x"78",x"66",x"c4"),
   408 => (x"c1",x"4a",x"73",x"83"),
   409 => (x"bf",x"97",x"e4",x"cf"),
   410 => (x"06",x"aa",x"b7",x"49"),
   411 => (x"c0",x"87",x"e9",x"fe"),
   412 => (x"d8",x"48",x"66",x"e0"),
   413 => (x"e4",x"c0",x"90",x"66"),
   414 => (x"1e",x"72",x"58",x"a6"),
   415 => (x"66",x"cc",x"49",x"70"),
   416 => (x"87",x"d3",x"f4",x"4a"),
   417 => (x"a6",x"dc",x"4a",x"26"),
   418 => (x"66",x"e0",x"c0",x"58"),
   419 => (x"89",x"66",x"c8",x"49"),
   420 => (x"48",x"71",x"91",x"c7"),
   421 => (x"c0",x"88",x"66",x"d8"),
   422 => (x"6e",x"58",x"a6",x"e4"),
   423 => (x"82",x"ca",x"4a",x"bf"),
   424 => (x"97",x"e0",x"cf",x"c1"),
   425 => (x"c1",x"c1",x"49",x"bf"),
   426 => (x"cc",x"c0",x"05",x"a9"),
   427 => (x"72",x"8a",x"c1",x"87"),
   428 => (x"d8",x"cf",x"c1",x"48"),
   429 => (x"08",x"6e",x"88",x"bf"),
   430 => (x"48",x"66",x"c4",x"78"),
   431 => (x"a6",x"c8",x"80",x"c1"),
   432 => (x"e8",x"e7",x"c0",x"58"),
   433 => (x"06",x"a8",x"b7",x"bf"),
   434 => (x"c3",x"87",x"e8",x"f7"),
   435 => (x"ff",x"48",x"c4",x"ef"),
   436 => (x"c0",x"78",x"bf",x"c8"),
   437 => (x"f1",x"1e",x"e8",x"f0"),
   438 => (x"f0",x"c0",x"87",x"c9"),
   439 => (x"c2",x"f1",x"1e",x"f8"),
   440 => (x"fc",x"f0",x"c0",x"87"),
   441 => (x"87",x"fb",x"f0",x"1e"),
   442 => (x"1e",x"f4",x"f1",x"c0"),
   443 => (x"c1",x"87",x"f4",x"f0"),
   444 => (x"1e",x"bf",x"d8",x"cf"),
   445 => (x"1e",x"f8",x"f1",x"c0"),
   446 => (x"c5",x"87",x"e8",x"f0"),
   447 => (x"d4",x"f2",x"c0",x"1e"),
   448 => (x"87",x"df",x"f0",x"1e"),
   449 => (x"bf",x"dc",x"cf",x"c1"),
   450 => (x"f0",x"f2",x"c0",x"1e"),
   451 => (x"87",x"d3",x"f0",x"1e"),
   452 => (x"f3",x"c0",x"1e",x"c1"),
   453 => (x"ca",x"f0",x"1e",x"cc"),
   454 => (x"e0",x"cf",x"c1",x"87"),
   455 => (x"1e",x"49",x"bf",x"97"),
   456 => (x"1e",x"e8",x"f3",x"c0"),
   457 => (x"c1",x"87",x"fc",x"ef"),
   458 => (x"f4",x"c0",x"1e",x"c1"),
   459 => (x"f2",x"ef",x"1e",x"c4"),
   460 => (x"e4",x"cf",x"c1",x"87"),
   461 => (x"1e",x"49",x"bf",x"97"),
   462 => (x"1e",x"e0",x"f4",x"c0"),
   463 => (x"c1",x"87",x"e4",x"ef"),
   464 => (x"f4",x"c0",x"1e",x"c2"),
   465 => (x"da",x"ef",x"1e",x"fc"),
   466 => (x"c8",x"d0",x"c1",x"87"),
   467 => (x"f5",x"c0",x"1e",x"bf"),
   468 => (x"ce",x"ef",x"1e",x"d8"),
   469 => (x"c0",x"1e",x"c7",x"87"),
   470 => (x"ef",x"1e",x"f4",x"f5"),
   471 => (x"ec",x"c1",x"87",x"c5"),
   472 => (x"c0",x"1e",x"bf",x"cc"),
   473 => (x"ee",x"1e",x"d0",x"f6"),
   474 => (x"f6",x"c0",x"87",x"f9"),
   475 => (x"f2",x"ee",x"1e",x"ec"),
   476 => (x"d8",x"f7",x"c0",x"87"),
   477 => (x"87",x"eb",x"ee",x"1e"),
   478 => (x"bf",x"d0",x"cf",x"c1"),
   479 => (x"f7",x"c0",x"1e",x"bf"),
   480 => (x"de",x"ee",x"1e",x"e4"),
   481 => (x"c0",x"f8",x"c0",x"87"),
   482 => (x"87",x"d7",x"ee",x"1e"),
   483 => (x"bf",x"d0",x"cf",x"c1"),
   484 => (x"69",x"81",x"c4",x"49"),
   485 => (x"f4",x"f8",x"c0",x"1e"),
   486 => (x"87",x"c7",x"ee",x"1e"),
   487 => (x"f9",x"c0",x"1e",x"c0"),
   488 => (x"fe",x"ed",x"1e",x"d0"),
   489 => (x"d0",x"cf",x"c1",x"87"),
   490 => (x"81",x"c8",x"49",x"bf"),
   491 => (x"f9",x"c0",x"1e",x"69"),
   492 => (x"ee",x"ed",x"1e",x"ec"),
   493 => (x"c0",x"1e",x"c2",x"87"),
   494 => (x"ed",x"1e",x"c8",x"fa"),
   495 => (x"cf",x"c1",x"87",x"e5"),
   496 => (x"cc",x"49",x"bf",x"d0"),
   497 => (x"c0",x"1e",x"69",x"81"),
   498 => (x"ed",x"1e",x"e4",x"fa"),
   499 => (x"1e",x"d1",x"87",x"d5"),
   500 => (x"1e",x"c0",x"fb",x"c0"),
   501 => (x"c1",x"87",x"cc",x"ed"),
   502 => (x"49",x"bf",x"d0",x"cf"),
   503 => (x"1e",x"71",x"81",x"d0"),
   504 => (x"1e",x"dc",x"fb",x"c0"),
   505 => (x"c0",x"87",x"fc",x"ec"),
   506 => (x"ec",x"1e",x"f8",x"fb"),
   507 => (x"fc",x"c0",x"87",x"f5"),
   508 => (x"ee",x"ec",x"1e",x"f0"),
   509 => (x"d4",x"cf",x"c1",x"87"),
   510 => (x"c0",x"1e",x"bf",x"bf"),
   511 => (x"ec",x"1e",x"c4",x"fd"),
   512 => (x"fd",x"c0",x"87",x"e1"),
   513 => (x"da",x"ec",x"1e",x"e0"),
   514 => (x"d4",x"cf",x"c1",x"87"),
   515 => (x"81",x"c4",x"49",x"bf"),
   516 => (x"fe",x"c0",x"1e",x"69"),
   517 => (x"ca",x"ec",x"1e",x"e0"),
   518 => (x"c0",x"1e",x"c0",x"87"),
   519 => (x"ec",x"1e",x"fc",x"fe"),
   520 => (x"cf",x"c1",x"87",x"c1"),
   521 => (x"c8",x"49",x"bf",x"d4"),
   522 => (x"c0",x"1e",x"69",x"81"),
   523 => (x"eb",x"1e",x"d8",x"ff"),
   524 => (x"1e",x"c1",x"87",x"f1"),
   525 => (x"1e",x"f4",x"ff",x"c0"),
   526 => (x"c1",x"87",x"e8",x"eb"),
   527 => (x"49",x"bf",x"d4",x"cf"),
   528 => (x"1e",x"69",x"81",x"cc"),
   529 => (x"1e",x"d0",x"c0",x"c1"),
   530 => (x"d2",x"87",x"d8",x"eb"),
   531 => (x"ec",x"c0",x"c1",x"1e"),
   532 => (x"87",x"cf",x"eb",x"1e"),
   533 => (x"bf",x"d4",x"cf",x"c1"),
   534 => (x"71",x"81",x"d0",x"49"),
   535 => (x"c8",x"c1",x"c1",x"1e"),
   536 => (x"87",x"ff",x"ea",x"1e"),
   537 => (x"1e",x"e4",x"c1",x"c1"),
   538 => (x"c4",x"87",x"f8",x"ea"),
   539 => (x"c1",x"1e",x"66",x"dc"),
   540 => (x"ea",x"1e",x"dc",x"c2"),
   541 => (x"1e",x"c5",x"87",x"ed"),
   542 => (x"1e",x"f8",x"c2",x"c1"),
   543 => (x"c4",x"87",x"e4",x"ea"),
   544 => (x"c1",x"1e",x"66",x"f4"),
   545 => (x"ea",x"1e",x"d4",x"c3"),
   546 => (x"1e",x"cd",x"87",x"d9"),
   547 => (x"1e",x"f0",x"c3",x"c1"),
   548 => (x"c4",x"87",x"d0",x"ea"),
   549 => (x"c1",x"1e",x"66",x"ec"),
   550 => (x"ea",x"1e",x"cc",x"c4"),
   551 => (x"1e",x"c7",x"87",x"c5"),
   552 => (x"1e",x"e8",x"c4",x"c1"),
   553 => (x"c5",x"87",x"fc",x"e9"),
   554 => (x"c1",x"1e",x"66",x"c4"),
   555 => (x"e9",x"1e",x"c4",x"c5"),
   556 => (x"1e",x"c1",x"87",x"f1"),
   557 => (x"1e",x"e0",x"c5",x"c1"),
   558 => (x"c3",x"87",x"e8",x"e9"),
   559 => (x"c1",x"1e",x"f8",x"f0"),
   560 => (x"e9",x"1e",x"fc",x"c5"),
   561 => (x"c6",x"c1",x"87",x"dd"),
   562 => (x"d6",x"e9",x"1e",x"d8"),
   563 => (x"d8",x"f1",x"c3",x"87"),
   564 => (x"d0",x"c7",x"c1",x"1e"),
   565 => (x"87",x"cb",x"e9",x"1e"),
   566 => (x"1e",x"ec",x"c7",x"c1"),
   567 => (x"c1",x"87",x"c4",x"e9"),
   568 => (x"e8",x"1e",x"e4",x"c8"),
   569 => (x"ef",x"c3",x"87",x"fd"),
   570 => (x"c3",x"49",x"bf",x"c4"),
   571 => (x"89",x"bf",x"c0",x"ef"),
   572 => (x"59",x"cc",x"ef",x"c3"),
   573 => (x"c8",x"c1",x"1e",x"71"),
   574 => (x"e6",x"e8",x"1e",x"e8"),
   575 => (x"86",x"e8",x"c5",x"87"),
   576 => (x"bf",x"c8",x"ef",x"c3"),
   577 => (x"b7",x"f8",x"c1",x"48"),
   578 => (x"d7",x"c0",x"03",x"a8"),
   579 => (x"d0",x"ea",x"c0",x"87"),
   580 => (x"87",x"cf",x"e8",x"1e"),
   581 => (x"1e",x"c8",x"eb",x"c0"),
   582 => (x"c0",x"87",x"c8",x"e8"),
   583 => (x"e8",x"1e",x"e8",x"eb"),
   584 => (x"86",x"cc",x"87",x"c1"),
   585 => (x"bf",x"c8",x"ef",x"c3"),
   586 => (x"e8",x"cf",x"4a",x"49"),
   587 => (x"72",x"1e",x"71",x"92"),
   588 => (x"c0",x"49",x"72",x"1e"),
   589 => (x"4a",x"bf",x"e8",x"e7"),
   590 => (x"26",x"87",x"dc",x"e9"),
   591 => (x"c3",x"49",x"26",x"4a"),
   592 => (x"c0",x"58",x"d0",x"ef"),
   593 => (x"4a",x"bf",x"e8",x"e7"),
   594 => (x"93",x"e8",x"cf",x"4b"),
   595 => (x"1e",x"72",x"1e",x"71"),
   596 => (x"e9",x"4a",x"09",x"73"),
   597 => (x"4a",x"26",x"87",x"c1"),
   598 => (x"ef",x"c3",x"49",x"26"),
   599 => (x"f9",x"c8",x"58",x"d4"),
   600 => (x"72",x"1e",x"71",x"92"),
   601 => (x"4a",x"09",x"72",x"1e"),
   602 => (x"26",x"87",x"ec",x"e8"),
   603 => (x"c3",x"49",x"26",x"4a"),
   604 => (x"c0",x"58",x"d8",x"ef"),
   605 => (x"e6",x"1e",x"ec",x"eb"),
   606 => (x"ef",x"c3",x"87",x"e9"),
   607 => (x"c0",x"1e",x"bf",x"cc"),
   608 => (x"e6",x"1e",x"dc",x"ec"),
   609 => (x"ec",x"c0",x"87",x"dd"),
   610 => (x"d6",x"e6",x"1e",x"e4"),
   611 => (x"d0",x"ef",x"c3",x"87"),
   612 => (x"ed",x"c0",x"1e",x"bf"),
   613 => (x"ca",x"e6",x"1e",x"d4"),
   614 => (x"d4",x"ef",x"c3",x"87"),
   615 => (x"ed",x"c0",x"1e",x"bf"),
   616 => (x"fe",x"e5",x"1e",x"dc"),
   617 => (x"fc",x"ed",x"c0",x"87"),
   618 => (x"87",x"f7",x"e5",x"1e"),
   619 => (x"f8",x"fe",x"48",x"c0"),
   620 => (x"26",x"4d",x"26",x"8e"),
   621 => (x"26",x"4b",x"26",x"4c"),
   622 => (x"4a",x"71",x"1e",x"4f"),
   623 => (x"bf",x"d0",x"cf",x"c1"),
   624 => (x"c1",x"87",x"c6",x"02"),
   625 => (x"bf",x"bf",x"d0",x"cf"),
   626 => (x"d0",x"cf",x"c1",x"7a"),
   627 => (x"81",x"cc",x"49",x"bf"),
   628 => (x"cf",x"c1",x"1e",x"71"),
   629 => (x"ca",x"1e",x"bf",x"d8"),
   630 => (x"f7",x"e2",x"c0",x"49"),
   631 => (x"26",x"8e",x"f8",x"87"),
   632 => (x"00",x"00",x"00",x"4f"),
   633 => (x"00",x"00",x"00",x"00"),
   634 => (x"00",x"00",x"61",x"a8"),
   635 => (x"67",x"6f",x"72",x"50"),
   636 => (x"20",x"6d",x"61",x"72"),
   637 => (x"70",x"6d",x"6f",x"63"),
   638 => (x"64",x"65",x"6c",x"69"),
   639 => (x"74",x"69",x"77",x"20"),
   640 => (x"72",x"27",x"20",x"68"),
   641 => (x"73",x"69",x"67",x"65"),
   642 => (x"27",x"72",x"65",x"74"),
   643 => (x"74",x"74",x"61",x"20"),
   644 => (x"75",x"62",x"69",x"72"),
   645 => (x"00",x"0a",x"65",x"74"),
   646 => (x"00",x"00",x"00",x"0a"),
   647 => (x"67",x"6f",x"72",x"50"),
   648 => (x"20",x"6d",x"61",x"72"),
   649 => (x"70",x"6d",x"6f",x"63"),
   650 => (x"64",x"65",x"6c",x"69"),
   651 => (x"74",x"69",x"77",x"20"),
   652 => (x"74",x"75",x"6f",x"68"),
   653 => (x"65",x"72",x"27",x"20"),
   654 => (x"74",x"73",x"69",x"67"),
   655 => (x"20",x"27",x"72",x"65"),
   656 => (x"72",x"74",x"74",x"61"),
   657 => (x"74",x"75",x"62",x"69"),
   658 => (x"00",x"00",x"0a",x"65"),
   659 => (x"00",x"00",x"00",x"0a"),
   660 => (x"59",x"52",x"48",x"44"),
   661 => (x"4e",x"4f",x"54",x"53"),
   662 => (x"52",x"50",x"20",x"45"),
   663 => (x"41",x"52",x"47",x"4f"),
   664 => (x"33",x"20",x"2c",x"4d"),
   665 => (x"20",x"44",x"52",x"27"),
   666 => (x"49",x"52",x"54",x"53"),
   667 => (x"00",x"00",x"47",x"4e"),
   668 => (x"59",x"52",x"48",x"44"),
   669 => (x"4e",x"4f",x"54",x"53"),
   670 => (x"52",x"50",x"20",x"45"),
   671 => (x"41",x"52",x"47",x"4f"),
   672 => (x"32",x"20",x"2c",x"4d"),
   673 => (x"20",x"44",x"4e",x"27"),
   674 => (x"49",x"52",x"54",x"53"),
   675 => (x"00",x"00",x"47",x"4e"),
   676 => (x"73",x"61",x"65",x"4d"),
   677 => (x"64",x"65",x"72",x"75"),
   678 => (x"6d",x"69",x"74",x"20"),
   679 => (x"6f",x"74",x"20",x"65"),
   680 => (x"6d",x"73",x"20",x"6f"),
   681 => (x"20",x"6c",x"6c",x"61"),
   682 => (x"6f",x"20",x"6f",x"74"),
   683 => (x"69",x"61",x"74",x"62"),
   684 => (x"65",x"6d",x"20",x"6e"),
   685 => (x"6e",x"69",x"6e",x"61"),
   686 => (x"6c",x"75",x"66",x"67"),
   687 => (x"73",x"65",x"72",x"20"),
   688 => (x"73",x"74",x"6c",x"75"),
   689 => (x"00",x"00",x"00",x"0a"),
   690 => (x"61",x"65",x"6c",x"50"),
   691 => (x"69",x"20",x"65",x"73"),
   692 => (x"65",x"72",x"63",x"6e"),
   693 => (x"20",x"65",x"73",x"61"),
   694 => (x"62",x"6d",x"75",x"6e"),
   695 => (x"6f",x"20",x"72",x"65"),
   696 => (x"75",x"72",x"20",x"66"),
   697 => (x"00",x"0a",x"73",x"6e"),
   698 => (x"00",x"00",x"00",x"0a"),
   699 => (x"72",x"63",x"69",x"4d"),
   700 => (x"63",x"65",x"73",x"6f"),
   701 => (x"73",x"64",x"6e",x"6f"),
   702 => (x"72",x"6f",x"66",x"20"),
   703 => (x"65",x"6e",x"6f",x"20"),
   704 => (x"6e",x"75",x"72",x"20"),
   705 => (x"72",x"68",x"74",x"20"),
   706 => (x"68",x"67",x"75",x"6f"),
   707 => (x"72",x"68",x"44",x"20"),
   708 => (x"6f",x"74",x"73",x"79"),
   709 => (x"20",x"3a",x"65",x"6e"),
   710 => (x"00",x"00",x"00",x"00"),
   711 => (x"0a",x"20",x"64",x"25"),
   712 => (x"00",x"00",x"00",x"00"),
   713 => (x"79",x"72",x"68",x"44"),
   714 => (x"6e",x"6f",x"74",x"73"),
   715 => (x"70",x"20",x"73",x"65"),
   716 => (x"53",x"20",x"72",x"65"),
   717 => (x"6e",x"6f",x"63",x"65"),
   718 => (x"20",x"20",x"3a",x"64"),
   719 => (x"20",x"20",x"20",x"20"),
   720 => (x"20",x"20",x"20",x"20"),
   721 => (x"20",x"20",x"20",x"20"),
   722 => (x"20",x"20",x"20",x"20"),
   723 => (x"20",x"20",x"20",x"20"),
   724 => (x"00",x"00",x"00",x"00"),
   725 => (x"0a",x"20",x"64",x"25"),
   726 => (x"00",x"00",x"00",x"00"),
   727 => (x"20",x"58",x"41",x"56"),
   728 => (x"53",x"50",x"49",x"4d"),
   729 => (x"74",x"61",x"72",x"20"),
   730 => (x"20",x"67",x"6e",x"69"),
   731 => (x"30",x"31",x"20",x"2a"),
   732 => (x"3d",x"20",x"30",x"30"),
   733 => (x"20",x"64",x"25",x"20"),
   734 => (x"00",x"00",x"00",x"0a"),
   735 => (x"00",x"00",x"00",x"0a"),
   736 => (x"59",x"52",x"48",x"44"),
   737 => (x"4e",x"4f",x"54",x"53"),
   738 => (x"52",x"50",x"20",x"45"),
   739 => (x"41",x"52",x"47",x"4f"),
   740 => (x"53",x"20",x"2c",x"4d"),
   741 => (x"20",x"45",x"4d",x"4f"),
   742 => (x"49",x"52",x"54",x"53"),
   743 => (x"00",x"00",x"47",x"4e"),
   744 => (x"59",x"52",x"48",x"44"),
   745 => (x"4e",x"4f",x"54",x"53"),
   746 => (x"52",x"50",x"20",x"45"),
   747 => (x"41",x"52",x"47",x"4f"),
   748 => (x"31",x"20",x"2c",x"4d"),
   749 => (x"20",x"54",x"53",x"27"),
   750 => (x"49",x"52",x"54",x"53"),
   751 => (x"00",x"00",x"47",x"4e"),
   752 => (x"00",x"00",x"00",x"0a"),
   753 => (x"79",x"72",x"68",x"44"),
   754 => (x"6e",x"6f",x"74",x"73"),
   755 => (x"65",x"42",x"20",x"65"),
   756 => (x"6d",x"68",x"63",x"6e"),
   757 => (x"2c",x"6b",x"72",x"61"),
   758 => (x"72",x"65",x"56",x"20"),
   759 => (x"6e",x"6f",x"69",x"73"),
   760 => (x"31",x"2e",x"32",x"20"),
   761 => (x"61",x"4c",x"28",x"20"),
   762 => (x"61",x"75",x"67",x"6e"),
   763 => (x"20",x"3a",x"65",x"67"),
   764 => (x"00",x"0a",x"29",x"43"),
   765 => (x"00",x"00",x"00",x"0a"),
   766 => (x"63",x"65",x"78",x"45"),
   767 => (x"6f",x"69",x"74",x"75"),
   768 => (x"74",x"73",x"20",x"6e"),
   769 => (x"73",x"74",x"72",x"61"),
   770 => (x"64",x"25",x"20",x"2c"),
   771 => (x"6e",x"75",x"72",x"20"),
   772 => (x"68",x"74",x"20",x"73"),
   773 => (x"67",x"75",x"6f",x"72"),
   774 => (x"68",x"44",x"20",x"68"),
   775 => (x"74",x"73",x"79",x"72"),
   776 => (x"0a",x"65",x"6e",x"6f"),
   777 => (x"00",x"00",x"00",x"00"),
   778 => (x"63",x"65",x"78",x"45"),
   779 => (x"6f",x"69",x"74",x"75"),
   780 => (x"6e",x"65",x"20",x"6e"),
   781 => (x"00",x"0a",x"73",x"64"),
   782 => (x"00",x"00",x"00",x"0a"),
   783 => (x"61",x"6e",x"69",x"46"),
   784 => (x"61",x"76",x"20",x"6c"),
   785 => (x"73",x"65",x"75",x"6c"),
   786 => (x"20",x"66",x"6f",x"20"),
   787 => (x"20",x"65",x"68",x"74"),
   788 => (x"69",x"72",x"61",x"76"),
   789 => (x"65",x"6c",x"62",x"61"),
   790 => (x"73",x"75",x"20",x"73"),
   791 => (x"69",x"20",x"64",x"65"),
   792 => (x"68",x"74",x"20",x"6e"),
   793 => (x"65",x"62",x"20",x"65"),
   794 => (x"6d",x"68",x"63",x"6e"),
   795 => (x"3a",x"6b",x"72",x"61"),
   796 => (x"00",x"00",x"00",x"0a"),
   797 => (x"00",x"00",x"00",x"0a"),
   798 => (x"5f",x"74",x"6e",x"49"),
   799 => (x"62",x"6f",x"6c",x"47"),
   800 => (x"20",x"20",x"20",x"3a"),
   801 => (x"20",x"20",x"20",x"20"),
   802 => (x"20",x"20",x"20",x"20"),
   803 => (x"0a",x"64",x"25",x"20"),
   804 => (x"00",x"00",x"00",x"00"),
   805 => (x"20",x"20",x"20",x"20"),
   806 => (x"20",x"20",x"20",x"20"),
   807 => (x"75",x"6f",x"68",x"73"),
   808 => (x"62",x"20",x"64",x"6c"),
   809 => (x"20",x"20",x"3a",x"65"),
   810 => (x"0a",x"64",x"25",x"20"),
   811 => (x"00",x"00",x"00",x"00"),
   812 => (x"6c",x"6f",x"6f",x"42"),
   813 => (x"6f",x"6c",x"47",x"5f"),
   814 => (x"20",x"20",x"3a",x"62"),
   815 => (x"20",x"20",x"20",x"20"),
   816 => (x"20",x"20",x"20",x"20"),
   817 => (x"0a",x"64",x"25",x"20"),
   818 => (x"00",x"00",x"00",x"00"),
   819 => (x"20",x"20",x"20",x"20"),
   820 => (x"20",x"20",x"20",x"20"),
   821 => (x"75",x"6f",x"68",x"73"),
   822 => (x"62",x"20",x"64",x"6c"),
   823 => (x"20",x"20",x"3a",x"65"),
   824 => (x"0a",x"64",x"25",x"20"),
   825 => (x"00",x"00",x"00",x"00"),
   826 => (x"31",x"5f",x"68",x"43"),
   827 => (x"6f",x"6c",x"47",x"5f"),
   828 => (x"20",x"20",x"3a",x"62"),
   829 => (x"20",x"20",x"20",x"20"),
   830 => (x"20",x"20",x"20",x"20"),
   831 => (x"0a",x"63",x"25",x"20"),
   832 => (x"00",x"00",x"00",x"00"),
   833 => (x"20",x"20",x"20",x"20"),
   834 => (x"20",x"20",x"20",x"20"),
   835 => (x"75",x"6f",x"68",x"73"),
   836 => (x"62",x"20",x"64",x"6c"),
   837 => (x"20",x"20",x"3a",x"65"),
   838 => (x"0a",x"63",x"25",x"20"),
   839 => (x"00",x"00",x"00",x"00"),
   840 => (x"32",x"5f",x"68",x"43"),
   841 => (x"6f",x"6c",x"47",x"5f"),
   842 => (x"20",x"20",x"3a",x"62"),
   843 => (x"20",x"20",x"20",x"20"),
   844 => (x"20",x"20",x"20",x"20"),
   845 => (x"0a",x"63",x"25",x"20"),
   846 => (x"00",x"00",x"00",x"00"),
   847 => (x"20",x"20",x"20",x"20"),
   848 => (x"20",x"20",x"20",x"20"),
   849 => (x"75",x"6f",x"68",x"73"),
   850 => (x"62",x"20",x"64",x"6c"),
   851 => (x"20",x"20",x"3a",x"65"),
   852 => (x"0a",x"63",x"25",x"20"),
   853 => (x"00",x"00",x"00",x"00"),
   854 => (x"5f",x"72",x"72",x"41"),
   855 => (x"6c",x"47",x"5f",x"31"),
   856 => (x"38",x"5b",x"62",x"6f"),
   857 => (x"20",x"20",x"3a",x"5d"),
   858 => (x"20",x"20",x"20",x"20"),
   859 => (x"0a",x"64",x"25",x"20"),
   860 => (x"00",x"00",x"00",x"00"),
   861 => (x"20",x"20",x"20",x"20"),
   862 => (x"20",x"20",x"20",x"20"),
   863 => (x"75",x"6f",x"68",x"73"),
   864 => (x"62",x"20",x"64",x"6c"),
   865 => (x"20",x"20",x"3a",x"65"),
   866 => (x"0a",x"64",x"25",x"20"),
   867 => (x"00",x"00",x"00",x"00"),
   868 => (x"5f",x"72",x"72",x"41"),
   869 => (x"6c",x"47",x"5f",x"32"),
   870 => (x"38",x"5b",x"62",x"6f"),
   871 => (x"5d",x"37",x"5b",x"5d"),
   872 => (x"20",x"20",x"20",x"3a"),
   873 => (x"0a",x"64",x"25",x"20"),
   874 => (x"00",x"00",x"00",x"00"),
   875 => (x"20",x"20",x"20",x"20"),
   876 => (x"20",x"20",x"20",x"20"),
   877 => (x"75",x"6f",x"68",x"73"),
   878 => (x"62",x"20",x"64",x"6c"),
   879 => (x"20",x"20",x"3a",x"65"),
   880 => (x"6d",x"75",x"4e",x"20"),
   881 => (x"5f",x"72",x"65",x"62"),
   882 => (x"52",x"5f",x"66",x"4f"),
   883 => (x"20",x"73",x"6e",x"75"),
   884 => (x"30",x"31",x"20",x"2b"),
   885 => (x"00",x"00",x"00",x"0a"),
   886 => (x"5f",x"72",x"74",x"50"),
   887 => (x"62",x"6f",x"6c",x"47"),
   888 => (x"00",x"0a",x"3e",x"2d"),
   889 => (x"74",x"50",x"20",x"20"),
   890 => (x"6f",x"43",x"5f",x"72"),
   891 => (x"20",x"3a",x"70",x"6d"),
   892 => (x"20",x"20",x"20",x"20"),
   893 => (x"20",x"20",x"20",x"20"),
   894 => (x"0a",x"64",x"25",x"20"),
   895 => (x"00",x"00",x"00",x"00"),
   896 => (x"20",x"20",x"20",x"20"),
   897 => (x"20",x"20",x"20",x"20"),
   898 => (x"75",x"6f",x"68",x"73"),
   899 => (x"62",x"20",x"64",x"6c"),
   900 => (x"20",x"20",x"3a",x"65"),
   901 => (x"6d",x"69",x"28",x"20"),
   902 => (x"6d",x"65",x"6c",x"70"),
   903 => (x"61",x"74",x"6e",x"65"),
   904 => (x"6e",x"6f",x"69",x"74"),
   905 => (x"70",x"65",x"64",x"2d"),
   906 => (x"65",x"64",x"6e",x"65"),
   907 => (x"0a",x"29",x"74",x"6e"),
   908 => (x"00",x"00",x"00",x"00"),
   909 => (x"69",x"44",x"20",x"20"),
   910 => (x"3a",x"72",x"63",x"73"),
   911 => (x"20",x"20",x"20",x"20"),
   912 => (x"20",x"20",x"20",x"20"),
   913 => (x"20",x"20",x"20",x"20"),
   914 => (x"0a",x"64",x"25",x"20"),
   915 => (x"00",x"00",x"00",x"00"),
   916 => (x"20",x"20",x"20",x"20"),
   917 => (x"20",x"20",x"20",x"20"),
   918 => (x"75",x"6f",x"68",x"73"),
   919 => (x"62",x"20",x"64",x"6c"),
   920 => (x"20",x"20",x"3a",x"65"),
   921 => (x"0a",x"64",x"25",x"20"),
   922 => (x"00",x"00",x"00",x"00"),
   923 => (x"6e",x"45",x"20",x"20"),
   924 => (x"43",x"5f",x"6d",x"75"),
   925 => (x"3a",x"70",x"6d",x"6f"),
   926 => (x"20",x"20",x"20",x"20"),
   927 => (x"20",x"20",x"20",x"20"),
   928 => (x"0a",x"64",x"25",x"20"),
   929 => (x"00",x"00",x"00",x"00"),
   930 => (x"20",x"20",x"20",x"20"),
   931 => (x"20",x"20",x"20",x"20"),
   932 => (x"75",x"6f",x"68",x"73"),
   933 => (x"62",x"20",x"64",x"6c"),
   934 => (x"20",x"20",x"3a",x"65"),
   935 => (x"0a",x"64",x"25",x"20"),
   936 => (x"00",x"00",x"00",x"00"),
   937 => (x"6e",x"49",x"20",x"20"),
   938 => (x"6f",x"43",x"5f",x"74"),
   939 => (x"20",x"3a",x"70",x"6d"),
   940 => (x"20",x"20",x"20",x"20"),
   941 => (x"20",x"20",x"20",x"20"),
   942 => (x"0a",x"64",x"25",x"20"),
   943 => (x"00",x"00",x"00",x"00"),
   944 => (x"20",x"20",x"20",x"20"),
   945 => (x"20",x"20",x"20",x"20"),
   946 => (x"75",x"6f",x"68",x"73"),
   947 => (x"62",x"20",x"64",x"6c"),
   948 => (x"20",x"20",x"3a",x"65"),
   949 => (x"0a",x"64",x"25",x"20"),
   950 => (x"00",x"00",x"00",x"00"),
   951 => (x"74",x"53",x"20",x"20"),
   952 => (x"6f",x"43",x"5f",x"72"),
   953 => (x"20",x"3a",x"70",x"6d"),
   954 => (x"20",x"20",x"20",x"20"),
   955 => (x"20",x"20",x"20",x"20"),
   956 => (x"0a",x"73",x"25",x"20"),
   957 => (x"00",x"00",x"00",x"00"),
   958 => (x"20",x"20",x"20",x"20"),
   959 => (x"20",x"20",x"20",x"20"),
   960 => (x"75",x"6f",x"68",x"73"),
   961 => (x"62",x"20",x"64",x"6c"),
   962 => (x"20",x"20",x"3a",x"65"),
   963 => (x"52",x"48",x"44",x"20"),
   964 => (x"4f",x"54",x"53",x"59"),
   965 => (x"50",x"20",x"45",x"4e"),
   966 => (x"52",x"47",x"4f",x"52"),
   967 => (x"20",x"2c",x"4d",x"41"),
   968 => (x"45",x"4d",x"4f",x"53"),
   969 => (x"52",x"54",x"53",x"20"),
   970 => (x"0a",x"47",x"4e",x"49"),
   971 => (x"00",x"00",x"00",x"00"),
   972 => (x"74",x"78",x"65",x"4e"),
   973 => (x"72",x"74",x"50",x"5f"),
   974 => (x"6f",x"6c",x"47",x"5f"),
   975 => (x"0a",x"3e",x"2d",x"62"),
   976 => (x"00",x"00",x"00",x"00"),
   977 => (x"74",x"50",x"20",x"20"),
   978 => (x"6f",x"43",x"5f",x"72"),
   979 => (x"20",x"3a",x"70",x"6d"),
   980 => (x"20",x"20",x"20",x"20"),
   981 => (x"20",x"20",x"20",x"20"),
   982 => (x"0a",x"64",x"25",x"20"),
   983 => (x"00",x"00",x"00",x"00"),
   984 => (x"20",x"20",x"20",x"20"),
   985 => (x"20",x"20",x"20",x"20"),
   986 => (x"75",x"6f",x"68",x"73"),
   987 => (x"62",x"20",x"64",x"6c"),
   988 => (x"20",x"20",x"3a",x"65"),
   989 => (x"6d",x"69",x"28",x"20"),
   990 => (x"6d",x"65",x"6c",x"70"),
   991 => (x"61",x"74",x"6e",x"65"),
   992 => (x"6e",x"6f",x"69",x"74"),
   993 => (x"70",x"65",x"64",x"2d"),
   994 => (x"65",x"64",x"6e",x"65"),
   995 => (x"2c",x"29",x"74",x"6e"),
   996 => (x"6d",x"61",x"73",x"20"),
   997 => (x"73",x"61",x"20",x"65"),
   998 => (x"6f",x"62",x"61",x"20"),
   999 => (x"00",x"0a",x"65",x"76"),
  1000 => (x"69",x"44",x"20",x"20"),
  1001 => (x"3a",x"72",x"63",x"73"),
  1002 => (x"20",x"20",x"20",x"20"),
  1003 => (x"20",x"20",x"20",x"20"),
  1004 => (x"20",x"20",x"20",x"20"),
  1005 => (x"0a",x"64",x"25",x"20"),
  1006 => (x"00",x"00",x"00",x"00"),
  1007 => (x"20",x"20",x"20",x"20"),
  1008 => (x"20",x"20",x"20",x"20"),
  1009 => (x"75",x"6f",x"68",x"73"),
  1010 => (x"62",x"20",x"64",x"6c"),
  1011 => (x"20",x"20",x"3a",x"65"),
  1012 => (x"0a",x"64",x"25",x"20"),
  1013 => (x"00",x"00",x"00",x"00"),
  1014 => (x"6e",x"45",x"20",x"20"),
  1015 => (x"43",x"5f",x"6d",x"75"),
  1016 => (x"3a",x"70",x"6d",x"6f"),
  1017 => (x"20",x"20",x"20",x"20"),
  1018 => (x"20",x"20",x"20",x"20"),
  1019 => (x"0a",x"64",x"25",x"20"),
  1020 => (x"00",x"00",x"00",x"00"),
  1021 => (x"20",x"20",x"20",x"20"),
  1022 => (x"20",x"20",x"20",x"20"),
  1023 => (x"75",x"6f",x"68",x"73"),
  1024 => (x"62",x"20",x"64",x"6c"),
  1025 => (x"20",x"20",x"3a",x"65"),
  1026 => (x"0a",x"64",x"25",x"20"),
  1027 => (x"00",x"00",x"00",x"00"),
  1028 => (x"6e",x"49",x"20",x"20"),
  1029 => (x"6f",x"43",x"5f",x"74"),
  1030 => (x"20",x"3a",x"70",x"6d"),
  1031 => (x"20",x"20",x"20",x"20"),
  1032 => (x"20",x"20",x"20",x"20"),
  1033 => (x"0a",x"64",x"25",x"20"),
  1034 => (x"00",x"00",x"00",x"00"),
  1035 => (x"20",x"20",x"20",x"20"),
  1036 => (x"20",x"20",x"20",x"20"),
  1037 => (x"75",x"6f",x"68",x"73"),
  1038 => (x"62",x"20",x"64",x"6c"),
  1039 => (x"20",x"20",x"3a",x"65"),
  1040 => (x"0a",x"64",x"25",x"20"),
  1041 => (x"00",x"00",x"00",x"00"),
  1042 => (x"74",x"53",x"20",x"20"),
  1043 => (x"6f",x"43",x"5f",x"72"),
  1044 => (x"20",x"3a",x"70",x"6d"),
  1045 => (x"20",x"20",x"20",x"20"),
  1046 => (x"20",x"20",x"20",x"20"),
  1047 => (x"0a",x"73",x"25",x"20"),
  1048 => (x"00",x"00",x"00",x"00"),
  1049 => (x"20",x"20",x"20",x"20"),
  1050 => (x"20",x"20",x"20",x"20"),
  1051 => (x"75",x"6f",x"68",x"73"),
  1052 => (x"62",x"20",x"64",x"6c"),
  1053 => (x"20",x"20",x"3a",x"65"),
  1054 => (x"52",x"48",x"44",x"20"),
  1055 => (x"4f",x"54",x"53",x"59"),
  1056 => (x"50",x"20",x"45",x"4e"),
  1057 => (x"52",x"47",x"4f",x"52"),
  1058 => (x"20",x"2c",x"4d",x"41"),
  1059 => (x"45",x"4d",x"4f",x"53"),
  1060 => (x"52",x"54",x"53",x"20"),
  1061 => (x"0a",x"47",x"4e",x"49"),
  1062 => (x"00",x"00",x"00",x"00"),
  1063 => (x"5f",x"74",x"6e",x"49"),
  1064 => (x"6f",x"4c",x"5f",x"31"),
  1065 => (x"20",x"20",x"3a",x"63"),
  1066 => (x"20",x"20",x"20",x"20"),
  1067 => (x"20",x"20",x"20",x"20"),
  1068 => (x"0a",x"64",x"25",x"20"),
  1069 => (x"00",x"00",x"00",x"00"),
  1070 => (x"20",x"20",x"20",x"20"),
  1071 => (x"20",x"20",x"20",x"20"),
  1072 => (x"75",x"6f",x"68",x"73"),
  1073 => (x"62",x"20",x"64",x"6c"),
  1074 => (x"20",x"20",x"3a",x"65"),
  1075 => (x"0a",x"64",x"25",x"20"),
  1076 => (x"00",x"00",x"00",x"00"),
  1077 => (x"5f",x"74",x"6e",x"49"),
  1078 => (x"6f",x"4c",x"5f",x"32"),
  1079 => (x"20",x"20",x"3a",x"63"),
  1080 => (x"20",x"20",x"20",x"20"),
  1081 => (x"20",x"20",x"20",x"20"),
  1082 => (x"0a",x"64",x"25",x"20"),
  1083 => (x"00",x"00",x"00",x"00"),
  1084 => (x"20",x"20",x"20",x"20"),
  1085 => (x"20",x"20",x"20",x"20"),
  1086 => (x"75",x"6f",x"68",x"73"),
  1087 => (x"62",x"20",x"64",x"6c"),
  1088 => (x"20",x"20",x"3a",x"65"),
  1089 => (x"0a",x"64",x"25",x"20"),
  1090 => (x"00",x"00",x"00",x"00"),
  1091 => (x"5f",x"74",x"6e",x"49"),
  1092 => (x"6f",x"4c",x"5f",x"33"),
  1093 => (x"20",x"20",x"3a",x"63"),
  1094 => (x"20",x"20",x"20",x"20"),
  1095 => (x"20",x"20",x"20",x"20"),
  1096 => (x"0a",x"64",x"25",x"20"),
  1097 => (x"00",x"00",x"00",x"00"),
  1098 => (x"20",x"20",x"20",x"20"),
  1099 => (x"20",x"20",x"20",x"20"),
  1100 => (x"75",x"6f",x"68",x"73"),
  1101 => (x"62",x"20",x"64",x"6c"),
  1102 => (x"20",x"20",x"3a",x"65"),
  1103 => (x"0a",x"64",x"25",x"20"),
  1104 => (x"00",x"00",x"00",x"00"),
  1105 => (x"6d",x"75",x"6e",x"45"),
  1106 => (x"63",x"6f",x"4c",x"5f"),
  1107 => (x"20",x"20",x"20",x"3a"),
  1108 => (x"20",x"20",x"20",x"20"),
  1109 => (x"20",x"20",x"20",x"20"),
  1110 => (x"0a",x"64",x"25",x"20"),
  1111 => (x"00",x"00",x"00",x"00"),
  1112 => (x"20",x"20",x"20",x"20"),
  1113 => (x"20",x"20",x"20",x"20"),
  1114 => (x"75",x"6f",x"68",x"73"),
  1115 => (x"62",x"20",x"64",x"6c"),
  1116 => (x"20",x"20",x"3a",x"65"),
  1117 => (x"0a",x"64",x"25",x"20"),
  1118 => (x"00",x"00",x"00",x"00"),
  1119 => (x"5f",x"72",x"74",x"53"),
  1120 => (x"6f",x"4c",x"5f",x"31"),
  1121 => (x"20",x"20",x"3a",x"63"),
  1122 => (x"20",x"20",x"20",x"20"),
  1123 => (x"20",x"20",x"20",x"20"),
  1124 => (x"0a",x"73",x"25",x"20"),
  1125 => (x"00",x"00",x"00",x"00"),
  1126 => (x"20",x"20",x"20",x"20"),
  1127 => (x"20",x"20",x"20",x"20"),
  1128 => (x"75",x"6f",x"68",x"73"),
  1129 => (x"62",x"20",x"64",x"6c"),
  1130 => (x"20",x"20",x"3a",x"65"),
  1131 => (x"52",x"48",x"44",x"20"),
  1132 => (x"4f",x"54",x"53",x"59"),
  1133 => (x"50",x"20",x"45",x"4e"),
  1134 => (x"52",x"47",x"4f",x"52"),
  1135 => (x"20",x"2c",x"4d",x"41"),
  1136 => (x"54",x"53",x"27",x"31"),
  1137 => (x"52",x"54",x"53",x"20"),
  1138 => (x"0a",x"47",x"4e",x"49"),
  1139 => (x"00",x"00",x"00",x"00"),
  1140 => (x"5f",x"72",x"74",x"53"),
  1141 => (x"6f",x"4c",x"5f",x"32"),
  1142 => (x"20",x"20",x"3a",x"63"),
  1143 => (x"20",x"20",x"20",x"20"),
  1144 => (x"20",x"20",x"20",x"20"),
  1145 => (x"0a",x"73",x"25",x"20"),
  1146 => (x"00",x"00",x"00",x"00"),
  1147 => (x"20",x"20",x"20",x"20"),
  1148 => (x"20",x"20",x"20",x"20"),
  1149 => (x"75",x"6f",x"68",x"73"),
  1150 => (x"62",x"20",x"64",x"6c"),
  1151 => (x"20",x"20",x"3a",x"65"),
  1152 => (x"52",x"48",x"44",x"20"),
  1153 => (x"4f",x"54",x"53",x"59"),
  1154 => (x"50",x"20",x"45",x"4e"),
  1155 => (x"52",x"47",x"4f",x"52"),
  1156 => (x"20",x"2c",x"4d",x"41"),
  1157 => (x"44",x"4e",x"27",x"32"),
  1158 => (x"52",x"54",x"53",x"20"),
  1159 => (x"0a",x"47",x"4e",x"49"),
  1160 => (x"00",x"00",x"00",x"00"),
  1161 => (x"00",x"00",x"00",x"0a"),
  1162 => (x"72",x"65",x"73",x"55"),
  1163 => (x"6d",x"69",x"74",x"20"),
  1164 => (x"25",x"20",x"3a",x"65"),
  1165 => (x"1e",x"00",x"0a",x"64"),
  1166 => (x"1e",x"74",x"1e",x"73"),
  1167 => (x"66",x"cc",x"4b",x"71"),
  1168 => (x"c2",x"7a",x"73",x"4a"),
  1169 => (x"87",x"c4",x"05",x"ab"),
  1170 => (x"87",x"c2",x"4c",x"c1"),
  1171 => (x"9c",x"74",x"4c",x"c0"),
  1172 => (x"c3",x"87",x"c2",x"05"),
  1173 => (x"02",x"9b",x"73",x"7a"),
  1174 => (x"c1",x"49",x"87",x"d6"),
  1175 => (x"87",x"d4",x"02",x"89"),
  1176 => (x"e3",x"c0",x"02",x"89"),
  1177 => (x"c0",x"02",x"89",x"87"),
  1178 => (x"02",x"89",x"87",x"e4"),
  1179 => (x"87",x"de",x"87",x"de"),
  1180 => (x"87",x"da",x"7a",x"c0"),
  1181 => (x"bf",x"d8",x"cf",x"c1"),
  1182 => (x"b7",x"e4",x"c1",x"48"),
  1183 => (x"87",x"c4",x"06",x"a8"),
  1184 => (x"87",x"ca",x"7a",x"c0"),
  1185 => (x"87",x"c6",x"7a",x"c3"),
  1186 => (x"87",x"c2",x"7a",x"c1"),
  1187 => (x"4c",x"26",x"7a",x"c2"),
  1188 => (x"4f",x"26",x"4b",x"26"),
  1189 => (x"49",x"4a",x"71",x"1e"),
  1190 => (x"66",x"c4",x"81",x"c2"),
  1191 => (x"c8",x"80",x"71",x"48"),
  1192 => (x"26",x"78",x"08",x"66"),
  1193 => (x"5b",x"5e",x"0e",x"4f"),
  1194 => (x"f4",x"0e",x"5d",x"5c"),
  1195 => (x"59",x"a6",x"c4",x"86"),
  1196 => (x"4c",x"66",x"e0",x"c0"),
  1197 => (x"48",x"74",x"84",x"c5"),
  1198 => (x"a6",x"c8",x"90",x"c4"),
  1199 => (x"70",x"4d",x"6e",x"58"),
  1200 => (x"66",x"e4",x"c0",x"85"),
  1201 => (x"49",x"a5",x"c4",x"7d"),
  1202 => (x"79",x"66",x"e4",x"c0"),
  1203 => (x"49",x"a5",x"f8",x"c1"),
  1204 => (x"a6",x"c8",x"79",x"74"),
  1205 => (x"78",x"a4",x"c1",x"48"),
  1206 => (x"dd",x"01",x"ac",x"b7"),
  1207 => (x"c3",x"49",x"74",x"87"),
  1208 => (x"66",x"dc",x"91",x"c8"),
  1209 => (x"c4",x"82",x"71",x"4a"),
  1210 => (x"66",x"c8",x"82",x"66"),
  1211 => (x"c1",x"8b",x"74",x"4b"),
  1212 => (x"c4",x"7a",x"74",x"83"),
  1213 => (x"01",x"8b",x"c1",x"82"),
  1214 => (x"49",x"74",x"87",x"f7"),
  1215 => (x"dc",x"91",x"c8",x"c3"),
  1216 => (x"4a",x"71",x"81",x"66"),
  1217 => (x"c4",x"82",x"66",x"c4"),
  1218 => (x"c1",x"48",x"6a",x"8a"),
  1219 => (x"c0",x"7a",x"70",x"80"),
  1220 => (x"c4",x"81",x"e0",x"fe"),
  1221 => (x"79",x"6d",x"81",x"66"),
  1222 => (x"48",x"d8",x"cf",x"c1"),
  1223 => (x"8e",x"f4",x"78",x"c5"),
  1224 => (x"4c",x"26",x"4d",x"26"),
  1225 => (x"4f",x"26",x"4b",x"26"),
  1226 => (x"74",x"1e",x"73",x"1e"),
  1227 => (x"4c",x"4b",x"71",x"1e"),
  1228 => (x"49",x"66",x"cc",x"4a"),
  1229 => (x"c4",x"02",x"aa",x"b7"),
  1230 => (x"c7",x"48",x"c0",x"87"),
  1231 => (x"e4",x"cf",x"c1",x"87"),
  1232 => (x"48",x"c1",x"5c",x"97"),
  1233 => (x"4b",x"26",x"4c",x"26"),
  1234 => (x"5e",x"0e",x"4f",x"26"),
  1235 => (x"0e",x"5d",x"5c",x"5b"),
  1236 => (x"a6",x"c4",x"86",x"f4"),
  1237 => (x"dc",x"4d",x"c2",x"59"),
  1238 => (x"81",x"c1",x"49",x"66"),
  1239 => (x"84",x"c2",x"4c",x"6e"),
  1240 => (x"49",x"6b",x"4b",x"a1"),
  1241 => (x"c4",x"99",x"ff",x"c3"),
  1242 => (x"50",x"6c",x"48",x"a6"),
  1243 => (x"4a",x"66",x"97",x"c4"),
  1244 => (x"02",x"aa",x"b7",x"71"),
  1245 => (x"a6",x"c8",x"87",x"c7"),
  1246 => (x"cd",x"78",x"c0",x"48"),
  1247 => (x"e0",x"cf",x"c1",x"87"),
  1248 => (x"66",x"97",x"c4",x"48"),
  1249 => (x"48",x"a6",x"c8",x"50"),
  1250 => (x"66",x"c8",x"78",x"c1"),
  1251 => (x"c1",x"87",x"c4",x"05"),
  1252 => (x"c2",x"84",x"83",x"85"),
  1253 => (x"ff",x"06",x"ad",x"b7"),
  1254 => (x"4a",x"6e",x"87",x"c8"),
  1255 => (x"fe",x"49",x"66",x"dc"),
  1256 => (x"c0",x"87",x"ef",x"fe"),
  1257 => (x"cb",x"06",x"a8",x"b7"),
  1258 => (x"d8",x"cf",x"c1",x"87"),
  1259 => (x"78",x"a5",x"c7",x"48"),
  1260 => (x"87",x"c2",x"48",x"c1"),
  1261 => (x"8e",x"f4",x"48",x"c0"),
  1262 => (x"4c",x"26",x"4d",x"26"),
  1263 => (x"4f",x"26",x"4b",x"26"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
