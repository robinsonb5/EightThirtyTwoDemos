
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"44",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"36"),
    10 => (x"c0",x"c0",x"c2",x"4f"),
    11 => (x"15",x"01",x"27",x"4e"),
    12 => (x"00",x"0f",x"00",x"00"),
    13 => (x"f0",x"c1",x"87",x"fd"),
    14 => (x"43",x"27",x"4e",x"c0"),
    15 => (x"0f",x"00",x"00",x"00"),
    16 => (x"4f",x"87",x"fd",x"00"),
    17 => (x"ff",x"1e",x"1e",x"4f"),
    18 => (x"48",x"69",x"49",x"c0"),
    19 => (x"c4",x"98",x"c0",x"c4"),
    20 => (x"02",x"6e",x"58",x"a6"),
    21 => (x"c8",x"87",x"f3",x"ff"),
    22 => (x"26",x"48",x"79",x"66"),
    23 => (x"87",x"c6",x"c0",x"c0"),
    24 => (x"4c",x"26",x"4d",x"26"),
    25 => (x"4f",x"26",x"4b",x"26"),
    26 => (x"5c",x"5b",x"5e",x"0e"),
    27 => (x"4c",x"66",x"cc",x"0e"),
    28 => (x"4a",x"14",x"4b",x"c0"),
    29 => (x"72",x"9a",x"ff",x"c3"),
    30 => (x"d9",x"c0",x"02",x"9a"),
    31 => (x"71",x"49",x"72",x"87"),
    32 => (x"00",x"45",x"27",x"1e"),
    33 => (x"c4",x"0f",x"00",x"00"),
    34 => (x"14",x"83",x"c1",x"86"),
    35 => (x"9a",x"ff",x"c3",x"4a"),
    36 => (x"ff",x"05",x"9a",x"72"),
    37 => (x"48",x"73",x"87",x"e7"),
    38 => (x"87",x"c6",x"ff",x"ff"),
    39 => (x"5c",x"5b",x"5e",x"0e"),
    40 => (x"86",x"f0",x"0e",x"5d"),
    41 => (x"a6",x"c4",x"4b",x"c0"),
    42 => (x"c0",x"78",x"c0",x"48"),
    43 => (x"c0",x"4c",x"a6",x"e4"),
    44 => (x"48",x"49",x"66",x"e0"),
    45 => (x"e4",x"c0",x"80",x"c1"),
    46 => (x"4a",x"11",x"58",x"a6"),
    47 => (x"ba",x"82",x"c0",x"fe"),
    48 => (x"c4",x"02",x"9a",x"72"),
    49 => (x"66",x"c4",x"87",x"ee"),
    50 => (x"87",x"f8",x"c3",x"02"),
    51 => (x"c0",x"48",x"a6",x"c4"),
    52 => (x"c0",x"49",x"72",x"78"),
    53 => (x"c3",x"02",x"aa",x"f0"),
    54 => (x"e3",x"c1",x"87",x"c0"),
    55 => (x"c1",x"c3",x"02",x"a9"),
    56 => (x"a9",x"e4",x"c1",x"87"),
    57 => (x"87",x"e3",x"c0",x"02"),
    58 => (x"02",x"a9",x"ec",x"c1"),
    59 => (x"c1",x"87",x"eb",x"c2"),
    60 => (x"c0",x"02",x"a9",x"f0"),
    61 => (x"f3",x"c1",x"87",x"d5"),
    62 => (x"c7",x"c2",x"02",x"a9"),
    63 => (x"a9",x"f5",x"c1",x"87"),
    64 => (x"87",x"c7",x"c0",x"02"),
    65 => (x"05",x"a9",x"f8",x"c1"),
    66 => (x"c4",x"87",x"ec",x"c2"),
    67 => (x"c4",x"49",x"74",x"84"),
    68 => (x"69",x"48",x"76",x"89"),
    69 => (x"c1",x"02",x"6e",x"78"),
    70 => (x"a6",x"c8",x"87",x"da"),
    71 => (x"cc",x"78",x"c0",x"48"),
    72 => (x"78",x"c0",x"48",x"a6"),
    73 => (x"b7",x"dc",x"49",x"6e"),
    74 => (x"cf",x"4a",x"71",x"29"),
    75 => (x"c4",x"48",x"6e",x"9a"),
    76 => (x"72",x"58",x"a6",x"30"),
    77 => (x"c5",x"c0",x"02",x"9a"),
    78 => (x"48",x"a6",x"c8",x"87"),
    79 => (x"aa",x"c9",x"78",x"c1"),
    80 => (x"87",x"c6",x"c0",x"06"),
    81 => (x"c0",x"82",x"f7",x"c0"),
    82 => (x"f0",x"c0",x"87",x"c3"),
    83 => (x"02",x"66",x"c8",x"82"),
    84 => (x"72",x"87",x"cc",x"c0"),
    85 => (x"00",x"45",x"27",x"1e"),
    86 => (x"c4",x"0f",x"00",x"00"),
    87 => (x"cc",x"83",x"c1",x"86"),
    88 => (x"80",x"c1",x"48",x"66"),
    89 => (x"cc",x"58",x"a6",x"d0"),
    90 => (x"b7",x"c8",x"48",x"66"),
    91 => (x"f3",x"fe",x"04",x"a8"),
    92 => (x"87",x"e9",x"c1",x"87"),
    93 => (x"27",x"1e",x"f0",x"c0"),
    94 => (x"00",x"00",x"00",x"45"),
    95 => (x"c1",x"86",x"c4",x"0f"),
    96 => (x"87",x"d9",x"c1",x"83"),
    97 => (x"49",x"74",x"84",x"c4"),
    98 => (x"1e",x"69",x"89",x"c4"),
    99 => (x"00",x"00",x"68",x"27"),
   100 => (x"86",x"c4",x"0f",x"00"),
   101 => (x"c1",x"83",x"49",x"70"),
   102 => (x"a6",x"c4",x"87",x"c3"),
   103 => (x"c0",x"78",x"c1",x"48"),
   104 => (x"84",x"c4",x"87",x"fb"),
   105 => (x"89",x"c4",x"49",x"74"),
   106 => (x"45",x"27",x"1e",x"69"),
   107 => (x"0f",x"00",x"00",x"00"),
   108 => (x"83",x"c1",x"86",x"c4"),
   109 => (x"72",x"87",x"e6",x"c0"),
   110 => (x"00",x"45",x"27",x"1e"),
   111 => (x"c4",x"0f",x"00",x"00"),
   112 => (x"87",x"d9",x"c0",x"86"),
   113 => (x"05",x"aa",x"e5",x"c0"),
   114 => (x"c4",x"87",x"c8",x"c0"),
   115 => (x"78",x"c1",x"48",x"a6"),
   116 => (x"72",x"87",x"ca",x"c0"),
   117 => (x"00",x"45",x"27",x"1e"),
   118 => (x"c4",x"0f",x"00",x"00"),
   119 => (x"66",x"e0",x"c0",x"86"),
   120 => (x"80",x"c1",x"48",x"49"),
   121 => (x"58",x"a6",x"e4",x"c0"),
   122 => (x"c0",x"fe",x"4a",x"11"),
   123 => (x"9a",x"72",x"ba",x"82"),
   124 => (x"87",x"d2",x"fb",x"05"),
   125 => (x"8e",x"f0",x"48",x"73"),
   126 => (x"4c",x"26",x"4d",x"26"),
   127 => (x"4f",x"26",x"4b",x"26"),
   128 => (x"00",x"00",x"00",x"00"),
   129 => (x"ff",x"1e",x"75",x"1e"),
   130 => (x"ff",x"c3",x"4d",x"d4"),
   131 => (x"48",x"6d",x"7d",x"49"),
   132 => (x"7d",x"71",x"38",x"c8"),
   133 => (x"38",x"c8",x"b0",x"6d"),
   134 => (x"b0",x"6d",x"7d",x"71"),
   135 => (x"7d",x"71",x"38",x"c8"),
   136 => (x"38",x"c8",x"b0",x"6d"),
   137 => (x"4f",x"26",x"4d",x"26"),
   138 => (x"ff",x"1e",x"75",x"1e"),
   139 => (x"ff",x"c3",x"4d",x"d4"),
   140 => (x"48",x"6d",x"7d",x"49"),
   141 => (x"7d",x"71",x"30",x"c8"),
   142 => (x"30",x"c8",x"b0",x"6d"),
   143 => (x"b0",x"6d",x"7d",x"71"),
   144 => (x"7d",x"71",x"30",x"c8"),
   145 => (x"4d",x"26",x"b0",x"6d"),
   146 => (x"75",x"1e",x"4f",x"26"),
   147 => (x"4d",x"d4",x"ff",x"1e"),
   148 => (x"c8",x"49",x"66",x"cc"),
   149 => (x"fe",x"7d",x"48",x"66"),
   150 => (x"c9",x"02",x"67",x"e6"),
   151 => (x"39",x"d8",x"07",x"31"),
   152 => (x"39",x"09",x"7d",x"09"),
   153 => (x"39",x"09",x"7d",x"09"),
   154 => (x"39",x"09",x"7d",x"09"),
   155 => (x"38",x"d0",x"7d",x"09"),
   156 => (x"f1",x"c9",x"7d",x"70"),
   157 => (x"ff",x"c3",x"49",x"c0"),
   158 => (x"a8",x"08",x"6d",x"48"),
   159 => (x"08",x"87",x"c7",x"05"),
   160 => (x"05",x"89",x"c1",x"7d"),
   161 => (x"4d",x"26",x"87",x"f3"),
   162 => (x"ff",x"1e",x"4f",x"26"),
   163 => (x"c8",x"c3",x"49",x"d4"),
   164 => (x"80",x"79",x"ff",x"48"),
   165 => (x"26",x"87",x"fa",x"05"),
   166 => (x"5a",x"5e",x"0e",x"4f"),
   167 => (x"0e",x"5d",x"5c",x"5b"),
   168 => (x"c1",x"f0",x"ff",x"c0"),
   169 => (x"c0",x"c1",x"4d",x"f7"),
   170 => (x"c0",x"c0",x"c0",x"c0"),
   171 => (x"02",x"8a",x"27",x"4b"),
   172 => (x"c4",x"0f",x"00",x"00"),
   173 => (x"c0",x"4c",x"df",x"f8"),
   174 => (x"27",x"1e",x"75",x"1e"),
   175 => (x"00",x"00",x"02",x"4a"),
   176 => (x"70",x"86",x"c8",x"0f"),
   177 => (x"aa",x"b7",x"c1",x"4a"),
   178 => (x"87",x"ef",x"c0",x"05"),
   179 => (x"c3",x"49",x"d4",x"ff"),
   180 => (x"1e",x"73",x"79",x"ff"),
   181 => (x"c1",x"f0",x"e1",x"c0"),
   182 => (x"4a",x"27",x"1e",x"e9"),
   183 => (x"0f",x"00",x"00",x"02"),
   184 => (x"4a",x"70",x"86",x"c8"),
   185 => (x"c0",x"05",x"9a",x"72"),
   186 => (x"d4",x"ff",x"87",x"cb"),
   187 => (x"79",x"ff",x"c3",x"49"),
   188 => (x"d0",x"c0",x"48",x"c1"),
   189 => (x"02",x"8a",x"27",x"87"),
   190 => (x"c1",x"0f",x"00",x"00"),
   191 => (x"05",x"9c",x"74",x"8c"),
   192 => (x"c0",x"87",x"f4",x"fe"),
   193 => (x"26",x"4d",x"26",x"48"),
   194 => (x"26",x"4b",x"26",x"4c"),
   195 => (x"0e",x"4f",x"26",x"4a"),
   196 => (x"5c",x"5b",x"5a",x"5e"),
   197 => (x"f0",x"ff",x"c0",x"0e"),
   198 => (x"ff",x"4c",x"c1",x"c1"),
   199 => (x"ff",x"c3",x"49",x"d4"),
   200 => (x"16",x"41",x"27",x"79"),
   201 => (x"27",x"1e",x"00",x"00"),
   202 => (x"00",x"00",x"00",x"68"),
   203 => (x"d3",x"86",x"c4",x"0f"),
   204 => (x"74",x"1e",x"c0",x"4b"),
   205 => (x"02",x"4a",x"27",x"1e"),
   206 => (x"c8",x"0f",x"00",x"00"),
   207 => (x"72",x"4a",x"70",x"86"),
   208 => (x"cb",x"c0",x"05",x"9a"),
   209 => (x"49",x"d4",x"ff",x"87"),
   210 => (x"c1",x"79",x"ff",x"c3"),
   211 => (x"87",x"d0",x"c0",x"48"),
   212 => (x"00",x"02",x"8a",x"27"),
   213 => (x"8b",x"c1",x"0f",x"00"),
   214 => (x"ff",x"05",x"9b",x"73"),
   215 => (x"48",x"c0",x"87",x"d3"),
   216 => (x"4b",x"26",x"4c",x"26"),
   217 => (x"4f",x"26",x"4a",x"26"),
   218 => (x"5b",x"5a",x"5e",x"0e"),
   219 => (x"1e",x"0e",x"5d",x"5c"),
   220 => (x"ff",x"4d",x"ff",x"c3"),
   221 => (x"8a",x"27",x"4c",x"d4"),
   222 => (x"0f",x"00",x"00",x"02"),
   223 => (x"c0",x"1e",x"ea",x"c6"),
   224 => (x"c8",x"c1",x"f0",x"e1"),
   225 => (x"02",x"4a",x"27",x"1e"),
   226 => (x"c8",x"0f",x"00",x"00"),
   227 => (x"72",x"4a",x"70",x"86"),
   228 => (x"04",x"c7",x"27",x"1e"),
   229 => (x"27",x"1e",x"00",x"00"),
   230 => (x"00",x"00",x"00",x"9c"),
   231 => (x"c1",x"86",x"c8",x"0f"),
   232 => (x"c0",x"02",x"aa",x"b7"),
   233 => (x"0f",x"27",x"87",x"cb"),
   234 => (x"0f",x"00",x"00",x"03"),
   235 => (x"c9",x"c3",x"48",x"c0"),
   236 => (x"02",x"28",x"27",x"87"),
   237 => (x"70",x"0f",x"00",x"00"),
   238 => (x"ff",x"ff",x"cf",x"4a"),
   239 => (x"b7",x"ea",x"c6",x"9a"),
   240 => (x"cb",x"c0",x"02",x"aa"),
   241 => (x"03",x"0f",x"27",x"87"),
   242 => (x"c0",x"0f",x"00",x"00"),
   243 => (x"87",x"ea",x"c2",x"48"),
   244 => (x"49",x"76",x"7c",x"75"),
   245 => (x"27",x"79",x"f1",x"c0"),
   246 => (x"00",x"00",x"02",x"99"),
   247 => (x"72",x"4a",x"70",x"0f"),
   248 => (x"eb",x"c1",x"02",x"9a"),
   249 => (x"c0",x"1e",x"c0",x"87"),
   250 => (x"fa",x"c1",x"f0",x"ff"),
   251 => (x"02",x"4a",x"27",x"1e"),
   252 => (x"c8",x"0f",x"00",x"00"),
   253 => (x"73",x"4b",x"70",x"86"),
   254 => (x"c3",x"c1",x"05",x"9b"),
   255 => (x"27",x"1e",x"73",x"87"),
   256 => (x"00",x"00",x"04",x"85"),
   257 => (x"00",x"9c",x"27",x"1e"),
   258 => (x"c8",x"0f",x"00",x"00"),
   259 => (x"6c",x"7c",x"75",x"86"),
   260 => (x"73",x"9b",x"75",x"4b"),
   261 => (x"04",x"91",x"27",x"1e"),
   262 => (x"27",x"1e",x"00",x"00"),
   263 => (x"00",x"00",x"00",x"9c"),
   264 => (x"75",x"86",x"c8",x"0f"),
   265 => (x"75",x"7c",x"75",x"7c"),
   266 => (x"73",x"7c",x"75",x"7c"),
   267 => (x"9a",x"c0",x"c1",x"4a"),
   268 => (x"c0",x"02",x"9a",x"72"),
   269 => (x"48",x"c1",x"87",x"c5"),
   270 => (x"c0",x"87",x"ff",x"c0"),
   271 => (x"87",x"fa",x"c0",x"48"),
   272 => (x"9f",x"27",x"1e",x"73"),
   273 => (x"1e",x"00",x"00",x"04"),
   274 => (x"00",x"00",x"9c",x"27"),
   275 => (x"86",x"c8",x"0f",x"00"),
   276 => (x"b7",x"c2",x"49",x"6e"),
   277 => (x"d3",x"c0",x"05",x"a9"),
   278 => (x"04",x"ab",x"27",x"87"),
   279 => (x"27",x"1e",x"00",x"00"),
   280 => (x"00",x"00",x"00",x"9c"),
   281 => (x"c0",x"86",x"c4",x"0f"),
   282 => (x"87",x"ce",x"c0",x"48"),
   283 => (x"88",x"c1",x"48",x"6e"),
   284 => (x"6e",x"58",x"a6",x"c4"),
   285 => (x"87",x"df",x"fd",x"05"),
   286 => (x"26",x"26",x"48",x"c0"),
   287 => (x"26",x"4c",x"26",x"4d"),
   288 => (x"26",x"4a",x"26",x"4b"),
   289 => (x"44",x"4d",x"43",x"4f"),
   290 => (x"25",x"20",x"38",x"35"),
   291 => (x"20",x"20",x"0a",x"64"),
   292 => (x"44",x"4d",x"43",x"00"),
   293 => (x"32",x"5f",x"38",x"35"),
   294 => (x"0a",x"64",x"25",x"20"),
   295 => (x"43",x"00",x"20",x"20"),
   296 => (x"38",x"35",x"44",x"4d"),
   297 => (x"0a",x"64",x"25",x"20"),
   298 => (x"53",x"00",x"20",x"20"),
   299 => (x"20",x"43",x"48",x"44"),
   300 => (x"74",x"69",x"6e",x"49"),
   301 => (x"69",x"6c",x"61",x"69"),
   302 => (x"69",x"74",x"61",x"7a"),
   303 => (x"65",x"20",x"6e",x"6f"),
   304 => (x"72",x"6f",x"72",x"72"),
   305 => (x"63",x"00",x"0a",x"21"),
   306 => (x"43",x"5f",x"64",x"6d"),
   307 => (x"20",x"38",x"44",x"4d"),
   308 => (x"70",x"73",x"65",x"72"),
   309 => (x"65",x"73",x"6e",x"6f"),
   310 => (x"64",x"25",x"20",x"3a"),
   311 => (x"5e",x"0e",x"00",x"0a"),
   312 => (x"5d",x"5c",x"5b",x"5a"),
   313 => (x"d0",x"ff",x"1e",x"0e"),
   314 => (x"c0",x"c0",x"c8",x"4c"),
   315 => (x"02",x"00",x"27",x"4b"),
   316 => (x"c1",x"49",x"00",x"00"),
   317 => (x"05",x"fb",x"27",x"79"),
   318 => (x"27",x"1e",x"00",x"00"),
   319 => (x"00",x"00",x"00",x"68"),
   320 => (x"c7",x"86",x"c4",x"0f"),
   321 => (x"73",x"48",x"6c",x"4d"),
   322 => (x"58",x"a6",x"c4",x"98"),
   323 => (x"cc",x"c0",x"02",x"6e"),
   324 => (x"73",x"48",x"6c",x"87"),
   325 => (x"58",x"a6",x"c4",x"98"),
   326 => (x"f4",x"ff",x"05",x"6e"),
   327 => (x"27",x"7c",x"c0",x"87"),
   328 => (x"00",x"00",x"02",x"8a"),
   329 => (x"73",x"48",x"6c",x"0f"),
   330 => (x"58",x"a6",x"c4",x"98"),
   331 => (x"cc",x"c0",x"02",x"6e"),
   332 => (x"73",x"48",x"6c",x"87"),
   333 => (x"58",x"a6",x"c4",x"98"),
   334 => (x"f4",x"ff",x"05",x"6e"),
   335 => (x"c0",x"7c",x"c1",x"87"),
   336 => (x"d0",x"e5",x"c0",x"1e"),
   337 => (x"27",x"1e",x"c0",x"c1"),
   338 => (x"00",x"00",x"02",x"4a"),
   339 => (x"70",x"86",x"c8",x"0f"),
   340 => (x"aa",x"b7",x"c1",x"4a"),
   341 => (x"87",x"c2",x"c0",x"05"),
   342 => (x"b7",x"c2",x"4d",x"c1"),
   343 => (x"d3",x"c0",x"05",x"ad"),
   344 => (x"05",x"f6",x"27",x"87"),
   345 => (x"27",x"1e",x"00",x"00"),
   346 => (x"00",x"00",x"00",x"68"),
   347 => (x"c0",x"86",x"c4",x"0f"),
   348 => (x"87",x"f7",x"c1",x"48"),
   349 => (x"9d",x"75",x"8d",x"c1"),
   350 => (x"87",x"c9",x"fe",x"05"),
   351 => (x"00",x"03",x"68",x"27"),
   352 => (x"04",x"27",x"0f",x"00"),
   353 => (x"58",x"00",x"00",x"02"),
   354 => (x"00",x"02",x"00",x"27"),
   355 => (x"c0",x"05",x"bf",x"00"),
   356 => (x"1e",x"c1",x"87",x"d0"),
   357 => (x"c1",x"f0",x"ff",x"c0"),
   358 => (x"4a",x"27",x"1e",x"d0"),
   359 => (x"0f",x"00",x"00",x"02"),
   360 => (x"d4",x"ff",x"86",x"c8"),
   361 => (x"79",x"ff",x"c3",x"49"),
   362 => (x"00",x"08",x"91",x"27"),
   363 => (x"e0",x"27",x"0f",x"00"),
   364 => (x"58",x"00",x"00",x"17"),
   365 => (x"00",x"17",x"dc",x"27"),
   366 => (x"27",x"1e",x"bf",x"00"),
   367 => (x"00",x"00",x"05",x"ff"),
   368 => (x"00",x"9c",x"27",x"1e"),
   369 => (x"c8",x"0f",x"00",x"00"),
   370 => (x"73",x"48",x"6c",x"86"),
   371 => (x"58",x"a6",x"c4",x"98"),
   372 => (x"cc",x"c0",x"02",x"6e"),
   373 => (x"73",x"48",x"6c",x"87"),
   374 => (x"58",x"a6",x"c4",x"98"),
   375 => (x"f4",x"ff",x"05",x"6e"),
   376 => (x"ff",x"7c",x"c0",x"87"),
   377 => (x"ff",x"c3",x"49",x"d4"),
   378 => (x"26",x"48",x"c1",x"79"),
   379 => (x"4c",x"26",x"4d",x"26"),
   380 => (x"4a",x"26",x"4b",x"26"),
   381 => (x"45",x"49",x"4f",x"26"),
   382 => (x"53",x"00",x"52",x"52"),
   383 => (x"53",x"00",x"49",x"50"),
   384 => (x"61",x"63",x"20",x"44"),
   385 => (x"73",x"20",x"64",x"72"),
   386 => (x"20",x"65",x"7a",x"69"),
   387 => (x"25",x"20",x"73",x"69"),
   388 => (x"0e",x"00",x"0a",x"64"),
   389 => (x"5c",x"5b",x"5a",x"5e"),
   390 => (x"c3",x"1e",x"0e",x"5d"),
   391 => (x"d4",x"ff",x"4d",x"ff"),
   392 => (x"ff",x"7c",x"75",x"4c"),
   393 => (x"c8",x"48",x"bf",x"d0"),
   394 => (x"c4",x"98",x"c0",x"c0"),
   395 => (x"02",x"6e",x"58",x"a6"),
   396 => (x"c8",x"87",x"d2",x"c0"),
   397 => (x"ff",x"4a",x"c0",x"c0"),
   398 => (x"72",x"48",x"bf",x"d0"),
   399 => (x"58",x"a6",x"c4",x"98"),
   400 => (x"f2",x"ff",x"05",x"6e"),
   401 => (x"49",x"d0",x"ff",x"87"),
   402 => (x"75",x"79",x"c1",x"c4"),
   403 => (x"1e",x"66",x"d8",x"7c"),
   404 => (x"c1",x"f0",x"ff",x"c0"),
   405 => (x"4a",x"27",x"1e",x"d8"),
   406 => (x"0f",x"00",x"00",x"02"),
   407 => (x"4a",x"70",x"86",x"c8"),
   408 => (x"c0",x"02",x"9a",x"72"),
   409 => (x"1b",x"27",x"87",x"d3"),
   410 => (x"1e",x"00",x"00",x"07"),
   411 => (x"00",x"00",x"68",x"27"),
   412 => (x"86",x"c4",x"0f",x"00"),
   413 => (x"d7",x"c2",x"48",x"c1"),
   414 => (x"c3",x"7c",x"75",x"87"),
   415 => (x"49",x"76",x"7c",x"fe"),
   416 => (x"66",x"dc",x"79",x"c0"),
   417 => (x"4b",x"72",x"4a",x"bf"),
   418 => (x"73",x"2b",x"b7",x"d8"),
   419 => (x"70",x"98",x"75",x"48"),
   420 => (x"d0",x"4b",x"72",x"7c"),
   421 => (x"48",x"73",x"2b",x"b7"),
   422 => (x"7c",x"70",x"98",x"75"),
   423 => (x"b7",x"c8",x"4b",x"72"),
   424 => (x"75",x"48",x"73",x"2b"),
   425 => (x"72",x"7c",x"70",x"98"),
   426 => (x"70",x"98",x"75",x"48"),
   427 => (x"48",x"66",x"dc",x"7c"),
   428 => (x"e0",x"c0",x"80",x"c4"),
   429 => (x"48",x"6e",x"58",x"a6"),
   430 => (x"a6",x"c4",x"80",x"c1"),
   431 => (x"c2",x"49",x"6e",x"58"),
   432 => (x"04",x"a9",x"b7",x"c0"),
   433 => (x"75",x"87",x"fb",x"fe"),
   434 => (x"75",x"7c",x"75",x"7c"),
   435 => (x"e0",x"da",x"d8",x"7c"),
   436 => (x"6c",x"7c",x"75",x"4b"),
   437 => (x"72",x"9a",x"75",x"4a"),
   438 => (x"c8",x"c0",x"05",x"9a"),
   439 => (x"73",x"8b",x"c1",x"87"),
   440 => (x"ec",x"ff",x"05",x"9b"),
   441 => (x"ff",x"7c",x"75",x"87"),
   442 => (x"c8",x"48",x"bf",x"d0"),
   443 => (x"c4",x"98",x"c0",x"c0"),
   444 => (x"02",x"6e",x"58",x"a6"),
   445 => (x"c8",x"87",x"d2",x"c0"),
   446 => (x"ff",x"4a",x"c0",x"c0"),
   447 => (x"72",x"48",x"bf",x"d0"),
   448 => (x"58",x"a6",x"c4",x"98"),
   449 => (x"f2",x"ff",x"05",x"6e"),
   450 => (x"49",x"d0",x"ff",x"87"),
   451 => (x"48",x"c0",x"79",x"c0"),
   452 => (x"26",x"4d",x"26",x"26"),
   453 => (x"26",x"4b",x"26",x"4c"),
   454 => (x"57",x"4f",x"26",x"4a"),
   455 => (x"65",x"74",x"69",x"72"),
   456 => (x"69",x"61",x"66",x"20"),
   457 => (x"0a",x"64",x"65",x"6c"),
   458 => (x"5a",x"5e",x"0e",x"00"),
   459 => (x"0e",x"5d",x"5c",x"5b"),
   460 => (x"4c",x"66",x"d8",x"1e"),
   461 => (x"76",x"4b",x"66",x"dc"),
   462 => (x"c5",x"79",x"c0",x"49"),
   463 => (x"4d",x"df",x"cd",x"ee"),
   464 => (x"c3",x"49",x"d4",x"ff"),
   465 => (x"d4",x"ff",x"79",x"ff"),
   466 => (x"ff",x"c3",x"4a",x"bf"),
   467 => (x"b7",x"fe",x"c3",x"9a"),
   468 => (x"e5",x"c1",x"05",x"aa"),
   469 => (x"17",x"d8",x"27",x"87"),
   470 => (x"c0",x"49",x"00",x"00"),
   471 => (x"ab",x"b7",x"c4",x"79"),
   472 => (x"87",x"e4",x"c0",x"04"),
   473 => (x"00",x"02",x"04",x"27"),
   474 => (x"4a",x"70",x"0f",x"00"),
   475 => (x"84",x"c4",x"7c",x"72"),
   476 => (x"00",x"17",x"d8",x"27"),
   477 => (x"72",x"48",x"bf",x"00"),
   478 => (x"17",x"dc",x"27",x"80"),
   479 => (x"c4",x"58",x"00",x"00"),
   480 => (x"ab",x"b7",x"c4",x"8b"),
   481 => (x"87",x"dc",x"ff",x"03"),
   482 => (x"06",x"ab",x"b7",x"c0"),
   483 => (x"ff",x"87",x"e5",x"c0"),
   484 => (x"ff",x"c3",x"4d",x"d4"),
   485 => (x"72",x"4a",x"6d",x"7d"),
   486 => (x"84",x"c1",x"7c",x"97"),
   487 => (x"00",x"17",x"d8",x"27"),
   488 => (x"72",x"48",x"bf",x"00"),
   489 => (x"17",x"dc",x"27",x"80"),
   490 => (x"c1",x"58",x"00",x"00"),
   491 => (x"ab",x"b7",x"c0",x"8b"),
   492 => (x"87",x"de",x"ff",x"01"),
   493 => (x"49",x"76",x"4d",x"c1"),
   494 => (x"8d",x"c1",x"79",x"c1"),
   495 => (x"fd",x"05",x"9d",x"75"),
   496 => (x"d4",x"ff",x"87",x"fe"),
   497 => (x"79",x"ff",x"c3",x"49"),
   498 => (x"26",x"26",x"48",x"6e"),
   499 => (x"26",x"4c",x"26",x"4d"),
   500 => (x"26",x"4a",x"26",x"4b"),
   501 => (x"5a",x"5e",x"0e",x"4f"),
   502 => (x"0e",x"5d",x"5c",x"5b"),
   503 => (x"4b",x"d0",x"ff",x"1e"),
   504 => (x"4a",x"c0",x"c0",x"c8"),
   505 => (x"d4",x"ff",x"4c",x"c0"),
   506 => (x"79",x"ff",x"c3",x"49"),
   507 => (x"98",x"72",x"48",x"6b"),
   508 => (x"6e",x"58",x"a6",x"c4"),
   509 => (x"87",x"cc",x"c0",x"02"),
   510 => (x"98",x"72",x"48",x"6b"),
   511 => (x"6e",x"58",x"a6",x"c4"),
   512 => (x"87",x"f4",x"ff",x"05"),
   513 => (x"ff",x"7b",x"c1",x"c4"),
   514 => (x"ff",x"c3",x"49",x"d4"),
   515 => (x"1e",x"66",x"d8",x"79"),
   516 => (x"c1",x"f0",x"ff",x"c0"),
   517 => (x"4a",x"27",x"1e",x"d1"),
   518 => (x"0f",x"00",x"00",x"02"),
   519 => (x"4d",x"70",x"86",x"c8"),
   520 => (x"c0",x"02",x"9d",x"75"),
   521 => (x"1e",x"75",x"87",x"d6"),
   522 => (x"27",x"1e",x"66",x"dc"),
   523 => (x"00",x"00",x"08",x"71"),
   524 => (x"00",x"9c",x"27",x"1e"),
   525 => (x"cc",x"0f",x"00",x"00"),
   526 => (x"87",x"e8",x"c0",x"86"),
   527 => (x"c0",x"1e",x"c0",x"c8"),
   528 => (x"fb",x"1e",x"66",x"e0"),
   529 => (x"86",x"c8",x"87",x"e3"),
   530 => (x"48",x"6b",x"4c",x"70"),
   531 => (x"a6",x"c4",x"98",x"72"),
   532 => (x"c0",x"02",x"6e",x"58"),
   533 => (x"48",x"6b",x"87",x"cc"),
   534 => (x"a6",x"c4",x"98",x"72"),
   535 => (x"ff",x"05",x"6e",x"58"),
   536 => (x"7b",x"c0",x"87",x"f4"),
   537 => (x"26",x"26",x"48",x"74"),
   538 => (x"26",x"4c",x"26",x"4d"),
   539 => (x"26",x"4a",x"26",x"4b"),
   540 => (x"61",x"65",x"52",x"4f"),
   541 => (x"6f",x"63",x"20",x"64"),
   542 => (x"6e",x"61",x"6d",x"6d"),
   543 => (x"61",x"66",x"20",x"64"),
   544 => (x"64",x"65",x"6c",x"69"),
   545 => (x"20",x"74",x"61",x"20"),
   546 => (x"28",x"20",x"64",x"25"),
   547 => (x"0a",x"29",x"64",x"25"),
   548 => (x"5a",x"5e",x"0e",x"00"),
   549 => (x"0e",x"5d",x"5c",x"5b"),
   550 => (x"c0",x"1e",x"c0",x"1e"),
   551 => (x"c9",x"c1",x"f0",x"ff"),
   552 => (x"02",x"4a",x"27",x"1e"),
   553 => (x"c8",x"0f",x"00",x"00"),
   554 => (x"27",x"1e",x"d2",x"86"),
   555 => (x"00",x"00",x"17",x"e8"),
   556 => (x"87",x"f5",x"f9",x"1e"),
   557 => (x"4d",x"c0",x"86",x"c8"),
   558 => (x"b7",x"d2",x"85",x"c1"),
   559 => (x"f7",x"ff",x"04",x"ad"),
   560 => (x"17",x"e8",x"27",x"87"),
   561 => (x"bf",x"97",x"00",x"00"),
   562 => (x"9a",x"c0",x"c3",x"4a"),
   563 => (x"aa",x"b7",x"c0",x"c1"),
   564 => (x"87",x"f2",x"c0",x"05"),
   565 => (x"00",x"17",x"ef",x"27"),
   566 => (x"4a",x"bf",x"97",x"00"),
   567 => (x"f0",x"27",x"32",x"d0"),
   568 => (x"97",x"00",x"00",x"17"),
   569 => (x"33",x"c8",x"4b",x"bf"),
   570 => (x"b2",x"73",x"4a",x"72"),
   571 => (x"00",x"17",x"f1",x"27"),
   572 => (x"4b",x"bf",x"97",x"00"),
   573 => (x"b2",x"73",x"4a",x"72"),
   574 => (x"ff",x"ff",x"ff",x"cf"),
   575 => (x"c1",x"4d",x"72",x"9a"),
   576 => (x"c3",x"35",x"ca",x"85"),
   577 => (x"f1",x"27",x"87",x"cb"),
   578 => (x"97",x"00",x"00",x"17"),
   579 => (x"32",x"c1",x"4a",x"bf"),
   580 => (x"f2",x"27",x"9a",x"c6"),
   581 => (x"97",x"00",x"00",x"17"),
   582 => (x"b7",x"c7",x"4b",x"bf"),
   583 => (x"73",x"4a",x"72",x"2b"),
   584 => (x"17",x"ed",x"27",x"b2"),
   585 => (x"bf",x"97",x"00",x"00"),
   586 => (x"cf",x"48",x"73",x"4b"),
   587 => (x"58",x"a6",x"c4",x"98"),
   588 => (x"00",x"17",x"ee",x"27"),
   589 => (x"4b",x"bf",x"97",x"00"),
   590 => (x"33",x"ca",x"9b",x"c3"),
   591 => (x"00",x"17",x"ef",x"27"),
   592 => (x"4c",x"bf",x"97",x"00"),
   593 => (x"4b",x"73",x"34",x"c2"),
   594 => (x"f0",x"27",x"b3",x"74"),
   595 => (x"97",x"00",x"00",x"17"),
   596 => (x"c0",x"c3",x"4c",x"bf"),
   597 => (x"2c",x"b7",x"c6",x"9c"),
   598 => (x"b3",x"74",x"4b",x"73"),
   599 => (x"66",x"c4",x"1e",x"73"),
   600 => (x"27",x"1e",x"72",x"1e"),
   601 => (x"00",x"00",x"09",x"de"),
   602 => (x"00",x"9c",x"27",x"1e"),
   603 => (x"d0",x"0f",x"00",x"00"),
   604 => (x"c1",x"82",x"c2",x"86"),
   605 => (x"70",x"30",x"72",x"48"),
   606 => (x"27",x"1e",x"72",x"4a"),
   607 => (x"00",x"00",x"0a",x"0b"),
   608 => (x"00",x"9c",x"27",x"1e"),
   609 => (x"c8",x"0f",x"00",x"00"),
   610 => (x"6e",x"48",x"c1",x"86"),
   611 => (x"58",x"a6",x"c4",x"30"),
   612 => (x"4d",x"73",x"83",x"c1"),
   613 => (x"1e",x"6e",x"95",x"72"),
   614 => (x"14",x"27",x"1e",x"75"),
   615 => (x"1e",x"00",x"00",x"0a"),
   616 => (x"00",x"00",x"9c",x"27"),
   617 => (x"86",x"cc",x"0f",x"00"),
   618 => (x"c0",x"c8",x"49",x"6e"),
   619 => (x"c0",x"06",x"a9",x"b7"),
   620 => (x"4a",x"6e",x"87",x"cf"),
   621 => (x"b7",x"c1",x"35",x"c1"),
   622 => (x"b7",x"c0",x"c8",x"2a"),
   623 => (x"f3",x"ff",x"01",x"aa"),
   624 => (x"27",x"1e",x"75",x"87"),
   625 => (x"00",x"00",x"0a",x"2a"),
   626 => (x"00",x"9c",x"27",x"1e"),
   627 => (x"c8",x"0f",x"00",x"00"),
   628 => (x"26",x"48",x"75",x"86"),
   629 => (x"4c",x"26",x"4d",x"26"),
   630 => (x"4a",x"26",x"4b",x"26"),
   631 => (x"5f",x"63",x"4f",x"26"),
   632 => (x"65",x"7a",x"69",x"73"),
   633 => (x"6c",x"75",x"6d",x"5f"),
   634 => (x"25",x"20",x"3a",x"74"),
   635 => (x"72",x"20",x"2c",x"64"),
   636 => (x"5f",x"64",x"61",x"65"),
   637 => (x"6c",x"5f",x"6c",x"62"),
   638 => (x"20",x"3a",x"6e",x"65"),
   639 => (x"20",x"2c",x"64",x"25"),
   640 => (x"7a",x"69",x"73",x"63"),
   641 => (x"25",x"20",x"3a",x"65"),
   642 => (x"4d",x"00",x"0a",x"64"),
   643 => (x"20",x"74",x"6c",x"75"),
   644 => (x"00",x"0a",x"64",x"25"),
   645 => (x"62",x"20",x"64",x"25"),
   646 => (x"6b",x"63",x"6f",x"6c"),
   647 => (x"66",x"6f",x"20",x"73"),
   648 => (x"7a",x"69",x"73",x"20"),
   649 => (x"64",x"25",x"20",x"65"),
   650 => (x"64",x"25",x"00",x"0a"),
   651 => (x"6f",x"6c",x"62",x"20"),
   652 => (x"20",x"73",x"6b",x"63"),
   653 => (x"35",x"20",x"66",x"6f"),
   654 => (x"62",x"20",x"32",x"31"),
   655 => (x"73",x"65",x"74",x"79"),
   656 => (x"5e",x"0e",x"00",x"0a"),
   657 => (x"4b",x"c0",x"0e",x"5b"),
   658 => (x"c0",x"48",x"66",x"d0"),
   659 => (x"c0",x"06",x"a8",x"b7"),
   660 => (x"66",x"c8",x"87",x"f8"),
   661 => (x"fe",x"4a",x"bf",x"97"),
   662 => (x"c8",x"ba",x"82",x"c0"),
   663 => (x"80",x"c1",x"48",x"66"),
   664 => (x"cc",x"58",x"a6",x"cc"),
   665 => (x"49",x"bf",x"97",x"66"),
   666 => (x"b9",x"81",x"c0",x"fe"),
   667 => (x"c1",x"48",x"66",x"cc"),
   668 => (x"58",x"a6",x"d0",x"80"),
   669 => (x"02",x"aa",x"b7",x"71"),
   670 => (x"c1",x"87",x"c5",x"c0"),
   671 => (x"87",x"cc",x"c0",x"48"),
   672 => (x"66",x"d0",x"83",x"c1"),
   673 => (x"ff",x"04",x"ab",x"b7"),
   674 => (x"48",x"c0",x"87",x"c8"),
   675 => (x"87",x"c4",x"c0",x"c0"),
   676 => (x"4c",x"26",x"4d",x"26"),
   677 => (x"4f",x"26",x"4b",x"26"),
   678 => (x"5c",x"5b",x"5e",x"0e"),
   679 => (x"08",x"27",x"0e",x"5d"),
   680 => (x"48",x"00",x"00",x"18"),
   681 => (x"19",x"27",x"78",x"c0"),
   682 => (x"1e",x"00",x"00",x"17"),
   683 => (x"00",x"00",x"68",x"27"),
   684 => (x"86",x"c4",x"0f",x"00"),
   685 => (x"00",x"18",x"48",x"27"),
   686 => (x"1e",x"c0",x"1e",x"00"),
   687 => (x"00",x"07",x"d5",x"27"),
   688 => (x"86",x"c8",x"0f",x"00"),
   689 => (x"c0",x"05",x"98",x"70"),
   690 => (x"45",x"27",x"87",x"d3"),
   691 => (x"1e",x"00",x"00",x"16"),
   692 => (x"00",x"00",x"68",x"27"),
   693 => (x"86",x"c4",x"0f",x"00"),
   694 => (x"d9",x"ce",x"48",x"c0"),
   695 => (x"17",x"26",x"27",x"87"),
   696 => (x"27",x"1e",x"00",x"00"),
   697 => (x"00",x"00",x"00",x"68"),
   698 => (x"c0",x"86",x"c4",x"0f"),
   699 => (x"18",x"34",x"27",x"4b"),
   700 => (x"c1",x"48",x"00",x"00"),
   701 => (x"27",x"1e",x"c8",x"78"),
   702 => (x"00",x"00",x"17",x"3d"),
   703 => (x"18",x"7e",x"27",x"1e"),
   704 => (x"27",x"1e",x"00",x"00"),
   705 => (x"00",x"00",x"0a",x"42"),
   706 => (x"70",x"86",x"cc",x"0f"),
   707 => (x"c8",x"c0",x"05",x"98"),
   708 => (x"18",x"34",x"27",x"87"),
   709 => (x"c0",x"48",x"00",x"00"),
   710 => (x"27",x"1e",x"c8",x"78"),
   711 => (x"00",x"00",x"17",x"46"),
   712 => (x"18",x"9a",x"27",x"1e"),
   713 => (x"27",x"1e",x"00",x"00"),
   714 => (x"00",x"00",x"0a",x"42"),
   715 => (x"70",x"86",x"cc",x"0f"),
   716 => (x"c8",x"c0",x"05",x"98"),
   717 => (x"18",x"34",x"27",x"87"),
   718 => (x"c0",x"48",x"00",x"00"),
   719 => (x"18",x"34",x"27",x"78"),
   720 => (x"1e",x"bf",x"00",x"00"),
   721 => (x"00",x"17",x"4f",x"27"),
   722 => (x"9c",x"27",x"1e",x"00"),
   723 => (x"0f",x"00",x"00",x"00"),
   724 => (x"34",x"27",x"86",x"c8"),
   725 => (x"bf",x"00",x"00",x"18"),
   726 => (x"87",x"fc",x"c2",x"02"),
   727 => (x"00",x"18",x"48",x"27"),
   728 => (x"06",x"27",x"4d",x"00"),
   729 => (x"4c",x"00",x"00",x"1a"),
   730 => (x"00",x"1a",x"46",x"27"),
   731 => (x"49",x"bf",x"9f",x"00"),
   732 => (x"46",x"27",x"1e",x"71"),
   733 => (x"49",x"00",x"00",x"1a"),
   734 => (x"00",x"18",x"48",x"27"),
   735 => (x"1e",x"71",x"89",x"00"),
   736 => (x"c0",x"c8",x"1e",x"d0"),
   737 => (x"16",x"77",x"27",x"1e"),
   738 => (x"27",x"1e",x"00",x"00"),
   739 => (x"00",x"00",x"00",x"9c"),
   740 => (x"74",x"86",x"d4",x"0f"),
   741 => (x"69",x"81",x"c8",x"49"),
   742 => (x"1a",x"46",x"27",x"4b"),
   743 => (x"bf",x"9f",x"00",x"00"),
   744 => (x"ea",x"d6",x"c5",x"49"),
   745 => (x"d3",x"c0",x"05",x"a9"),
   746 => (x"c8",x"49",x"74",x"87"),
   747 => (x"27",x"1e",x"69",x"81"),
   748 => (x"00",x"00",x"11",x"8a"),
   749 => (x"70",x"86",x"c4",x"0f"),
   750 => (x"87",x"e3",x"c0",x"4b"),
   751 => (x"fe",x"c7",x"49",x"75"),
   752 => (x"49",x"69",x"9f",x"81"),
   753 => (x"a9",x"d5",x"e9",x"ca"),
   754 => (x"87",x"d3",x"c0",x"02"),
   755 => (x"00",x"16",x"59",x"27"),
   756 => (x"68",x"27",x"1e",x"00"),
   757 => (x"0f",x"00",x"00",x"00"),
   758 => (x"48",x"c0",x"86",x"c4"),
   759 => (x"73",x"87",x"d7",x"ca"),
   760 => (x"16",x"b4",x"27",x"1e"),
   761 => (x"27",x"1e",x"00",x"00"),
   762 => (x"00",x"00",x"00",x"9c"),
   763 => (x"27",x"86",x"c8",x"0f"),
   764 => (x"00",x"00",x"18",x"48"),
   765 => (x"27",x"1e",x"73",x"1e"),
   766 => (x"00",x"00",x"07",x"d5"),
   767 => (x"70",x"86",x"c8",x"0f"),
   768 => (x"c5",x"c0",x"05",x"98"),
   769 => (x"c9",x"48",x"c0",x"87"),
   770 => (x"cc",x"27",x"87",x"ec"),
   771 => (x"1e",x"00",x"00",x"16"),
   772 => (x"00",x"00",x"68",x"27"),
   773 => (x"86",x"c4",x"0f",x"00"),
   774 => (x"00",x"17",x"62",x"27"),
   775 => (x"9c",x"27",x"1e",x"00"),
   776 => (x"0f",x"00",x"00",x"00"),
   777 => (x"1e",x"c8",x"86",x"c4"),
   778 => (x"00",x"17",x"7a",x"27"),
   779 => (x"9a",x"27",x"1e",x"00"),
   780 => (x"1e",x"00",x"00",x"18"),
   781 => (x"00",x"0a",x"42",x"27"),
   782 => (x"86",x"cc",x"0f",x"00"),
   783 => (x"c0",x"05",x"98",x"70"),
   784 => (x"08",x"27",x"87",x"cb"),
   785 => (x"48",x"00",x"00",x"18"),
   786 => (x"ef",x"c0",x"78",x"c1"),
   787 => (x"27",x"1e",x"c8",x"87"),
   788 => (x"00",x"00",x"17",x"83"),
   789 => (x"18",x"7e",x"27",x"1e"),
   790 => (x"27",x"1e",x"00",x"00"),
   791 => (x"00",x"00",x"0a",x"42"),
   792 => (x"70",x"86",x"cc",x"0f"),
   793 => (x"d3",x"c0",x"02",x"98"),
   794 => (x"16",x"f3",x"27",x"87"),
   795 => (x"27",x"1e",x"00",x"00"),
   796 => (x"00",x"00",x"00",x"9c"),
   797 => (x"c0",x"86",x"c4",x"0f"),
   798 => (x"87",x"fa",x"c7",x"48"),
   799 => (x"00",x"1a",x"46",x"27"),
   800 => (x"49",x"bf",x"97",x"00"),
   801 => (x"05",x"a9",x"d5",x"c1"),
   802 => (x"27",x"87",x"cf",x"c0"),
   803 => (x"00",x"00",x"1a",x"47"),
   804 => (x"c2",x"49",x"bf",x"97"),
   805 => (x"c0",x"02",x"a9",x"ea"),
   806 => (x"48",x"c0",x"87",x"c5"),
   807 => (x"27",x"87",x"d7",x"c7"),
   808 => (x"00",x"00",x"18",x"48"),
   809 => (x"c3",x"49",x"bf",x"97"),
   810 => (x"c0",x"02",x"a9",x"e9"),
   811 => (x"48",x"27",x"87",x"d4"),
   812 => (x"97",x"00",x"00",x"18"),
   813 => (x"eb",x"c3",x"49",x"bf"),
   814 => (x"c5",x"c0",x"02",x"a9"),
   815 => (x"c6",x"48",x"c0",x"87"),
   816 => (x"53",x"27",x"87",x"f4"),
   817 => (x"97",x"00",x"00",x"18"),
   818 => (x"99",x"71",x"49",x"bf"),
   819 => (x"87",x"ce",x"c0",x"05"),
   820 => (x"00",x"18",x"54",x"27"),
   821 => (x"49",x"bf",x"97",x"00"),
   822 => (x"c0",x"02",x"a9",x"c2"),
   823 => (x"48",x"c0",x"87",x"c5"),
   824 => (x"27",x"87",x"d3",x"c6"),
   825 => (x"00",x"00",x"18",x"55"),
   826 => (x"27",x"48",x"bf",x"97"),
   827 => (x"00",x"00",x"18",x"04"),
   828 => (x"18",x"00",x"27",x"58"),
   829 => (x"49",x"bf",x"00",x"00"),
   830 => (x"8a",x"c1",x"4a",x"71"),
   831 => (x"00",x"18",x"08",x"27"),
   832 => (x"1e",x"72",x"5a",x"00"),
   833 => (x"8c",x"27",x"1e",x"71"),
   834 => (x"1e",x"00",x"00",x"17"),
   835 => (x"00",x"00",x"9c",x"27"),
   836 => (x"86",x"cc",x"0f",x"00"),
   837 => (x"00",x"18",x"56",x"27"),
   838 => (x"49",x"bf",x"97",x"00"),
   839 => (x"57",x"27",x"81",x"73"),
   840 => (x"97",x"00",x"00",x"18"),
   841 => (x"32",x"c8",x"4a",x"bf"),
   842 => (x"80",x"71",x"48",x"72"),
   843 => (x"00",x"18",x"18",x"27"),
   844 => (x"58",x"27",x"58",x"00"),
   845 => (x"97",x"00",x"00",x"18"),
   846 => (x"2c",x"27",x"48",x"bf"),
   847 => (x"58",x"00",x"00",x"18"),
   848 => (x"00",x"18",x"08",x"27"),
   849 => (x"c3",x"02",x"bf",x"00"),
   850 => (x"1e",x"c8",x"87",x"c3"),
   851 => (x"00",x"17",x"10",x"27"),
   852 => (x"9a",x"27",x"1e",x"00"),
   853 => (x"1e",x"00",x"00",x"18"),
   854 => (x"00",x"0a",x"42",x"27"),
   855 => (x"86",x"cc",x"0f",x"00"),
   856 => (x"c0",x"02",x"98",x"70"),
   857 => (x"48",x"c0",x"87",x"c5"),
   858 => (x"27",x"87",x"cb",x"c4"),
   859 => (x"00",x"00",x"18",x"00"),
   860 => (x"48",x"72",x"4a",x"bf"),
   861 => (x"30",x"27",x"30",x"c4"),
   862 => (x"58",x"00",x"00",x"18"),
   863 => (x"00",x"18",x"28",x"27"),
   864 => (x"6d",x"27",x"5a",x"00"),
   865 => (x"97",x"00",x"00",x"18"),
   866 => (x"31",x"c8",x"49",x"bf"),
   867 => (x"00",x"18",x"6c",x"27"),
   868 => (x"4b",x"bf",x"97",x"00"),
   869 => (x"6e",x"27",x"81",x"73"),
   870 => (x"97",x"00",x"00",x"18"),
   871 => (x"33",x"d0",x"4b",x"bf"),
   872 => (x"6f",x"27",x"81",x"73"),
   873 => (x"97",x"00",x"00",x"18"),
   874 => (x"33",x"d8",x"4b",x"bf"),
   875 => (x"34",x"27",x"81",x"73"),
   876 => (x"59",x"00",x"00",x"18"),
   877 => (x"00",x"18",x"28",x"27"),
   878 => (x"27",x"91",x"bf",x"00"),
   879 => (x"00",x"00",x"18",x"14"),
   880 => (x"1c",x"27",x"81",x"bf"),
   881 => (x"59",x"00",x"00",x"18"),
   882 => (x"00",x"18",x"75",x"27"),
   883 => (x"4b",x"bf",x"97",x"00"),
   884 => (x"74",x"27",x"33",x"c8"),
   885 => (x"97",x"00",x"00",x"18"),
   886 => (x"83",x"74",x"4c",x"bf"),
   887 => (x"00",x"18",x"76",x"27"),
   888 => (x"4c",x"bf",x"97",x"00"),
   889 => (x"83",x"74",x"34",x"d0"),
   890 => (x"00",x"18",x"77",x"27"),
   891 => (x"4c",x"bf",x"97",x"00"),
   892 => (x"34",x"d8",x"9c",x"cf"),
   893 => (x"20",x"27",x"83",x"74"),
   894 => (x"5b",x"00",x"00",x"18"),
   895 => (x"92",x"73",x"8b",x"c2"),
   896 => (x"80",x"71",x"48",x"72"),
   897 => (x"00",x"18",x"24",x"27"),
   898 => (x"e7",x"c1",x"58",x"00"),
   899 => (x"18",x"5a",x"27",x"87"),
   900 => (x"bf",x"97",x"00",x"00"),
   901 => (x"27",x"31",x"c8",x"49"),
   902 => (x"00",x"00",x"18",x"59"),
   903 => (x"72",x"4a",x"bf",x"97"),
   904 => (x"18",x"30",x"27",x"81"),
   905 => (x"c5",x"59",x"00",x"00"),
   906 => (x"81",x"ff",x"c7",x"31"),
   907 => (x"28",x"27",x"29",x"c9"),
   908 => (x"59",x"00",x"00",x"18"),
   909 => (x"00",x"18",x"5f",x"27"),
   910 => (x"4a",x"bf",x"97",x"00"),
   911 => (x"5e",x"27",x"32",x"c8"),
   912 => (x"97",x"00",x"00",x"18"),
   913 => (x"82",x"73",x"4b",x"bf"),
   914 => (x"00",x"18",x"34",x"27"),
   915 => (x"28",x"27",x"5a",x"00"),
   916 => (x"bf",x"00",x"00",x"18"),
   917 => (x"18",x"14",x"27",x"92"),
   918 => (x"82",x"bf",x"00",x"00"),
   919 => (x"00",x"18",x"24",x"27"),
   920 => (x"1c",x"27",x"5a",x"00"),
   921 => (x"48",x"00",x"00",x"18"),
   922 => (x"48",x"72",x"78",x"c0"),
   923 => (x"1c",x"27",x"80",x"71"),
   924 => (x"58",x"00",x"00",x"18"),
   925 => (x"f0",x"ff",x"48",x"c1"),
   926 => (x"5e",x"0e",x"87",x"d6"),
   927 => (x"27",x"0e",x"5c",x"5b"),
   928 => (x"00",x"00",x"18",x"08"),
   929 => (x"cf",x"c0",x"02",x"bf"),
   930 => (x"4a",x"66",x"cc",x"87"),
   931 => (x"cc",x"2a",x"b7",x"c7"),
   932 => (x"ff",x"c1",x"4b",x"66"),
   933 => (x"87",x"cc",x"c0",x"9b"),
   934 => (x"c8",x"4a",x"66",x"cc"),
   935 => (x"66",x"cc",x"2a",x"b7"),
   936 => (x"9b",x"ff",x"c3",x"4b"),
   937 => (x"00",x"18",x"48",x"27"),
   938 => (x"14",x"27",x"1e",x"00"),
   939 => (x"bf",x"00",x"00",x"18"),
   940 => (x"71",x"81",x"72",x"49"),
   941 => (x"07",x"d5",x"27",x"1e"),
   942 => (x"c8",x"0f",x"00",x"00"),
   943 => (x"05",x"98",x"70",x"86"),
   944 => (x"c0",x"87",x"c5",x"c0"),
   945 => (x"87",x"f0",x"c0",x"48"),
   946 => (x"00",x"18",x"08",x"27"),
   947 => (x"c0",x"02",x"bf",x"00"),
   948 => (x"49",x"73",x"87",x"d6"),
   949 => (x"27",x"91",x"b7",x"c4"),
   950 => (x"00",x"00",x"18",x"48"),
   951 => (x"cf",x"4c",x"69",x"81"),
   952 => (x"ff",x"ff",x"ff",x"ff"),
   953 => (x"87",x"ce",x"c0",x"9c"),
   954 => (x"b7",x"c2",x"49",x"73"),
   955 => (x"18",x"48",x"27",x"91"),
   956 => (x"9f",x"81",x"00",x"00"),
   957 => (x"48",x"74",x"4c",x"69"),
   958 => (x"87",x"d6",x"ee",x"ff"),
   959 => (x"5c",x"5b",x"5e",x"0e"),
   960 => (x"86",x"f4",x"0e",x"5d"),
   961 => (x"48",x"76",x"4b",x"c0"),
   962 => (x"00",x"18",x"1c",x"27"),
   963 => (x"c4",x"78",x"bf",x"00"),
   964 => (x"20",x"27",x"48",x"a6"),
   965 => (x"bf",x"00",x"00",x"18"),
   966 => (x"18",x"08",x"27",x"78"),
   967 => (x"02",x"bf",x"00",x"00"),
   968 => (x"27",x"87",x"cc",x"c0"),
   969 => (x"00",x"00",x"18",x"00"),
   970 => (x"31",x"c4",x"49",x"bf"),
   971 => (x"27",x"87",x"c9",x"c0"),
   972 => (x"00",x"00",x"18",x"24"),
   973 => (x"31",x"c4",x"49",x"bf"),
   974 => (x"c0",x"59",x"a6",x"cc"),
   975 => (x"48",x"66",x"c8",x"4d"),
   976 => (x"c3",x"06",x"a8",x"c0"),
   977 => (x"49",x"75",x"87",x"c2"),
   978 => (x"99",x"71",x"99",x"cf"),
   979 => (x"87",x"e2",x"c0",x"05"),
   980 => (x"00",x"18",x"48",x"27"),
   981 => (x"66",x"c8",x"1e",x"00"),
   982 => (x"80",x"c1",x"48",x"49"),
   983 => (x"71",x"58",x"a6",x"cc"),
   984 => (x"07",x"d5",x"27",x"1e"),
   985 => (x"c8",x"0f",x"00",x"00"),
   986 => (x"18",x"48",x"27",x"86"),
   987 => (x"c0",x"4b",x"00",x"00"),
   988 => (x"e0",x"c0",x"87",x"c3"),
   989 => (x"49",x"6b",x"97",x"83"),
   990 => (x"c2",x"02",x"99",x"71"),
   991 => (x"6b",x"97",x"87",x"c1"),
   992 => (x"a9",x"e5",x"c3",x"49"),
   993 => (x"87",x"f7",x"c1",x"02"),
   994 => (x"81",x"cb",x"49",x"73"),
   995 => (x"d8",x"49",x"69",x"97"),
   996 => (x"05",x"99",x"71",x"99"),
   997 => (x"73",x"87",x"e8",x"c1"),
   998 => (x"00",x"68",x"27",x"1e"),
   999 => (x"c4",x"0f",x"00",x"00"),
  1000 => (x"c0",x"1e",x"cb",x"86"),
  1001 => (x"73",x"1e",x"66",x"e4"),
  1002 => (x"0a",x"42",x"27",x"1e"),
  1003 => (x"cc",x"0f",x"00",x"00"),
  1004 => (x"05",x"98",x"70",x"86"),
  1005 => (x"73",x"87",x"c8",x"c1"),
  1006 => (x"66",x"82",x"dc",x"4a"),
  1007 => (x"6a",x"81",x"c4",x"49"),
  1008 => (x"da",x"4a",x"73",x"79"),
  1009 => (x"49",x"66",x"dc",x"82"),
  1010 => (x"6a",x"9f",x"81",x"c8"),
  1011 => (x"71",x"79",x"70",x"48"),
  1012 => (x"18",x"08",x"27",x"4c"),
  1013 => (x"02",x"bf",x"00",x"00"),
  1014 => (x"73",x"87",x"d2",x"c0"),
  1015 => (x"9f",x"81",x"d4",x"49"),
  1016 => (x"ff",x"c0",x"49",x"69"),
  1017 => (x"4a",x"71",x"99",x"ff"),
  1018 => (x"c2",x"c0",x"32",x"d0"),
  1019 => (x"72",x"4a",x"c0",x"87"),
  1020 => (x"70",x"80",x"6c",x"48"),
  1021 => (x"48",x"66",x"dc",x"7c"),
  1022 => (x"48",x"c1",x"78",x"c0"),
  1023 => (x"c1",x"87",x"c9",x"c1"),
  1024 => (x"ad",x"66",x"c8",x"85"),
  1025 => (x"87",x"fe",x"fc",x"04"),
  1026 => (x"00",x"18",x"08",x"27"),
  1027 => (x"c0",x"02",x"bf",x"00"),
  1028 => (x"1e",x"6e",x"87",x"f4"),
  1029 => (x"00",x"0e",x"7a",x"27"),
  1030 => (x"86",x"c4",x"0f",x"00"),
  1031 => (x"6e",x"58",x"a6",x"c4"),
  1032 => (x"ff",x"ff",x"cf",x"49"),
  1033 => (x"a9",x"99",x"f8",x"ff"),
  1034 => (x"87",x"da",x"c0",x"02"),
  1035 => (x"89",x"c2",x"49",x"6e"),
  1036 => (x"00",x"18",x"00",x"27"),
  1037 => (x"27",x"91",x"bf",x"00"),
  1038 => (x"00",x"00",x"18",x"18"),
  1039 => (x"80",x"71",x"48",x"bf"),
  1040 => (x"fb",x"58",x"a6",x"c8"),
  1041 => (x"48",x"c0",x"87",x"f5"),
  1042 => (x"e9",x"ff",x"8e",x"f4"),
  1043 => (x"73",x"1e",x"87",x"c2"),
  1044 => (x"bf",x"66",x"c8",x"1e"),
  1045 => (x"c8",x"81",x"c1",x"49"),
  1046 => (x"09",x"79",x"09",x"66"),
  1047 => (x"00",x"18",x"04",x"27"),
  1048 => (x"71",x"99",x"bf",x"00"),
  1049 => (x"d2",x"c0",x"05",x"99"),
  1050 => (x"4b",x"66",x"c8",x"87"),
  1051 => (x"1e",x"6b",x"83",x"c8"),
  1052 => (x"00",x"0e",x"7a",x"27"),
  1053 => (x"86",x"c4",x"0f",x"00"),
  1054 => (x"c1",x"7b",x"49",x"70"),
  1055 => (x"d3",x"e8",x"ff",x"48"),
  1056 => (x"18",x"27",x"1e",x"87"),
  1057 => (x"bf",x"00",x"00",x"18"),
  1058 => (x"4a",x"66",x"c4",x"49"),
  1059 => (x"4a",x"6a",x"82",x"c8"),
  1060 => (x"00",x"27",x"8a",x"c2"),
  1061 => (x"bf",x"00",x"00",x"18"),
  1062 => (x"27",x"81",x"72",x"92"),
  1063 => (x"00",x"00",x"18",x"04"),
  1064 => (x"66",x"c4",x"4a",x"bf"),
  1065 => (x"81",x"72",x"9a",x"bf"),
  1066 => (x"71",x"1e",x"66",x"c8"),
  1067 => (x"07",x"d5",x"27",x"1e"),
  1068 => (x"c8",x"0f",x"00",x"00"),
  1069 => (x"05",x"98",x"70",x"86"),
  1070 => (x"c0",x"87",x"c5",x"c0"),
  1071 => (x"87",x"c2",x"c0",x"48"),
  1072 => (x"e7",x"ff",x"48",x"c1"),
  1073 => (x"5e",x"0e",x"87",x"d0"),
  1074 => (x"cc",x"0e",x"5c",x"5b"),
  1075 => (x"38",x"27",x"1e",x"66"),
  1076 => (x"1e",x"00",x"00",x"18"),
  1077 => (x"00",x"0e",x"fc",x"27"),
  1078 => (x"86",x"c8",x"0f",x"00"),
  1079 => (x"c1",x"02",x"98",x"70"),
  1080 => (x"3c",x"27",x"87",x"e4"),
  1081 => (x"bf",x"00",x"00",x"18"),
  1082 => (x"81",x"ff",x"c7",x"49"),
  1083 => (x"4c",x"71",x"29",x"c9"),
  1084 => (x"62",x"27",x"4b",x"c0"),
  1085 => (x"1e",x"00",x"00",x"11"),
  1086 => (x"00",x"00",x"68",x"27"),
  1087 => (x"86",x"c4",x"0f",x"00"),
  1088 => (x"06",x"ac",x"b7",x"c0"),
  1089 => (x"d0",x"87",x"d5",x"c1"),
  1090 => (x"38",x"27",x"1e",x"66"),
  1091 => (x"1e",x"00",x"00",x"18"),
  1092 => (x"00",x"10",x"81",x"27"),
  1093 => (x"86",x"c8",x"0f",x"00"),
  1094 => (x"c0",x"05",x"98",x"70"),
  1095 => (x"48",x"c0",x"87",x"c5"),
  1096 => (x"27",x"87",x"fb",x"c0"),
  1097 => (x"00",x"00",x"18",x"38"),
  1098 => (x"10",x"4e",x"27",x"1e"),
  1099 => (x"c4",x"0f",x"00",x"00"),
  1100 => (x"48",x"66",x"d0",x"86"),
  1101 => (x"d4",x"80",x"c0",x"c8"),
  1102 => (x"83",x"c1",x"58",x"a6"),
  1103 => (x"04",x"ab",x"b7",x"74"),
  1104 => (x"c0",x"87",x"c4",x"ff"),
  1105 => (x"66",x"cc",x"87",x"d6"),
  1106 => (x"11",x"7b",x"27",x"1e"),
  1107 => (x"27",x"1e",x"00",x"00"),
  1108 => (x"00",x"00",x"00",x"9c"),
  1109 => (x"c0",x"86",x"c8",x"0f"),
  1110 => (x"87",x"c2",x"c0",x"48"),
  1111 => (x"e4",x"ff",x"48",x"c1"),
  1112 => (x"70",x"4f",x"87",x"f0"),
  1113 => (x"64",x"65",x"6e",x"65"),
  1114 => (x"6c",x"69",x"66",x"20"),
  1115 => (x"6c",x"20",x"2c",x"65"),
  1116 => (x"69",x"64",x"61",x"6f"),
  1117 => (x"2e",x"2e",x"67",x"6e"),
  1118 => (x"43",x"00",x"0a",x"2e"),
  1119 => (x"74",x"27",x"6e",x"61"),
  1120 => (x"65",x"70",x"6f",x"20"),
  1121 => (x"73",x"25",x"20",x"6e"),
  1122 => (x"c4",x"1e",x"00",x"0a"),
  1123 => (x"29",x"d8",x"49",x"66"),
  1124 => (x"c4",x"99",x"ff",x"c3"),
  1125 => (x"2a",x"c8",x"4a",x"66"),
  1126 => (x"9a",x"c0",x"fc",x"cf"),
  1127 => (x"66",x"c4",x"b1",x"72"),
  1128 => (x"c0",x"32",x"c8",x"4a"),
  1129 => (x"c0",x"c0",x"f0",x"ff"),
  1130 => (x"c4",x"b1",x"72",x"9a"),
  1131 => (x"32",x"d8",x"4a",x"66"),
  1132 => (x"c0",x"c0",x"c0",x"ff"),
  1133 => (x"b1",x"72",x"9a",x"c0"),
  1134 => (x"c0",x"c0",x"48",x"71"),
  1135 => (x"4d",x"26",x"87",x"c6"),
  1136 => (x"4b",x"26",x"4c",x"26"),
  1137 => (x"c4",x"1e",x"4f",x"26"),
  1138 => (x"2a",x"c8",x"4a",x"66"),
  1139 => (x"cf",x"9a",x"ff",x"c3"),
  1140 => (x"c4",x"9a",x"ff",x"ff"),
  1141 => (x"31",x"c8",x"49",x"66"),
  1142 => (x"99",x"c0",x"fc",x"cf"),
  1143 => (x"ff",x"cf",x"b1",x"72"),
  1144 => (x"48",x"71",x"99",x"ff"),
  1145 => (x"87",x"dc",x"ff",x"ff"),
  1146 => (x"49",x"66",x"c4",x"1e"),
  1147 => (x"ff",x"cf",x"29",x"d0"),
  1148 => (x"66",x"c4",x"99",x"ff"),
  1149 => (x"f0",x"32",x"d0",x"4a"),
  1150 => (x"72",x"9a",x"c0",x"c0"),
  1151 => (x"ff",x"48",x"71",x"b1"),
  1152 => (x"1e",x"87",x"c1",x"ff"),
  1153 => (x"c0",x"d0",x"1e",x"73"),
  1154 => (x"4b",x"c0",x"c0",x"c0"),
  1155 => (x"fd",x"ff",x"0f",x"73"),
  1156 => (x"c4",x"c0",x"c0",x"87"),
  1157 => (x"26",x"4d",x"26",x"87"),
  1158 => (x"26",x"4b",x"26",x"4c"),
  1159 => (x"66",x"c8",x"1e",x"4f"),
  1160 => (x"99",x"df",x"c3",x"49"),
  1161 => (x"c0",x"89",x"f7",x"c0"),
  1162 => (x"c0",x"03",x"a9",x"b7"),
  1163 => (x"e7",x"c0",x"87",x"c3"),
  1164 => (x"48",x"66",x"c4",x"81"),
  1165 => (x"a6",x"c8",x"30",x"c4"),
  1166 => (x"48",x"66",x"c4",x"58"),
  1167 => (x"a6",x"c8",x"b0",x"71"),
  1168 => (x"48",x"66",x"c4",x"58"),
  1169 => (x"87",x"d3",x"ff",x"ff"),
  1170 => (x"5c",x"5b",x"5e",x"0e"),
  1171 => (x"c0",x"c0",x"d0",x"0e"),
  1172 => (x"27",x"4c",x"c0",x"c0"),
  1173 => (x"00",x"00",x"1a",x"48"),
  1174 => (x"80",x"c1",x"48",x"bf"),
  1175 => (x"00",x"1a",x"4c",x"27"),
  1176 => (x"cc",x"97",x"58",x"00"),
  1177 => (x"c0",x"fe",x"49",x"66"),
  1178 => (x"d3",x"c1",x"b9",x"81"),
  1179 => (x"e9",x"c0",x"05",x"a9"),
  1180 => (x"1a",x"48",x"27",x"87"),
  1181 => (x"c0",x"48",x"00",x"00"),
  1182 => (x"1a",x"4c",x"27",x"78"),
  1183 => (x"c0",x"48",x"00",x"00"),
  1184 => (x"1a",x"54",x"27",x"78"),
  1185 => (x"c0",x"48",x"00",x"00"),
  1186 => (x"1a",x"58",x"27",x"78"),
  1187 => (x"c0",x"48",x"00",x"00"),
  1188 => (x"48",x"c0",x"ff",x"78"),
  1189 => (x"c9",x"78",x"d3",x"c1"),
  1190 => (x"48",x"27",x"87",x"e3"),
  1191 => (x"bf",x"00",x"00",x"1a"),
  1192 => (x"05",x"a8",x"c1",x"48"),
  1193 => (x"ff",x"87",x"d4",x"c1"),
  1194 => (x"f4",x"c1",x"48",x"c0"),
  1195 => (x"66",x"cc",x"97",x"78"),
  1196 => (x"81",x"c0",x"fe",x"49"),
  1197 => (x"27",x"1e",x"71",x"b9"),
  1198 => (x"00",x"00",x"1a",x"58"),
  1199 => (x"1d",x"27",x"1e",x"bf"),
  1200 => (x"0f",x"00",x"00",x"12"),
  1201 => (x"5c",x"27",x"86",x"c8"),
  1202 => (x"58",x"00",x"00",x"1a"),
  1203 => (x"00",x"1a",x"58",x"27"),
  1204 => (x"c3",x"4a",x"bf",x"00"),
  1205 => (x"c0",x"06",x"aa",x"b7"),
  1206 => (x"48",x"ca",x"87",x"c6"),
  1207 => (x"4a",x"70",x"88",x"72"),
  1208 => (x"81",x"c1",x"49",x"72"),
  1209 => (x"30",x"c1",x"48",x"71"),
  1210 => (x"00",x"1a",x"54",x"27"),
  1211 => (x"48",x"72",x"58",x"00"),
  1212 => (x"ff",x"80",x"f0",x"c0"),
  1213 => (x"08",x"78",x"08",x"c0"),
  1214 => (x"27",x"87",x"c2",x"c8"),
  1215 => (x"00",x"00",x"1a",x"58"),
  1216 => (x"b7",x"c9",x"48",x"bf"),
  1217 => (x"f4",x"c7",x"01",x"a8"),
  1218 => (x"1a",x"58",x"27",x"87"),
  1219 => (x"48",x"bf",x"00",x"00"),
  1220 => (x"06",x"a8",x"b7",x"c0"),
  1221 => (x"27",x"87",x"e6",x"c7"),
  1222 => (x"00",x"00",x"1a",x"58"),
  1223 => (x"f0",x"c0",x"48",x"bf"),
  1224 => (x"08",x"c0",x"ff",x"80"),
  1225 => (x"48",x"27",x"08",x"78"),
  1226 => (x"bf",x"00",x"00",x"1a"),
  1227 => (x"a8",x"b7",x"c3",x"48"),
  1228 => (x"87",x"e2",x"c0",x"01"),
  1229 => (x"49",x"66",x"cc",x"97"),
  1230 => (x"b9",x"81",x"c0",x"fe"),
  1231 => (x"54",x"27",x"1e",x"71"),
  1232 => (x"bf",x"00",x"00",x"1a"),
  1233 => (x"12",x"1d",x"27",x"1e"),
  1234 => (x"c8",x"0f",x"00",x"00"),
  1235 => (x"1a",x"58",x"27",x"86"),
  1236 => (x"c6",x"58",x"00",x"00"),
  1237 => (x"50",x"27",x"87",x"e7"),
  1238 => (x"bf",x"00",x"00",x"1a"),
  1239 => (x"27",x"81",x"c3",x"49"),
  1240 => (x"00",x"00",x"1a",x"48"),
  1241 => (x"04",x"a9",x"b7",x"bf"),
  1242 => (x"97",x"87",x"ea",x"c0"),
  1243 => (x"fe",x"49",x"66",x"cc"),
  1244 => (x"71",x"b9",x"81",x"c0"),
  1245 => (x"1a",x"4c",x"27",x"1e"),
  1246 => (x"1e",x"bf",x"00",x"00"),
  1247 => (x"00",x"12",x"1d",x"27"),
  1248 => (x"86",x"c8",x"0f",x"00"),
  1249 => (x"00",x"1a",x"50",x"27"),
  1250 => (x"5c",x"27",x"58",x"00"),
  1251 => (x"48",x"00",x"00",x"1a"),
  1252 => (x"e8",x"c5",x"78",x"c1"),
  1253 => (x"1a",x"58",x"27",x"87"),
  1254 => (x"48",x"bf",x"00",x"00"),
  1255 => (x"06",x"a8",x"b7",x"c0"),
  1256 => (x"27",x"87",x"c4",x"c3"),
  1257 => (x"00",x"00",x"1a",x"58"),
  1258 => (x"b7",x"c3",x"48",x"bf"),
  1259 => (x"f6",x"c2",x"01",x"a8"),
  1260 => (x"1a",x"54",x"27",x"87"),
  1261 => (x"49",x"bf",x"00",x"00"),
  1262 => (x"27",x"81",x"31",x"c1"),
  1263 => (x"00",x"00",x"1a",x"48"),
  1264 => (x"04",x"a9",x"b7",x"bf"),
  1265 => (x"97",x"87",x"fa",x"c1"),
  1266 => (x"fe",x"49",x"66",x"cc"),
  1267 => (x"71",x"b9",x"81",x"c0"),
  1268 => (x"1a",x"60",x"27",x"1e"),
  1269 => (x"1e",x"bf",x"00",x"00"),
  1270 => (x"00",x"12",x"1d",x"27"),
  1271 => (x"86",x"c8",x"0f",x"00"),
  1272 => (x"00",x"1a",x"64",x"27"),
  1273 => (x"5c",x"27",x"58",x"00"),
  1274 => (x"bf",x"00",x"00",x"1a"),
  1275 => (x"27",x"89",x"c1",x"49"),
  1276 => (x"00",x"00",x"1a",x"60"),
  1277 => (x"a9",x"b7",x"c0",x"59"),
  1278 => (x"87",x"c1",x"c4",x"03"),
  1279 => (x"00",x"1a",x"4c",x"27"),
  1280 => (x"27",x"49",x"bf",x"00"),
  1281 => (x"00",x"00",x"1a",x"60"),
  1282 => (x"c3",x"51",x"bf",x"97"),
  1283 => (x"4c",x"27",x"98",x"ff"),
  1284 => (x"bf",x"00",x"00",x"1a"),
  1285 => (x"27",x"81",x"c1",x"49"),
  1286 => (x"00",x"00",x"1a",x"50"),
  1287 => (x"1a",x"64",x"27",x"59"),
  1288 => (x"b7",x"bf",x"00",x"00"),
  1289 => (x"cd",x"c0",x"06",x"a9"),
  1290 => (x"1a",x"64",x"27",x"87"),
  1291 => (x"27",x"48",x"00",x"00"),
  1292 => (x"00",x"00",x"1a",x"4c"),
  1293 => (x"5c",x"27",x"78",x"bf"),
  1294 => (x"48",x"00",x"00",x"1a"),
  1295 => (x"fc",x"c2",x"78",x"c1"),
  1296 => (x"1a",x"5c",x"27",x"87"),
  1297 => (x"05",x"bf",x"00",x"00"),
  1298 => (x"27",x"87",x"f2",x"c2"),
  1299 => (x"00",x"00",x"1a",x"60"),
  1300 => (x"31",x"c4",x"49",x"bf"),
  1301 => (x"00",x"1a",x"64",x"27"),
  1302 => (x"4c",x"27",x"59",x"00"),
  1303 => (x"bf",x"00",x"00",x"1a"),
  1304 => (x"09",x"79",x"97",x"09"),
  1305 => (x"27",x"87",x"d6",x"c2"),
  1306 => (x"00",x"00",x"1a",x"58"),
  1307 => (x"b7",x"c7",x"48",x"bf"),
  1308 => (x"f9",x"c1",x"04",x"a8"),
  1309 => (x"fe",x"4b",x"c0",x"87"),
  1310 => (x"78",x"c1",x"48",x"f4"),
  1311 => (x"00",x"1a",x"64",x"27"),
  1312 => (x"74",x"1e",x"bf",x"00"),
  1313 => (x"17",x"b0",x"27",x"1e"),
  1314 => (x"27",x"1e",x"00",x"00"),
  1315 => (x"00",x"00",x"00",x"9c"),
  1316 => (x"27",x"86",x"cc",x"0f"),
  1317 => (x"00",x"00",x"1a",x"50"),
  1318 => (x"1a",x"4c",x"27",x"5c"),
  1319 => (x"48",x"bf",x"00",x"00"),
  1320 => (x"00",x"1a",x"64",x"27"),
  1321 => (x"a8",x"b7",x"bf",x"00"),
  1322 => (x"87",x"e3",x"c0",x"03"),
  1323 => (x"00",x"1a",x"4c",x"27"),
  1324 => (x"83",x"bf",x"bf",x"00"),
  1325 => (x"00",x"1a",x"4c",x"27"),
  1326 => (x"c4",x"49",x"bf",x"00"),
  1327 => (x"1a",x"50",x"27",x"81"),
  1328 => (x"27",x"59",x"00",x"00"),
  1329 => (x"00",x"00",x"1a",x"64"),
  1330 => (x"04",x"a9",x"b7",x"bf"),
  1331 => (x"73",x"87",x"dd",x"ff"),
  1332 => (x"17",x"cf",x"27",x"1e"),
  1333 => (x"27",x"1e",x"00",x"00"),
  1334 => (x"00",x"00",x"00",x"9c"),
  1335 => (x"ff",x"86",x"c8",x"0f"),
  1336 => (x"c2",x"c1",x"48",x"c0"),
  1337 => (x"12",x"03",x"27",x"78"),
  1338 => (x"c0",x"0f",x"00",x"00"),
  1339 => (x"58",x"27",x"87",x"cf"),
  1340 => (x"bf",x"00",x"00",x"1a"),
  1341 => (x"80",x"f0",x"c0",x"48"),
  1342 => (x"78",x"08",x"c0",x"ff"),
  1343 => (x"d6",x"f4",x"ff",x"08"),
  1344 => (x"5b",x"5e",x"0e",x"87"),
  1345 => (x"27",x"0e",x"5d",x"5c"),
  1346 => (x"00",x"00",x"16",x"03"),
  1347 => (x"00",x"68",x"27",x"1e"),
  1348 => (x"c4",x"0f",x"00",x"00"),
  1349 => (x"04",x"de",x"27",x"86"),
  1350 => (x"70",x"0f",x"00",x"00"),
  1351 => (x"d1",x"c0",x"02",x"98"),
  1352 => (x"0a",x"98",x"27",x"87"),
  1353 => (x"70",x"0f",x"00",x"00"),
  1354 => (x"c5",x"c0",x"02",x"98"),
  1355 => (x"c0",x"49",x"c1",x"87"),
  1356 => (x"49",x"c0",x"87",x"c2"),
  1357 => (x"19",x"27",x"4d",x"71"),
  1358 => (x"1e",x"00",x"00",x"16"),
  1359 => (x"00",x"00",x"68",x"27"),
  1360 => (x"86",x"c4",x"0f",x"00"),
  1361 => (x"00",x"1a",x"64",x"27"),
  1362 => (x"78",x"c0",x"48",x"00"),
  1363 => (x"27",x"1e",x"ee",x"c0"),
  1364 => (x"00",x"00",x"00",x"45"),
  1365 => (x"c3",x"86",x"c4",x"0f"),
  1366 => (x"4a",x"ff",x"c8",x"f4"),
  1367 => (x"4c",x"bf",x"c0",x"ff"),
  1368 => (x"c0",x"c8",x"49",x"74"),
  1369 => (x"02",x"99",x"71",x"99"),
  1370 => (x"74",x"87",x"df",x"c1"),
  1371 => (x"9b",x"ff",x"c3",x"4b"),
  1372 => (x"c1",x"05",x"ab",x"db"),
  1373 => (x"9d",x"75",x"87",x"c5"),
  1374 => (x"87",x"f1",x"c0",x"02"),
  1375 => (x"c0",x"c0",x"c0",x"d0"),
  1376 => (x"e7",x"27",x"1e",x"c0"),
  1377 => (x"1e",x"00",x"00",x"15"),
  1378 => (x"00",x"10",x"c6",x"27"),
  1379 => (x"86",x"c8",x"0f",x"00"),
  1380 => (x"c0",x"02",x"98",x"70"),
  1381 => (x"db",x"27",x"87",x"d7"),
  1382 => (x"1e",x"00",x"00",x"15"),
  1383 => (x"00",x"00",x"68",x"27"),
  1384 => (x"86",x"c4",x"0f",x"00"),
  1385 => (x"00",x"12",x"03",x"27"),
  1386 => (x"ce",x"c0",x"0f",x"00"),
  1387 => (x"15",x"f3",x"27",x"87"),
  1388 => (x"27",x"1e",x"00",x"00"),
  1389 => (x"00",x"00",x"00",x"68"),
  1390 => (x"73",x"86",x"c4",x"0f"),
  1391 => (x"12",x"48",x"27",x"1e"),
  1392 => (x"c4",x"0f",x"00",x"00"),
  1393 => (x"c9",x"f4",x"c3",x"86"),
  1394 => (x"49",x"72",x"4a",x"c0"),
  1395 => (x"99",x"71",x"8a",x"c1"),
  1396 => (x"87",x"c8",x"fe",x"05"),
  1397 => (x"ff",x"87",x"f5",x"fd"),
  1398 => (x"42",x"87",x"fa",x"f0"),
  1399 => (x"69",x"74",x"6f",x"6f"),
  1400 => (x"2e",x"2e",x"67",x"6e"),
  1401 => (x"42",x"00",x"0a",x"2e"),
  1402 => (x"38",x"54",x"4f",x"4f"),
  1403 => (x"42",x"20",x"32",x"33"),
  1404 => (x"53",x"00",x"4e",x"49"),
  1405 => (x"6f",x"62",x"20",x"44"),
  1406 => (x"66",x"20",x"74",x"6f"),
  1407 => (x"65",x"6c",x"69",x"61"),
  1408 => (x"49",x"00",x"0a",x"64"),
  1409 => (x"69",x"74",x"69",x"6e"),
  1410 => (x"7a",x"69",x"6c",x"61"),
  1411 => (x"20",x"67",x"6e",x"69"),
  1412 => (x"63",x"20",x"44",x"53"),
  1413 => (x"0a",x"64",x"72",x"61"),
  1414 => (x"32",x"53",x"52",x"00"),
  1415 => (x"62",x"20",x"32",x"33"),
  1416 => (x"20",x"74",x"6f",x"6f"),
  1417 => (x"72",x"70",x"20",x"2d"),
  1418 => (x"20",x"73",x"73",x"65"),
  1419 => (x"20",x"43",x"53",x"45"),
  1420 => (x"62",x"20",x"6f",x"74"),
  1421 => (x"20",x"74",x"6f",x"6f"),
  1422 => (x"6d",x"6f",x"72",x"66"),
  1423 => (x"2e",x"44",x"53",x"20"),
  1424 => (x"44",x"4d",x"43",x"00"),
  1425 => (x"61",x"65",x"52",x"00"),
  1426 => (x"66",x"6f",x"20",x"64"),
  1427 => (x"52",x"42",x"4d",x"20"),
  1428 => (x"69",x"61",x"66",x"20"),
  1429 => (x"0a",x"64",x"65",x"6c"),
  1430 => (x"20",x"6f",x"4e",x"00"),
  1431 => (x"74",x"72",x"61",x"70"),
  1432 => (x"6f",x"69",x"74",x"69"),
  1433 => (x"69",x"73",x"20",x"6e"),
  1434 => (x"74",x"61",x"6e",x"67"),
  1435 => (x"20",x"65",x"72",x"75"),
  1436 => (x"6e",x"75",x"6f",x"66"),
  1437 => (x"4d",x"00",x"0a",x"64"),
  1438 => (x"69",x"73",x"52",x"42"),
  1439 => (x"20",x"3a",x"65",x"7a"),
  1440 => (x"20",x"2c",x"64",x"25"),
  1441 => (x"74",x"72",x"61",x"70"),
  1442 => (x"6f",x"69",x"74",x"69"),
  1443 => (x"7a",x"69",x"73",x"6e"),
  1444 => (x"25",x"20",x"3a",x"65"),
  1445 => (x"6f",x"20",x"2c",x"64"),
  1446 => (x"65",x"73",x"66",x"66"),
  1447 => (x"66",x"6f",x"20",x"74"),
  1448 => (x"67",x"69",x"73",x"20"),
  1449 => (x"64",x"25",x"20",x"3a"),
  1450 => (x"69",x"73",x"20",x"2c"),
  1451 => (x"78",x"30",x"20",x"67"),
  1452 => (x"00",x"0a",x"78",x"25"),
  1453 => (x"64",x"61",x"65",x"52"),
  1454 => (x"20",x"67",x"6e",x"69"),
  1455 => (x"74",x"6f",x"6f",x"62"),
  1456 => (x"63",x"65",x"73",x"20"),
  1457 => (x"20",x"72",x"6f",x"74"),
  1458 => (x"00",x"0a",x"64",x"25"),
  1459 => (x"64",x"61",x"65",x"52"),
  1460 => (x"6f",x"6f",x"62",x"20"),
  1461 => (x"65",x"73",x"20",x"74"),
  1462 => (x"72",x"6f",x"74",x"63"),
  1463 => (x"6f",x"72",x"66",x"20"),
  1464 => (x"69",x"66",x"20",x"6d"),
  1465 => (x"20",x"74",x"73",x"72"),
  1466 => (x"74",x"72",x"61",x"70"),
  1467 => (x"6f",x"69",x"74",x"69"),
  1468 => (x"55",x"00",x"0a",x"6e"),
  1469 => (x"70",x"75",x"73",x"6e"),
  1470 => (x"74",x"72",x"6f",x"70"),
  1471 => (x"70",x"20",x"64",x"65"),
  1472 => (x"69",x"74",x"72",x"61"),
  1473 => (x"6e",x"6f",x"69",x"74"),
  1474 => (x"70",x"79",x"74",x"20"),
  1475 => (x"00",x"0d",x"21",x"65"),
  1476 => (x"33",x"54",x"41",x"46"),
  1477 => (x"20",x"20",x"20",x"32"),
  1478 => (x"61",x"65",x"52",x"00"),
  1479 => (x"67",x"6e",x"69",x"64"),
  1480 => (x"52",x"42",x"4d",x"20"),
  1481 => (x"42",x"4d",x"00",x"0a"),
  1482 => (x"75",x"73",x"20",x"52"),
  1483 => (x"73",x"65",x"63",x"63"),
  1484 => (x"6c",x"75",x"66",x"73"),
  1485 => (x"72",x"20",x"79",x"6c"),
  1486 => (x"0a",x"64",x"61",x"65"),
  1487 => (x"54",x"41",x"46",x"00"),
  1488 => (x"20",x"20",x"36",x"31"),
  1489 => (x"41",x"46",x"00",x"20"),
  1490 => (x"20",x"32",x"33",x"54"),
  1491 => (x"50",x"00",x"20",x"20"),
  1492 => (x"69",x"74",x"72",x"61"),
  1493 => (x"6e",x"6f",x"69",x"74"),
  1494 => (x"6e",x"75",x"6f",x"63"),
  1495 => (x"64",x"25",x"20",x"74"),
  1496 => (x"75",x"48",x"00",x"0a"),
  1497 => (x"6e",x"69",x"74",x"6e"),
  1498 => (x"6f",x"66",x"20",x"67"),
  1499 => (x"69",x"66",x"20",x"72"),
  1500 => (x"79",x"73",x"65",x"6c"),
  1501 => (x"6d",x"65",x"74",x"73"),
  1502 => (x"41",x"46",x"00",x"0a"),
  1503 => (x"20",x"32",x"33",x"54"),
  1504 => (x"46",x"00",x"20",x"20"),
  1505 => (x"36",x"31",x"54",x"41"),
  1506 => (x"00",x"20",x"20",x"20"),
  1507 => (x"73",x"75",x"6c",x"43"),
  1508 => (x"20",x"72",x"65",x"74"),
  1509 => (x"65",x"7a",x"69",x"73"),
  1510 => (x"64",x"25",x"20",x"3a"),
  1511 => (x"6c",x"43",x"20",x"2c"),
  1512 => (x"65",x"74",x"73",x"75"),
  1513 => (x"61",x"6d",x"20",x"72"),
  1514 => (x"20",x"2c",x"6b",x"73"),
  1515 => (x"00",x"0a",x"64",x"25"),
  1516 => (x"63",x"65",x"68",x"43"),
  1517 => (x"6d",x"75",x"73",x"6b"),
  1518 => (x"67",x"6e",x"69",x"6d"),
  1519 => (x"6f",x"72",x"66",x"20"),
  1520 => (x"64",x"25",x"20",x"6d"),
  1521 => (x"20",x"6f",x"74",x"20"),
  1522 => (x"2e",x"2e",x"64",x"25"),
  1523 => (x"25",x"00",x"20",x"2e"),
  1524 => (x"25",x"00",x"0a",x"64"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
