
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"3b",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"38"),
    10 => (x"20",x"00",x"27",x"4f"),
    11 => (x"27",x"4e",x"00",x"00"),
    12 => (x"00",x"00",x"13",x"ce"),
    13 => (x"87",x"fd",x"00",x"0f"),
    14 => (x"4f",x"87",x"fd",x"00"),
    15 => (x"ff",x"86",x"fc",x"1e"),
    16 => (x"48",x"69",x"49",x"c0"),
    17 => (x"c4",x"98",x"c0",x"c4"),
    18 => (x"02",x"6e",x"58",x"a6"),
    19 => (x"66",x"c8",x"87",x"f4"),
    20 => (x"8e",x"fc",x"48",x"79"),
    21 => (x"5e",x"0e",x"4f",x"26"),
    22 => (x"0e",x"5d",x"5c",x"5b"),
    23 => (x"c0",x"4b",x"66",x"d0"),
    24 => (x"c3",x"49",x"13",x"4c"),
    25 => (x"99",x"71",x"99",x"ff"),
    26 => (x"71",x"87",x"dd",x"02"),
    27 => (x"4a",x"c0",x"ff",x"4d"),
    28 => (x"c0",x"c4",x"49",x"6a"),
    29 => (x"02",x"99",x"71",x"99"),
    30 => (x"7a",x"75",x"87",x"f6"),
    31 => (x"49",x"13",x"84",x"c1"),
    32 => (x"71",x"99",x"ff",x"c3"),
    33 => (x"87",x"e3",x"05",x"99"),
    34 => (x"4d",x"26",x"48",x"74"),
    35 => (x"4b",x"26",x"4c",x"26"),
    36 => (x"5e",x"0e",x"4f",x"26"),
    37 => (x"0e",x"5d",x"5c",x"5b"),
    38 => (x"4b",x"c0",x"86",x"f0"),
    39 => (x"c0",x"48",x"a6",x"c4"),
    40 => (x"a6",x"e4",x"c0",x"78"),
    41 => (x"66",x"e0",x"c0",x"4c"),
    42 => (x"80",x"c1",x"48",x"49"),
    43 => (x"58",x"a6",x"e4",x"c0"),
    44 => (x"c0",x"fe",x"4a",x"11"),
    45 => (x"9a",x"72",x"ba",x"82"),
    46 => (x"87",x"d3",x"c4",x"02"),
    47 => (x"c3",x"02",x"66",x"c4"),
    48 => (x"a6",x"c4",x"87",x"e2"),
    49 => (x"72",x"78",x"c0",x"48"),
    50 => (x"aa",x"f0",x"c0",x"49"),
    51 => (x"87",x"f2",x"c2",x"02"),
    52 => (x"02",x"a9",x"e3",x"c1"),
    53 => (x"c1",x"87",x"f3",x"c2"),
    54 => (x"c0",x"02",x"a9",x"e4"),
    55 => (x"ec",x"c1",x"87",x"e1"),
    56 => (x"dd",x"c2",x"02",x"a9"),
    57 => (x"a9",x"f0",x"c1",x"87"),
    58 => (x"c1",x"87",x"d4",x"02"),
    59 => (x"c1",x"02",x"a9",x"f3"),
    60 => (x"f5",x"c1",x"87",x"fc"),
    61 => (x"87",x"c7",x"02",x"a9"),
    62 => (x"05",x"a9",x"f8",x"c1"),
    63 => (x"c4",x"87",x"dc",x"c2"),
    64 => (x"c4",x"49",x"74",x"84"),
    65 => (x"69",x"48",x"76",x"89"),
    66 => (x"c1",x"02",x"6e",x"78"),
    67 => (x"80",x"c8",x"87",x"d3"),
    68 => (x"a6",x"cc",x"78",x"c0"),
    69 => (x"6e",x"78",x"c0",x"48"),
    70 => (x"29",x"b7",x"dc",x"49"),
    71 => (x"9a",x"cf",x"4a",x"71"),
    72 => (x"30",x"c4",x"48",x"6e"),
    73 => (x"72",x"58",x"a6",x"c4"),
    74 => (x"87",x"c5",x"02",x"9a"),
    75 => (x"c1",x"48",x"a6",x"c8"),
    76 => (x"06",x"aa",x"c9",x"78"),
    77 => (x"f7",x"c0",x"87",x"c5"),
    78 => (x"c0",x"87",x"c3",x"82"),
    79 => (x"66",x"c8",x"82",x"f0"),
    80 => (x"72",x"87",x"c9",x"02"),
    81 => (x"87",x"f4",x"fb",x"1e"),
    82 => (x"83",x"c1",x"86",x"c4"),
    83 => (x"c1",x"48",x"66",x"cc"),
    84 => (x"58",x"a6",x"d0",x"80"),
    85 => (x"c8",x"48",x"66",x"cc"),
    86 => (x"fe",x"04",x"a8",x"b7"),
    87 => (x"d7",x"c1",x"87",x"f9"),
    88 => (x"1e",x"f0",x"c0",x"87"),
    89 => (x"c4",x"87",x"d5",x"fb"),
    90 => (x"c1",x"83",x"c1",x"86"),
    91 => (x"84",x"c4",x"87",x"ca"),
    92 => (x"89",x"c4",x"49",x"74"),
    93 => (x"dd",x"fb",x"1e",x"69"),
    94 => (x"70",x"86",x"c4",x"87"),
    95 => (x"c0",x"83",x"71",x"49"),
    96 => (x"a6",x"c4",x"87",x"f6"),
    97 => (x"c0",x"78",x"c1",x"48"),
    98 => (x"84",x"c4",x"87",x"ee"),
    99 => (x"89",x"c4",x"49",x"74"),
   100 => (x"e7",x"fa",x"1e",x"69"),
   101 => (x"c1",x"86",x"c4",x"87"),
   102 => (x"72",x"87",x"dd",x"83"),
   103 => (x"87",x"dc",x"fa",x"1e"),
   104 => (x"87",x"d4",x"86",x"c4"),
   105 => (x"05",x"aa",x"e5",x"c0"),
   106 => (x"a6",x"c4",x"87",x"c7"),
   107 => (x"c7",x"78",x"c1",x"48"),
   108 => (x"fa",x"1e",x"72",x"87"),
   109 => (x"86",x"c4",x"87",x"c6"),
   110 => (x"49",x"66",x"e0",x"c0"),
   111 => (x"c0",x"80",x"c1",x"48"),
   112 => (x"11",x"58",x"a6",x"e4"),
   113 => (x"82",x"c0",x"fe",x"4a"),
   114 => (x"05",x"9a",x"72",x"ba"),
   115 => (x"73",x"87",x"ed",x"fb"),
   116 => (x"26",x"8e",x"f0",x"48"),
   117 => (x"26",x"4c",x"26",x"4d"),
   118 => (x"0e",x"4f",x"26",x"4b"),
   119 => (x"86",x"e8",x"0e",x"5e"),
   120 => (x"c3",x"4a",x"d4",x"ff"),
   121 => (x"49",x"6a",x"7a",x"ff"),
   122 => (x"6a",x"7a",x"ff",x"c3"),
   123 => (x"c4",x"30",x"c8",x"48"),
   124 => (x"a6",x"c8",x"58",x"a6"),
   125 => (x"c3",x"b1",x"6e",x"59"),
   126 => (x"48",x"6a",x"7a",x"ff"),
   127 => (x"a6",x"cc",x"30",x"d0"),
   128 => (x"59",x"a6",x"d0",x"58"),
   129 => (x"c3",x"b1",x"66",x"c8"),
   130 => (x"48",x"6a",x"7a",x"ff"),
   131 => (x"a6",x"d4",x"30",x"d8"),
   132 => (x"59",x"a6",x"d8",x"58"),
   133 => (x"71",x"b1",x"66",x"d0"),
   134 => (x"c6",x"8e",x"e8",x"48"),
   135 => (x"26",x"4d",x"26",x"87"),
   136 => (x"26",x"4b",x"26",x"4c"),
   137 => (x"0e",x"5e",x"0e",x"4f"),
   138 => (x"d4",x"ff",x"86",x"f4"),
   139 => (x"7a",x"ff",x"c3",x"4a"),
   140 => (x"ff",x"c3",x"49",x"6a"),
   141 => (x"c8",x"48",x"71",x"7a"),
   142 => (x"58",x"a6",x"c4",x"30"),
   143 => (x"b1",x"6e",x"49",x"6a"),
   144 => (x"71",x"7a",x"ff",x"c3"),
   145 => (x"c8",x"30",x"c8",x"48"),
   146 => (x"49",x"6a",x"58",x"a6"),
   147 => (x"c3",x"b1",x"66",x"c4"),
   148 => (x"48",x"71",x"7a",x"ff"),
   149 => (x"a6",x"cc",x"30",x"c8"),
   150 => (x"c8",x"49",x"6a",x"58"),
   151 => (x"48",x"71",x"b1",x"66"),
   152 => (x"fe",x"fe",x"8e",x"f4"),
   153 => (x"5b",x"5e",x"0e",x"87"),
   154 => (x"d4",x"ff",x"0e",x"5c"),
   155 => (x"48",x"66",x"cc",x"4c"),
   156 => (x"70",x"98",x"ff",x"c3"),
   157 => (x"d4",x"d4",x"c1",x"7c"),
   158 => (x"87",x"c8",x"05",x"bf"),
   159 => (x"c9",x"48",x"66",x"d0"),
   160 => (x"58",x"a6",x"d4",x"30"),
   161 => (x"d8",x"49",x"66",x"d0"),
   162 => (x"c3",x"48",x"71",x"29"),
   163 => (x"7c",x"70",x"98",x"ff"),
   164 => (x"d0",x"49",x"66",x"d0"),
   165 => (x"c3",x"48",x"71",x"29"),
   166 => (x"7c",x"70",x"98",x"ff"),
   167 => (x"c8",x"49",x"66",x"d0"),
   168 => (x"c3",x"48",x"71",x"29"),
   169 => (x"7c",x"70",x"98",x"ff"),
   170 => (x"c3",x"48",x"66",x"d0"),
   171 => (x"7c",x"70",x"98",x"ff"),
   172 => (x"d0",x"49",x"66",x"cc"),
   173 => (x"c3",x"48",x"71",x"29"),
   174 => (x"7c",x"70",x"98",x"ff"),
   175 => (x"f0",x"c9",x"4a",x"6c"),
   176 => (x"ff",x"c3",x"4b",x"ff"),
   177 => (x"87",x"d2",x"05",x"aa"),
   178 => (x"6c",x"7c",x"ff",x"c3"),
   179 => (x"73",x"8b",x"c1",x"4a"),
   180 => (x"87",x"c6",x"02",x"9b"),
   181 => (x"02",x"aa",x"ff",x"c3"),
   182 => (x"48",x"72",x"87",x"ee"),
   183 => (x"1e",x"87",x"c0",x"fd"),
   184 => (x"d4",x"ff",x"49",x"c0"),
   185 => (x"78",x"ff",x"c3",x"48"),
   186 => (x"c8",x"c3",x"81",x"c1"),
   187 => (x"f1",x"04",x"a9",x"b7"),
   188 => (x"87",x"ef",x"fc",x"87"),
   189 => (x"0e",x"5b",x"5e",x"0e"),
   190 => (x"f8",x"c4",x"87",x"e5"),
   191 => (x"1e",x"c0",x"4b",x"df"),
   192 => (x"c1",x"f0",x"ff",x"c0"),
   193 => (x"dc",x"fd",x"1e",x"f7"),
   194 => (x"c1",x"86",x"c8",x"87"),
   195 => (x"ea",x"c0",x"05",x"a8"),
   196 => (x"48",x"d4",x"ff",x"87"),
   197 => (x"c1",x"78",x"ff",x"c3"),
   198 => (x"c0",x"c0",x"c0",x"c0"),
   199 => (x"e1",x"c0",x"1e",x"c0"),
   200 => (x"1e",x"e9",x"c1",x"f0"),
   201 => (x"c8",x"87",x"fe",x"fc"),
   202 => (x"05",x"98",x"70",x"86"),
   203 => (x"d4",x"ff",x"87",x"ca"),
   204 => (x"78",x"ff",x"c3",x"48"),
   205 => (x"87",x"cd",x"48",x"c1"),
   206 => (x"c1",x"87",x"e4",x"fe"),
   207 => (x"05",x"9b",x"73",x"8b"),
   208 => (x"c0",x"87",x"fb",x"fe"),
   209 => (x"87",x"d9",x"fb",x"48"),
   210 => (x"0e",x"5b",x"5e",x"0e"),
   211 => (x"c3",x"48",x"d4",x"ff"),
   212 => (x"e5",x"c0",x"78",x"ff"),
   213 => (x"fd",x"f3",x"1e",x"d5"),
   214 => (x"d3",x"86",x"c4",x"87"),
   215 => (x"c0",x"1e",x"c0",x"4b"),
   216 => (x"c1",x"c1",x"f0",x"ff"),
   217 => (x"87",x"fd",x"fb",x"1e"),
   218 => (x"98",x"70",x"86",x"c8"),
   219 => (x"ff",x"87",x"ca",x"05"),
   220 => (x"ff",x"c3",x"48",x"d4"),
   221 => (x"cd",x"48",x"c1",x"78"),
   222 => (x"87",x"e3",x"fd",x"87"),
   223 => (x"9b",x"73",x"8b",x"c1"),
   224 => (x"87",x"d9",x"ff",x"05"),
   225 => (x"d8",x"fa",x"48",x"c0"),
   226 => (x"5b",x"5e",x"0e",x"87"),
   227 => (x"ff",x"0e",x"5d",x"5c"),
   228 => (x"ca",x"fd",x"4d",x"d4"),
   229 => (x"1e",x"ea",x"c6",x"87"),
   230 => (x"c1",x"f0",x"e1",x"c0"),
   231 => (x"c4",x"fb",x"1e",x"c8"),
   232 => (x"70",x"86",x"c8",x"87"),
   233 => (x"d2",x"1e",x"73",x"4b"),
   234 => (x"e5",x"f3",x"1e",x"d4"),
   235 => (x"c1",x"86",x"c8",x"87"),
   236 => (x"87",x"c8",x"02",x"ab"),
   237 => (x"c0",x"87",x"d1",x"fe"),
   238 => (x"87",x"d3",x"c2",x"48"),
   239 => (x"70",x"87",x"e6",x"f9"),
   240 => (x"ff",x"ff",x"cf",x"49"),
   241 => (x"a9",x"ea",x"c6",x"99"),
   242 => (x"fd",x"87",x"c8",x"02"),
   243 => (x"48",x"c0",x"87",x"fa"),
   244 => (x"c3",x"87",x"fc",x"c1"),
   245 => (x"f1",x"c0",x"7d",x"ff"),
   246 => (x"87",x"d8",x"fc",x"4c"),
   247 => (x"c1",x"02",x"98",x"70"),
   248 => (x"1e",x"c0",x"87",x"d2"),
   249 => (x"c1",x"f0",x"ff",x"c0"),
   250 => (x"f8",x"f9",x"1e",x"fa"),
   251 => (x"70",x"86",x"c8",x"87"),
   252 => (x"05",x"9b",x"73",x"4b"),
   253 => (x"73",x"87",x"f3",x"c0"),
   254 => (x"1e",x"d2",x"d1",x"1e"),
   255 => (x"c8",x"87",x"d3",x"f2"),
   256 => (x"7d",x"ff",x"c3",x"86"),
   257 => (x"1e",x"73",x"4b",x"6d"),
   258 => (x"f2",x"1e",x"de",x"d1"),
   259 => (x"86",x"c8",x"87",x"c4"),
   260 => (x"7d",x"7d",x"ff",x"c3"),
   261 => (x"49",x"73",x"7d",x"7d"),
   262 => (x"71",x"99",x"c0",x"c1"),
   263 => (x"87",x"c5",x"02",x"99"),
   264 => (x"ea",x"c0",x"48",x"c1"),
   265 => (x"c0",x"48",x"c0",x"87"),
   266 => (x"1e",x"73",x"87",x"e5"),
   267 => (x"f1",x"1e",x"ec",x"d1"),
   268 => (x"86",x"c8",x"87",x"e0"),
   269 => (x"cc",x"05",x"ac",x"c2"),
   270 => (x"1e",x"f8",x"d1",x"87"),
   271 => (x"c4",x"87",x"d3",x"f1"),
   272 => (x"ca",x"48",x"c0",x"86"),
   273 => (x"74",x"8c",x"c1",x"87"),
   274 => (x"cc",x"fe",x"05",x"9c"),
   275 => (x"f7",x"48",x"c0",x"87"),
   276 => (x"4d",x"43",x"87",x"cb"),
   277 => (x"20",x"38",x"35",x"44"),
   278 => (x"20",x"0a",x"64",x"25"),
   279 => (x"4d",x"43",x"00",x"20"),
   280 => (x"5f",x"38",x"35",x"44"),
   281 => (x"64",x"25",x"20",x"32"),
   282 => (x"00",x"20",x"20",x"0a"),
   283 => (x"35",x"44",x"4d",x"43"),
   284 => (x"64",x"25",x"20",x"38"),
   285 => (x"00",x"20",x"20",x"0a"),
   286 => (x"43",x"48",x"44",x"53"),
   287 => (x"69",x"6e",x"49",x"20"),
   288 => (x"6c",x"61",x"69",x"74"),
   289 => (x"74",x"61",x"7a",x"69"),
   290 => (x"20",x"6e",x"6f",x"69"),
   291 => (x"6f",x"72",x"72",x"65"),
   292 => (x"00",x"0a",x"21",x"72"),
   293 => (x"5f",x"64",x"6d",x"63"),
   294 => (x"38",x"44",x"4d",x"43"),
   295 => (x"73",x"65",x"72",x"20"),
   296 => (x"73",x"6e",x"6f",x"70"),
   297 => (x"25",x"20",x"3a",x"65"),
   298 => (x"0e",x"00",x"0a",x"64"),
   299 => (x"5d",x"5c",x"5b",x"5e"),
   300 => (x"d0",x"ff",x"1e",x"0e"),
   301 => (x"c0",x"c0",x"c8",x"4d"),
   302 => (x"d4",x"d4",x"c1",x"4b"),
   303 => (x"d6",x"78",x"c1",x"48"),
   304 => (x"d1",x"ee",x"1e",x"d1"),
   305 => (x"c7",x"86",x"c4",x"87"),
   306 => (x"73",x"48",x"6d",x"4c"),
   307 => (x"58",x"a6",x"c4",x"98"),
   308 => (x"cc",x"c0",x"02",x"6e"),
   309 => (x"73",x"48",x"6d",x"87"),
   310 => (x"58",x"a6",x"c4",x"98"),
   311 => (x"f4",x"ff",x"05",x"6e"),
   312 => (x"f7",x"7d",x"c0",x"87"),
   313 => (x"48",x"6d",x"87",x"f9"),
   314 => (x"a6",x"c4",x"98",x"73"),
   315 => (x"c0",x"02",x"6e",x"58"),
   316 => (x"48",x"6d",x"87",x"cc"),
   317 => (x"a6",x"c4",x"98",x"73"),
   318 => (x"ff",x"05",x"6e",x"58"),
   319 => (x"7d",x"c1",x"87",x"f4"),
   320 => (x"e5",x"c0",x"1e",x"c0"),
   321 => (x"1e",x"c0",x"c1",x"d0"),
   322 => (x"c8",x"87",x"da",x"f5"),
   323 => (x"05",x"a8",x"c1",x"86"),
   324 => (x"c1",x"87",x"c2",x"c0"),
   325 => (x"05",x"ac",x"c2",x"4c"),
   326 => (x"d6",x"87",x"cd",x"c0"),
   327 => (x"f5",x"ec",x"1e",x"cc"),
   328 => (x"c0",x"86",x"c4",x"87"),
   329 => (x"87",x"e0",x"c1",x"48"),
   330 => (x"9c",x"74",x"8c",x"c1"),
   331 => (x"87",x"d9",x"fe",x"05"),
   332 => (x"c1",x"87",x"d6",x"f9"),
   333 => (x"c1",x"58",x"d8",x"d4"),
   334 => (x"05",x"bf",x"d4",x"d4"),
   335 => (x"c1",x"87",x"cd",x"c0"),
   336 => (x"f0",x"ff",x"c0",x"1e"),
   337 => (x"f4",x"1e",x"d0",x"c1"),
   338 => (x"86",x"c8",x"87",x"db"),
   339 => (x"c3",x"48",x"d4",x"ff"),
   340 => (x"c4",x"ca",x"78",x"ff"),
   341 => (x"dc",x"d4",x"c1",x"87"),
   342 => (x"d8",x"d4",x"c1",x"58"),
   343 => (x"d5",x"d6",x"1e",x"bf"),
   344 => (x"87",x"ee",x"ec",x"1e"),
   345 => (x"48",x"6d",x"86",x"c8"),
   346 => (x"a6",x"c4",x"98",x"73"),
   347 => (x"c0",x"02",x"6e",x"58"),
   348 => (x"48",x"6d",x"87",x"cc"),
   349 => (x"a6",x"c4",x"98",x"73"),
   350 => (x"ff",x"05",x"6e",x"58"),
   351 => (x"7d",x"c0",x"87",x"f4"),
   352 => (x"c3",x"48",x"d4",x"ff"),
   353 => (x"48",x"c1",x"78",x"ff"),
   354 => (x"87",x"d1",x"f2",x"26"),
   355 => (x"52",x"52",x"45",x"49"),
   356 => (x"49",x"50",x"53",x"00"),
   357 => (x"20",x"44",x"53",x"00"),
   358 => (x"64",x"72",x"61",x"63"),
   359 => (x"7a",x"69",x"73",x"20"),
   360 => (x"73",x"69",x"20",x"65"),
   361 => (x"0a",x"64",x"25",x"20"),
   362 => (x"5b",x"5e",x"0e",x"00"),
   363 => (x"1e",x"0e",x"5d",x"5c"),
   364 => (x"ff",x"4c",x"ff",x"c3"),
   365 => (x"7b",x"74",x"4b",x"d4"),
   366 => (x"48",x"bf",x"d0",x"ff"),
   367 => (x"98",x"c0",x"c0",x"c8"),
   368 => (x"6e",x"58",x"a6",x"c4"),
   369 => (x"87",x"d0",x"c0",x"02"),
   370 => (x"48",x"bf",x"d0",x"ff"),
   371 => (x"98",x"c0",x"c0",x"c8"),
   372 => (x"6e",x"58",x"a6",x"c4"),
   373 => (x"87",x"f0",x"ff",x"05"),
   374 => (x"c4",x"48",x"d0",x"ff"),
   375 => (x"7b",x"74",x"78",x"c1"),
   376 => (x"c0",x"1e",x"66",x"d4"),
   377 => (x"d8",x"c1",x"f0",x"ff"),
   378 => (x"87",x"f9",x"f1",x"1e"),
   379 => (x"98",x"70",x"86",x"c8"),
   380 => (x"87",x"cd",x"c0",x"02"),
   381 => (x"e9",x"1e",x"ca",x"da"),
   382 => (x"86",x"c4",x"87",x"dc"),
   383 => (x"c5",x"c2",x"48",x"c1"),
   384 => (x"c3",x"7b",x"74",x"87"),
   385 => (x"4d",x"c0",x"7b",x"fe"),
   386 => (x"49",x"bf",x"66",x"d8"),
   387 => (x"b7",x"d8",x"4a",x"71"),
   388 => (x"74",x"48",x"72",x"2a"),
   389 => (x"71",x"7b",x"70",x"98"),
   390 => (x"2a",x"b7",x"d0",x"4a"),
   391 => (x"98",x"74",x"48",x"72"),
   392 => (x"4a",x"71",x"7b",x"70"),
   393 => (x"72",x"2a",x"b7",x"c8"),
   394 => (x"70",x"98",x"74",x"48"),
   395 => (x"74",x"48",x"71",x"7b"),
   396 => (x"d8",x"7b",x"70",x"98"),
   397 => (x"80",x"c4",x"48",x"66"),
   398 => (x"c1",x"58",x"a6",x"dc"),
   399 => (x"b7",x"c0",x"c2",x"85"),
   400 => (x"c3",x"ff",x"04",x"ad"),
   401 => (x"74",x"7b",x"74",x"87"),
   402 => (x"d8",x"7b",x"74",x"7b"),
   403 => (x"74",x"49",x"e0",x"da"),
   404 => (x"c0",x"05",x"6b",x"7b"),
   405 => (x"89",x"c1",x"87",x"c8"),
   406 => (x"ff",x"05",x"99",x"71"),
   407 => (x"7b",x"74",x"87",x"f1"),
   408 => (x"48",x"bf",x"d0",x"ff"),
   409 => (x"98",x"c0",x"c0",x"c8"),
   410 => (x"6e",x"58",x"a6",x"c4"),
   411 => (x"87",x"d0",x"c0",x"02"),
   412 => (x"48",x"bf",x"d0",x"ff"),
   413 => (x"98",x"c0",x"c0",x"c8"),
   414 => (x"6e",x"58",x"a6",x"c4"),
   415 => (x"87",x"f0",x"ff",x"05"),
   416 => (x"c0",x"48",x"d0",x"ff"),
   417 => (x"ee",x"26",x"48",x"78"),
   418 => (x"72",x"57",x"87",x"d3"),
   419 => (x"20",x"65",x"74",x"69"),
   420 => (x"6c",x"69",x"61",x"66"),
   421 => (x"00",x"0a",x"64",x"65"),
   422 => (x"5c",x"5b",x"5e",x"0e"),
   423 => (x"4c",x"66",x"d0",x"0e"),
   424 => (x"c0",x"4b",x"66",x"cc"),
   425 => (x"cd",x"ee",x"c5",x"4a"),
   426 => (x"d4",x"ff",x"49",x"df"),
   427 => (x"78",x"ff",x"c3",x"48"),
   428 => (x"c3",x"48",x"bf",x"70"),
   429 => (x"c1",x"05",x"a8",x"fe"),
   430 => (x"d4",x"c1",x"87",x"d8"),
   431 => (x"78",x"c0",x"48",x"d0"),
   432 => (x"04",x"ac",x"b7",x"c4"),
   433 => (x"ec",x"87",x"dc",x"c0"),
   434 => (x"49",x"70",x"87",x"d1"),
   435 => (x"83",x"c4",x"7b",x"71"),
   436 => (x"bf",x"d0",x"d4",x"c1"),
   437 => (x"c1",x"80",x"71",x"48"),
   438 => (x"c4",x"58",x"d4",x"d4"),
   439 => (x"03",x"ac",x"b7",x"8c"),
   440 => (x"c0",x"87",x"e4",x"ff"),
   441 => (x"c0",x"06",x"ac",x"b7"),
   442 => (x"d4",x"ff",x"87",x"e5"),
   443 => (x"78",x"ff",x"c3",x"48"),
   444 => (x"71",x"49",x"bf",x"70"),
   445 => (x"ff",x"c3",x"7b",x"97"),
   446 => (x"c1",x"83",x"c1",x"98"),
   447 => (x"48",x"bf",x"d0",x"d4"),
   448 => (x"d4",x"c1",x"80",x"71"),
   449 => (x"8c",x"c1",x"58",x"d4"),
   450 => (x"01",x"ac",x"b7",x"c0"),
   451 => (x"c1",x"87",x"db",x"ff"),
   452 => (x"89",x"c1",x"4a",x"49"),
   453 => (x"fe",x"05",x"99",x"71"),
   454 => (x"d4",x"ff",x"87",x"d0"),
   455 => (x"78",x"ff",x"c3",x"48"),
   456 => (x"fa",x"eb",x"48",x"72"),
   457 => (x"5b",x"5e",x"0e",x"87"),
   458 => (x"c8",x"1e",x"0e",x"5c"),
   459 => (x"c0",x"4c",x"c0",x"c0"),
   460 => (x"48",x"d4",x"ff",x"4b"),
   461 => (x"ff",x"78",x"ff",x"c3"),
   462 => (x"74",x"48",x"bf",x"d0"),
   463 => (x"58",x"a6",x"c4",x"98"),
   464 => (x"ce",x"c0",x"02",x"6e"),
   465 => (x"bf",x"d0",x"ff",x"87"),
   466 => (x"c4",x"98",x"74",x"48"),
   467 => (x"05",x"6e",x"58",x"a6"),
   468 => (x"ff",x"87",x"f2",x"ff"),
   469 => (x"c1",x"c4",x"48",x"d0"),
   470 => (x"48",x"d4",x"ff",x"78"),
   471 => (x"d0",x"78",x"ff",x"c3"),
   472 => (x"ff",x"c0",x"1e",x"66"),
   473 => (x"1e",x"d1",x"c1",x"f0"),
   474 => (x"c8",x"87",x"fa",x"eb"),
   475 => (x"71",x"49",x"70",x"86"),
   476 => (x"d0",x"c0",x"02",x"99"),
   477 => (x"d4",x"1e",x"71",x"87"),
   478 => (x"f9",x"de",x"1e",x"66"),
   479 => (x"87",x"d2",x"e4",x"1e"),
   480 => (x"ee",x"c0",x"86",x"cc"),
   481 => (x"1e",x"c0",x"c8",x"87"),
   482 => (x"fc",x"1e",x"66",x"d8"),
   483 => (x"86",x"c8",x"87",x"ca"),
   484 => (x"d0",x"ff",x"4b",x"70"),
   485 => (x"98",x"74",x"48",x"bf"),
   486 => (x"6e",x"58",x"a6",x"c4"),
   487 => (x"87",x"ce",x"c0",x"02"),
   488 => (x"48",x"bf",x"d0",x"ff"),
   489 => (x"a6",x"c4",x"98",x"74"),
   490 => (x"ff",x"05",x"6e",x"58"),
   491 => (x"d0",x"ff",x"87",x"f2"),
   492 => (x"73",x"78",x"c0",x"48"),
   493 => (x"e6",x"e9",x"26",x"48"),
   494 => (x"61",x"65",x"52",x"87"),
   495 => (x"6f",x"63",x"20",x"64"),
   496 => (x"6e",x"61",x"6d",x"6d"),
   497 => (x"61",x"66",x"20",x"64"),
   498 => (x"64",x"65",x"6c",x"69"),
   499 => (x"20",x"74",x"61",x"20"),
   500 => (x"28",x"20",x"64",x"25"),
   501 => (x"0a",x"29",x"64",x"25"),
   502 => (x"5b",x"5e",x"0e",x"00"),
   503 => (x"1e",x"0e",x"5d",x"5c"),
   504 => (x"ff",x"c0",x"1e",x"c0"),
   505 => (x"1e",x"c9",x"c1",x"f0"),
   506 => (x"c8",x"87",x"fa",x"e9"),
   507 => (x"c1",x"1e",x"d2",x"86"),
   508 => (x"fa",x"1e",x"e2",x"d4"),
   509 => (x"86",x"c8",x"87",x"e2"),
   510 => (x"85",x"c1",x"4d",x"c0"),
   511 => (x"04",x"ad",x"b7",x"d2"),
   512 => (x"c1",x"87",x"f7",x"ff"),
   513 => (x"bf",x"97",x"e2",x"d4"),
   514 => (x"99",x"c0",x"c3",x"49"),
   515 => (x"05",x"a9",x"c0",x"c1"),
   516 => (x"c1",x"87",x"e8",x"c0"),
   517 => (x"bf",x"97",x"e9",x"d4"),
   518 => (x"c1",x"31",x"d0",x"49"),
   519 => (x"bf",x"97",x"ea",x"d4"),
   520 => (x"72",x"32",x"c8",x"4a"),
   521 => (x"eb",x"d4",x"c1",x"b1"),
   522 => (x"72",x"4a",x"bf",x"97"),
   523 => (x"ff",x"ff",x"cf",x"b1"),
   524 => (x"4d",x"71",x"99",x"ff"),
   525 => (x"35",x"ca",x"85",x"c1"),
   526 => (x"c1",x"87",x"f0",x"c2"),
   527 => (x"bf",x"97",x"eb",x"d4"),
   528 => (x"c6",x"33",x"c1",x"4b"),
   529 => (x"ec",x"d4",x"c1",x"9b"),
   530 => (x"c7",x"49",x"bf",x"97"),
   531 => (x"b3",x"71",x"29",x"b7"),
   532 => (x"97",x"e7",x"d4",x"c1"),
   533 => (x"48",x"71",x"49",x"bf"),
   534 => (x"a6",x"c4",x"98",x"cf"),
   535 => (x"e8",x"d4",x"c1",x"58"),
   536 => (x"c3",x"4c",x"bf",x"97"),
   537 => (x"c1",x"34",x"ca",x"9c"),
   538 => (x"bf",x"97",x"e9",x"d4"),
   539 => (x"71",x"31",x"c2",x"49"),
   540 => (x"ea",x"d4",x"c1",x"b4"),
   541 => (x"c3",x"49",x"bf",x"97"),
   542 => (x"b7",x"c6",x"99",x"c0"),
   543 => (x"74",x"b4",x"71",x"29"),
   544 => (x"1e",x"66",x"c4",x"1e"),
   545 => (x"e3",x"c0",x"1e",x"73"),
   546 => (x"c5",x"e0",x"1e",x"f1"),
   547 => (x"c2",x"86",x"d0",x"87"),
   548 => (x"73",x"48",x"c1",x"83"),
   549 => (x"73",x"4b",x"70",x"30"),
   550 => (x"de",x"e4",x"c0",x"1e"),
   551 => (x"f1",x"df",x"ff",x"1e"),
   552 => (x"c1",x"86",x"c8",x"87"),
   553 => (x"c4",x"30",x"6e",x"48"),
   554 => (x"49",x"74",x"58",x"a6"),
   555 => (x"4d",x"71",x"81",x"c1"),
   556 => (x"6e",x"95",x"b7",x"73"),
   557 => (x"c0",x"1e",x"75",x"1e"),
   558 => (x"ff",x"1e",x"e7",x"e4"),
   559 => (x"cc",x"87",x"d3",x"df"),
   560 => (x"c8",x"48",x"6e",x"86"),
   561 => (x"06",x"a8",x"b7",x"c0"),
   562 => (x"c1",x"87",x"d4",x"c0"),
   563 => (x"c1",x"48",x"6e",x"35"),
   564 => (x"a6",x"c4",x"28",x"b7"),
   565 => (x"c8",x"48",x"6e",x"58"),
   566 => (x"01",x"a8",x"b7",x"c0"),
   567 => (x"75",x"87",x"ec",x"ff"),
   568 => (x"fd",x"e4",x"c0",x"1e"),
   569 => (x"e9",x"de",x"ff",x"1e"),
   570 => (x"75",x"86",x"c8",x"87"),
   571 => (x"ec",x"e4",x"26",x"48"),
   572 => (x"73",x"5f",x"63",x"87"),
   573 => (x"5f",x"65",x"7a",x"69"),
   574 => (x"74",x"6c",x"75",x"6d"),
   575 => (x"64",x"25",x"20",x"3a"),
   576 => (x"65",x"72",x"20",x"2c"),
   577 => (x"62",x"5f",x"64",x"61"),
   578 => (x"65",x"6c",x"5f",x"6c"),
   579 => (x"25",x"20",x"3a",x"6e"),
   580 => (x"63",x"20",x"2c",x"64"),
   581 => (x"65",x"7a",x"69",x"73"),
   582 => (x"64",x"25",x"20",x"3a"),
   583 => (x"75",x"4d",x"00",x"0a"),
   584 => (x"25",x"20",x"74",x"6c"),
   585 => (x"25",x"00",x"0a",x"64"),
   586 => (x"6c",x"62",x"20",x"64"),
   587 => (x"73",x"6b",x"63",x"6f"),
   588 => (x"20",x"66",x"6f",x"20"),
   589 => (x"65",x"7a",x"69",x"73"),
   590 => (x"0a",x"64",x"25",x"20"),
   591 => (x"20",x"64",x"25",x"00"),
   592 => (x"63",x"6f",x"6c",x"62"),
   593 => (x"6f",x"20",x"73",x"6b"),
   594 => (x"31",x"35",x"20",x"66"),
   595 => (x"79",x"62",x"20",x"32"),
   596 => (x"0a",x"73",x"65",x"74"),
   597 => (x"44",x"4d",x"43",x"00"),
   598 => (x"5b",x"5e",x"0e",x"00"),
   599 => (x"d0",x"4b",x"c0",x"0e"),
   600 => (x"b7",x"c0",x"48",x"66"),
   601 => (x"f6",x"c0",x"06",x"a8"),
   602 => (x"97",x"66",x"c8",x"87"),
   603 => (x"c0",x"fe",x"4a",x"bf"),
   604 => (x"66",x"c8",x"ba",x"82"),
   605 => (x"cc",x"80",x"c1",x"48"),
   606 => (x"66",x"cc",x"58",x"a6"),
   607 => (x"fe",x"49",x"bf",x"97"),
   608 => (x"cc",x"b9",x"81",x"c0"),
   609 => (x"80",x"c1",x"48",x"66"),
   610 => (x"71",x"58",x"a6",x"d0"),
   611 => (x"c4",x"02",x"aa",x"b7"),
   612 => (x"cc",x"48",x"c1",x"87"),
   613 => (x"d0",x"83",x"c1",x"87"),
   614 => (x"04",x"ab",x"b7",x"66"),
   615 => (x"c0",x"87",x"ca",x"ff"),
   616 => (x"26",x"87",x"c4",x"48"),
   617 => (x"26",x"4c",x"26",x"4d"),
   618 => (x"0e",x"4f",x"26",x"4b"),
   619 => (x"5d",x"5c",x"5b",x"5e"),
   620 => (x"fc",x"dc",x"c1",x"0e"),
   621 => (x"c1",x"78",x"c0",x"48"),
   622 => (x"ff",x"1e",x"c5",x"c1"),
   623 => (x"c4",x"87",x"d7",x"da"),
   624 => (x"f4",x"d4",x"c1",x"86"),
   625 => (x"f5",x"1e",x"c0",x"1e"),
   626 => (x"86",x"c8",x"87",x"db"),
   627 => (x"cf",x"05",x"98",x"70"),
   628 => (x"f1",x"fd",x"c0",x"87"),
   629 => (x"fd",x"d9",x"ff",x"1e"),
   630 => (x"c0",x"86",x"c4",x"87"),
   631 => (x"87",x"d6",x"cb",x"48"),
   632 => (x"1e",x"d2",x"c1",x"c1"),
   633 => (x"87",x"ee",x"d9",x"ff"),
   634 => (x"4b",x"c0",x"86",x"c4"),
   635 => (x"48",x"e8",x"dd",x"c1"),
   636 => (x"1e",x"c8",x"78",x"c1"),
   637 => (x"1e",x"e9",x"c1",x"c1"),
   638 => (x"1e",x"ea",x"d5",x"c1"),
   639 => (x"cc",x"87",x"da",x"fd"),
   640 => (x"05",x"98",x"70",x"86"),
   641 => (x"dd",x"c1",x"87",x"c6"),
   642 => (x"78",x"c0",x"48",x"e8"),
   643 => (x"c1",x"c1",x"1e",x"c8"),
   644 => (x"d6",x"c1",x"1e",x"f2"),
   645 => (x"c0",x"fd",x"1e",x"c6"),
   646 => (x"70",x"86",x"cc",x"87"),
   647 => (x"87",x"c6",x"05",x"98"),
   648 => (x"48",x"e8",x"dd",x"c1"),
   649 => (x"dd",x"c1",x"78",x"c0"),
   650 => (x"c1",x"1e",x"bf",x"e8"),
   651 => (x"ff",x"1e",x"fb",x"c1"),
   652 => (x"c8",x"87",x"df",x"d9"),
   653 => (x"e8",x"dd",x"c1",x"86"),
   654 => (x"d8",x"c2",x"02",x"bf"),
   655 => (x"f4",x"d4",x"c1",x"87"),
   656 => (x"f2",x"db",x"c1",x"4d"),
   657 => (x"f2",x"dc",x"c1",x"4c"),
   658 => (x"71",x"49",x"bf",x"9f"),
   659 => (x"f2",x"dc",x"c1",x"1e"),
   660 => (x"f4",x"d4",x"c1",x"49"),
   661 => (x"d0",x"1e",x"71",x"89"),
   662 => (x"1e",x"c0",x"c8",x"1e"),
   663 => (x"1e",x"e3",x"fe",x"c0"),
   664 => (x"87",x"ee",x"d8",x"ff"),
   665 => (x"49",x"74",x"86",x"d4"),
   666 => (x"4b",x"69",x"81",x"c8"),
   667 => (x"9f",x"f2",x"dc",x"c1"),
   668 => (x"d6",x"c5",x"49",x"bf"),
   669 => (x"c0",x"05",x"a9",x"ea"),
   670 => (x"49",x"74",x"87",x"d0"),
   671 => (x"1e",x"69",x"81",x"c8"),
   672 => (x"c4",x"87",x"d9",x"d9"),
   673 => (x"c0",x"4b",x"70",x"86"),
   674 => (x"49",x"75",x"87",x"df"),
   675 => (x"9f",x"81",x"fe",x"c7"),
   676 => (x"e9",x"ca",x"49",x"69"),
   677 => (x"c0",x"02",x"a9",x"d5"),
   678 => (x"fe",x"c0",x"87",x"cf"),
   679 => (x"d6",x"ff",x"1e",x"c5"),
   680 => (x"86",x"c4",x"87",x"f4"),
   681 => (x"cd",x"c8",x"48",x"c0"),
   682 => (x"c0",x"1e",x"73",x"87"),
   683 => (x"ff",x"1e",x"e0",x"ff"),
   684 => (x"c8",x"87",x"df",x"d7"),
   685 => (x"f4",x"d4",x"c1",x"86"),
   686 => (x"f1",x"1e",x"73",x"1e"),
   687 => (x"86",x"c8",x"87",x"e7"),
   688 => (x"c0",x"05",x"98",x"70"),
   689 => (x"48",x"c0",x"87",x"c5"),
   690 => (x"c0",x"87",x"eb",x"c7"),
   691 => (x"ff",x"1e",x"f8",x"ff"),
   692 => (x"c4",x"87",x"c3",x"d6"),
   693 => (x"ce",x"c2",x"c1",x"86"),
   694 => (x"f5",x"d6",x"ff",x"1e"),
   695 => (x"c8",x"86",x"c4",x"87"),
   696 => (x"e6",x"c2",x"c1",x"1e"),
   697 => (x"c6",x"d6",x"c1",x"1e"),
   698 => (x"87",x"ed",x"f9",x"1e"),
   699 => (x"98",x"70",x"86",x"cc"),
   700 => (x"87",x"c9",x"c0",x"05"),
   701 => (x"48",x"fc",x"dc",x"c1"),
   702 => (x"e4",x"c0",x"78",x"c1"),
   703 => (x"c1",x"1e",x"c8",x"87"),
   704 => (x"c1",x"1e",x"ef",x"c2"),
   705 => (x"f9",x"1e",x"ea",x"d5"),
   706 => (x"86",x"cc",x"87",x"cf"),
   707 => (x"c0",x"02",x"98",x"70"),
   708 => (x"c0",x"c1",x"87",x"cf"),
   709 => (x"d5",x"ff",x"1e",x"df"),
   710 => (x"86",x"c4",x"87",x"f8"),
   711 => (x"d5",x"c6",x"48",x"c0"),
   712 => (x"f2",x"dc",x"c1",x"87"),
   713 => (x"c1",x"49",x"bf",x"97"),
   714 => (x"c0",x"05",x"a9",x"d5"),
   715 => (x"dc",x"c1",x"87",x"cd"),
   716 => (x"49",x"bf",x"97",x"f3"),
   717 => (x"02",x"a9",x"ea",x"c2"),
   718 => (x"c0",x"87",x"c5",x"c0"),
   719 => (x"87",x"f6",x"c5",x"48"),
   720 => (x"97",x"f4",x"d4",x"c1"),
   721 => (x"e9",x"c3",x"49",x"bf"),
   722 => (x"d2",x"c0",x"02",x"a9"),
   723 => (x"f4",x"d4",x"c1",x"87"),
   724 => (x"c3",x"49",x"bf",x"97"),
   725 => (x"c0",x"02",x"a9",x"eb"),
   726 => (x"48",x"c0",x"87",x"c5"),
   727 => (x"c1",x"87",x"d7",x"c5"),
   728 => (x"bf",x"97",x"ff",x"d4"),
   729 => (x"05",x"99",x"71",x"49"),
   730 => (x"c1",x"87",x"cc",x"c0"),
   731 => (x"bf",x"97",x"c0",x"d5"),
   732 => (x"02",x"a9",x"c2",x"49"),
   733 => (x"c0",x"87",x"c5",x"c0"),
   734 => (x"87",x"fa",x"c4",x"48"),
   735 => (x"97",x"c1",x"d5",x"c1"),
   736 => (x"dc",x"c1",x"48",x"bf"),
   737 => (x"dc",x"c1",x"58",x"f8"),
   738 => (x"71",x"49",x"bf",x"f4"),
   739 => (x"c1",x"8a",x"c1",x"4a"),
   740 => (x"72",x"5a",x"fc",x"dc"),
   741 => (x"c1",x"1e",x"71",x"1e"),
   742 => (x"ff",x"1e",x"f8",x"c2"),
   743 => (x"cc",x"87",x"f3",x"d3"),
   744 => (x"c2",x"d5",x"c1",x"86"),
   745 => (x"73",x"49",x"bf",x"97"),
   746 => (x"c3",x"d5",x"c1",x"81"),
   747 => (x"c8",x"4a",x"bf",x"97"),
   748 => (x"71",x"48",x"72",x"32"),
   749 => (x"cc",x"dd",x"c1",x"80"),
   750 => (x"c4",x"d5",x"c1",x"58"),
   751 => (x"c1",x"48",x"bf",x"97"),
   752 => (x"c1",x"58",x"e0",x"dd"),
   753 => (x"02",x"bf",x"fc",x"dc"),
   754 => (x"c8",x"87",x"da",x"c2"),
   755 => (x"fc",x"c0",x"c1",x"1e"),
   756 => (x"c6",x"d6",x"c1",x"1e"),
   757 => (x"87",x"c1",x"f6",x"1e"),
   758 => (x"98",x"70",x"86",x"cc"),
   759 => (x"87",x"c5",x"c0",x"02"),
   760 => (x"d1",x"c3",x"48",x"c0"),
   761 => (x"f4",x"dc",x"c1",x"87"),
   762 => (x"48",x"72",x"4a",x"bf"),
   763 => (x"dd",x"c1",x"30",x"c4"),
   764 => (x"dd",x"c1",x"58",x"e4"),
   765 => (x"d5",x"c1",x"5a",x"dc"),
   766 => (x"49",x"bf",x"97",x"d9"),
   767 => (x"d5",x"c1",x"31",x"c8"),
   768 => (x"4b",x"bf",x"97",x"d8"),
   769 => (x"d5",x"c1",x"81",x"73"),
   770 => (x"4b",x"bf",x"97",x"da"),
   771 => (x"81",x"73",x"33",x"d0"),
   772 => (x"97",x"db",x"d5",x"c1"),
   773 => (x"33",x"d8",x"4b",x"bf"),
   774 => (x"dd",x"c1",x"81",x"73"),
   775 => (x"dd",x"c1",x"59",x"e8"),
   776 => (x"c1",x"91",x"bf",x"dc"),
   777 => (x"81",x"bf",x"c8",x"dd"),
   778 => (x"59",x"d0",x"dd",x"c1"),
   779 => (x"97",x"e1",x"d5",x"c1"),
   780 => (x"33",x"c8",x"4b",x"bf"),
   781 => (x"97",x"e0",x"d5",x"c1"),
   782 => (x"83",x"74",x"4c",x"bf"),
   783 => (x"97",x"e2",x"d5",x"c1"),
   784 => (x"34",x"d0",x"4c",x"bf"),
   785 => (x"d5",x"c1",x"83",x"74"),
   786 => (x"4c",x"bf",x"97",x"e3"),
   787 => (x"34",x"d8",x"9c",x"cf"),
   788 => (x"dd",x"c1",x"83",x"74"),
   789 => (x"8b",x"c2",x"5b",x"d4"),
   790 => (x"48",x"72",x"92",x"73"),
   791 => (x"dd",x"c1",x"80",x"71"),
   792 => (x"cf",x"c1",x"58",x"d8"),
   793 => (x"c6",x"d5",x"c1",x"87"),
   794 => (x"c8",x"49",x"bf",x"97"),
   795 => (x"c5",x"d5",x"c1",x"31"),
   796 => (x"72",x"4a",x"bf",x"97"),
   797 => (x"e4",x"dd",x"c1",x"81"),
   798 => (x"c7",x"31",x"c5",x"59"),
   799 => (x"29",x"c9",x"81",x"ff"),
   800 => (x"59",x"dc",x"dd",x"c1"),
   801 => (x"97",x"cb",x"d5",x"c1"),
   802 => (x"32",x"c8",x"4a",x"bf"),
   803 => (x"97",x"ca",x"d5",x"c1"),
   804 => (x"82",x"73",x"4b",x"bf"),
   805 => (x"5a",x"e8",x"dd",x"c1"),
   806 => (x"bf",x"dc",x"dd",x"c1"),
   807 => (x"c8",x"dd",x"c1",x"92"),
   808 => (x"dd",x"c1",x"82",x"bf"),
   809 => (x"dd",x"c1",x"5a",x"d8"),
   810 => (x"78",x"c0",x"48",x"d0"),
   811 => (x"80",x"71",x"48",x"72"),
   812 => (x"58",x"d0",x"dd",x"c1"),
   813 => (x"ea",x"f3",x"48",x"c1"),
   814 => (x"5b",x"5e",x"0e",x"87"),
   815 => (x"dc",x"c1",x"0e",x"5c"),
   816 => (x"c0",x"02",x"bf",x"fc"),
   817 => (x"66",x"cc",x"87",x"cf"),
   818 => (x"2a",x"b7",x"c7",x"4a"),
   819 => (x"c1",x"4b",x"66",x"cc"),
   820 => (x"cc",x"c0",x"9b",x"ff"),
   821 => (x"4a",x"66",x"cc",x"87"),
   822 => (x"cc",x"2a",x"b7",x"c8"),
   823 => (x"ff",x"c3",x"4b",x"66"),
   824 => (x"f4",x"d4",x"c1",x"9b"),
   825 => (x"c8",x"dd",x"c1",x"1e"),
   826 => (x"81",x"72",x"49",x"bf"),
   827 => (x"f4",x"e8",x"1e",x"71"),
   828 => (x"70",x"86",x"c8",x"87"),
   829 => (x"c5",x"c0",x"05",x"98"),
   830 => (x"c0",x"48",x"c0",x"87"),
   831 => (x"dc",x"c1",x"87",x"ea"),
   832 => (x"c0",x"02",x"bf",x"fc"),
   833 => (x"49",x"73",x"87",x"d4"),
   834 => (x"c1",x"91",x"b7",x"c4"),
   835 => (x"69",x"81",x"f4",x"d4"),
   836 => (x"ff",x"ff",x"cf",x"4c"),
   837 => (x"c0",x"9c",x"ff",x"ff"),
   838 => (x"49",x"73",x"87",x"cc"),
   839 => (x"c1",x"91",x"b7",x"c2"),
   840 => (x"9f",x"81",x"f4",x"d4"),
   841 => (x"48",x"74",x"4c",x"69"),
   842 => (x"0e",x"87",x"fa",x"f1"),
   843 => (x"5d",x"5c",x"5b",x"5e"),
   844 => (x"c0",x"86",x"f4",x"0e"),
   845 => (x"c1",x"48",x"76",x"4b"),
   846 => (x"78",x"bf",x"d0",x"dd"),
   847 => (x"dd",x"c1",x"80",x"c4"),
   848 => (x"c1",x"78",x"bf",x"d4"),
   849 => (x"02",x"bf",x"fc",x"dc"),
   850 => (x"c1",x"87",x"ca",x"c0"),
   851 => (x"49",x"bf",x"f4",x"dc"),
   852 => (x"c7",x"c0",x"31",x"c4"),
   853 => (x"d8",x"dd",x"c1",x"87"),
   854 => (x"31",x"c4",x"49",x"bf"),
   855 => (x"c0",x"59",x"a6",x"cc"),
   856 => (x"48",x"66",x"c8",x"4d"),
   857 => (x"c2",x"06",x"a8",x"c0"),
   858 => (x"49",x"75",x"87",x"f5"),
   859 => (x"99",x"71",x"99",x"cf"),
   860 => (x"87",x"db",x"c0",x"05"),
   861 => (x"1e",x"f4",x"d4",x"c1"),
   862 => (x"48",x"49",x"66",x"c8"),
   863 => (x"a6",x"cc",x"80",x"c1"),
   864 => (x"e6",x"1e",x"71",x"58"),
   865 => (x"86",x"c8",x"87",x"df"),
   866 => (x"4b",x"f4",x"d4",x"c1"),
   867 => (x"c0",x"87",x"c3",x"c0"),
   868 => (x"6b",x"97",x"83",x"e0"),
   869 => (x"02",x"99",x"71",x"49"),
   870 => (x"97",x"87",x"fb",x"c1"),
   871 => (x"e5",x"c3",x"49",x"6b"),
   872 => (x"f1",x"c1",x"02",x"a9"),
   873 => (x"cb",x"49",x"73",x"87"),
   874 => (x"49",x"69",x"97",x"81"),
   875 => (x"99",x"71",x"99",x"d8"),
   876 => (x"87",x"e2",x"c1",x"05"),
   877 => (x"ca",x"ff",x"1e",x"73"),
   878 => (x"86",x"c4",x"87",x"dc"),
   879 => (x"e4",x"c0",x"1e",x"cb"),
   880 => (x"1e",x"73",x"1e",x"66"),
   881 => (x"cc",x"87",x"d2",x"ee"),
   882 => (x"05",x"98",x"70",x"86"),
   883 => (x"73",x"87",x"c7",x"c1"),
   884 => (x"dc",x"82",x"dc",x"4a"),
   885 => (x"81",x"c4",x"49",x"66"),
   886 => (x"4a",x"73",x"79",x"6a"),
   887 => (x"66",x"dc",x"82",x"da"),
   888 => (x"9f",x"81",x"c8",x"49"),
   889 => (x"79",x"70",x"48",x"6a"),
   890 => (x"dc",x"c1",x"4c",x"71"),
   891 => (x"c0",x"02",x"bf",x"fc"),
   892 => (x"49",x"73",x"87",x"d2"),
   893 => (x"69",x"9f",x"81",x"d4"),
   894 => (x"ff",x"ff",x"c0",x"49"),
   895 => (x"d0",x"4a",x"71",x"99"),
   896 => (x"87",x"c2",x"c0",x"32"),
   897 => (x"48",x"72",x"4a",x"c0"),
   898 => (x"7c",x"70",x"80",x"6c"),
   899 => (x"c0",x"48",x"66",x"dc"),
   900 => (x"c1",x"48",x"c1",x"78"),
   901 => (x"85",x"c1",x"87",x"c0"),
   902 => (x"04",x"ad",x"66",x"c8"),
   903 => (x"c1",x"87",x"cb",x"fd"),
   904 => (x"02",x"bf",x"fc",x"dc"),
   905 => (x"6e",x"87",x"ed",x"c0"),
   906 => (x"87",x"cd",x"fa",x"1e"),
   907 => (x"a6",x"c4",x"86",x"c4"),
   908 => (x"cf",x"49",x"6e",x"58"),
   909 => (x"f8",x"ff",x"ff",x"ff"),
   910 => (x"c0",x"02",x"a9",x"99"),
   911 => (x"49",x"6e",x"87",x"d6"),
   912 => (x"dc",x"c1",x"89",x"c2"),
   913 => (x"c1",x"91",x"bf",x"f4"),
   914 => (x"48",x"bf",x"cc",x"dd"),
   915 => (x"a6",x"c8",x"80",x"71"),
   916 => (x"87",x"cb",x"fc",x"58"),
   917 => (x"8e",x"f4",x"48",x"c0"),
   918 => (x"0e",x"87",x"c8",x"ed"),
   919 => (x"c8",x"0e",x"5b",x"5e"),
   920 => (x"c1",x"49",x"bf",x"66"),
   921 => (x"09",x"66",x"c8",x"81"),
   922 => (x"dc",x"c1",x"09",x"79"),
   923 => (x"71",x"99",x"bf",x"f8"),
   924 => (x"d0",x"c0",x"05",x"99"),
   925 => (x"4b",x"66",x"c8",x"87"),
   926 => (x"1e",x"6b",x"83",x"c8"),
   927 => (x"c4",x"87",x"fa",x"f8"),
   928 => (x"71",x"49",x"70",x"86"),
   929 => (x"ec",x"48",x"c1",x"7b"),
   930 => (x"5e",x"0e",x"87",x"dd"),
   931 => (x"cc",x"dd",x"c1",x"0e"),
   932 => (x"66",x"c4",x"49",x"bf"),
   933 => (x"6a",x"82",x"c8",x"4a"),
   934 => (x"c1",x"8a",x"c2",x"4a"),
   935 => (x"92",x"bf",x"f4",x"dc"),
   936 => (x"dc",x"c1",x"81",x"72"),
   937 => (x"c4",x"4a",x"bf",x"f8"),
   938 => (x"72",x"9a",x"bf",x"66"),
   939 => (x"1e",x"66",x"c8",x"81"),
   940 => (x"f0",x"e1",x"1e",x"71"),
   941 => (x"70",x"86",x"c8",x"87"),
   942 => (x"c5",x"c0",x"05",x"98"),
   943 => (x"c0",x"48",x"c0",x"87"),
   944 => (x"48",x"c1",x"87",x"c2"),
   945 => (x"0e",x"87",x"e2",x"eb"),
   946 => (x"0e",x"5c",x"5b",x"5e"),
   947 => (x"c1",x"1e",x"66",x"cc"),
   948 => (x"f9",x"1e",x"ec",x"dd"),
   949 => (x"86",x"c8",x"87",x"d5"),
   950 => (x"c1",x"02",x"98",x"70"),
   951 => (x"dd",x"c1",x"87",x"d4"),
   952 => (x"c7",x"49",x"bf",x"f0"),
   953 => (x"29",x"c9",x"81",x"ff"),
   954 => (x"4b",x"c0",x"4c",x"71"),
   955 => (x"1e",x"c9",x"fd",x"c0"),
   956 => (x"87",x"e2",x"c5",x"ff"),
   957 => (x"b7",x"c0",x"86",x"c4"),
   958 => (x"c7",x"c1",x"06",x"ac"),
   959 => (x"1e",x"66",x"d0",x"87"),
   960 => (x"1e",x"ec",x"dd",x"c1"),
   961 => (x"c8",x"87",x"c3",x"fe"),
   962 => (x"05",x"98",x"70",x"86"),
   963 => (x"c0",x"87",x"c5",x"c0"),
   964 => (x"87",x"f2",x"c0",x"48"),
   965 => (x"1e",x"ec",x"dd",x"c1"),
   966 => (x"c4",x"87",x"c0",x"fd"),
   967 => (x"48",x"66",x"d0",x"86"),
   968 => (x"d4",x"80",x"c0",x"c8"),
   969 => (x"83",x"c1",x"58",x"a6"),
   970 => (x"04",x"ab",x"b7",x"74"),
   971 => (x"c0",x"87",x"ce",x"ff"),
   972 => (x"66",x"cc",x"87",x"d2"),
   973 => (x"e2",x"fd",x"c0",x"1e"),
   974 => (x"d5",x"c5",x"ff",x"1e"),
   975 => (x"c0",x"86",x"c8",x"87"),
   976 => (x"87",x"c2",x"c0",x"48"),
   977 => (x"dc",x"e9",x"48",x"c1"),
   978 => (x"65",x"70",x"4f",x"87"),
   979 => (x"20",x"64",x"65",x"6e"),
   980 => (x"65",x"6c",x"69",x"66"),
   981 => (x"6f",x"6c",x"20",x"2c"),
   982 => (x"6e",x"69",x"64",x"61"),
   983 => (x"2e",x"2e",x"2e",x"67"),
   984 => (x"61",x"43",x"00",x"0a"),
   985 => (x"20",x"74",x"27",x"6e"),
   986 => (x"6e",x"65",x"70",x"6f"),
   987 => (x"0a",x"73",x"25",x"20"),
   988 => (x"61",x"65",x"52",x"00"),
   989 => (x"66",x"6f",x"20",x"64"),
   990 => (x"52",x"42",x"4d",x"20"),
   991 => (x"69",x"61",x"66",x"20"),
   992 => (x"0a",x"64",x"65",x"6c"),
   993 => (x"20",x"6f",x"4e",x"00"),
   994 => (x"74",x"72",x"61",x"70"),
   995 => (x"6f",x"69",x"74",x"69"),
   996 => (x"69",x"73",x"20",x"6e"),
   997 => (x"74",x"61",x"6e",x"67"),
   998 => (x"20",x"65",x"72",x"75"),
   999 => (x"6e",x"75",x"6f",x"66"),
  1000 => (x"4d",x"00",x"0a",x"64"),
  1001 => (x"69",x"73",x"52",x"42"),
  1002 => (x"20",x"3a",x"65",x"7a"),
  1003 => (x"20",x"2c",x"64",x"25"),
  1004 => (x"74",x"72",x"61",x"70"),
  1005 => (x"6f",x"69",x"74",x"69"),
  1006 => (x"7a",x"69",x"73",x"6e"),
  1007 => (x"25",x"20",x"3a",x"65"),
  1008 => (x"6f",x"20",x"2c",x"64"),
  1009 => (x"65",x"73",x"66",x"66"),
  1010 => (x"66",x"6f",x"20",x"74"),
  1011 => (x"67",x"69",x"73",x"20"),
  1012 => (x"64",x"25",x"20",x"3a"),
  1013 => (x"69",x"73",x"20",x"2c"),
  1014 => (x"78",x"30",x"20",x"67"),
  1015 => (x"00",x"0a",x"78",x"25"),
  1016 => (x"64",x"61",x"65",x"52"),
  1017 => (x"20",x"67",x"6e",x"69"),
  1018 => (x"74",x"6f",x"6f",x"62"),
  1019 => (x"63",x"65",x"73",x"20"),
  1020 => (x"20",x"72",x"6f",x"74"),
  1021 => (x"00",x"0a",x"64",x"25"),
  1022 => (x"64",x"61",x"65",x"52"),
  1023 => (x"6f",x"6f",x"62",x"20"),
  1024 => (x"65",x"73",x"20",x"74"),
  1025 => (x"72",x"6f",x"74",x"63"),
  1026 => (x"6f",x"72",x"66",x"20"),
  1027 => (x"69",x"66",x"20",x"6d"),
  1028 => (x"20",x"74",x"73",x"72"),
  1029 => (x"74",x"72",x"61",x"70"),
  1030 => (x"6f",x"69",x"74",x"69"),
  1031 => (x"55",x"00",x"0a",x"6e"),
  1032 => (x"70",x"75",x"73",x"6e"),
  1033 => (x"74",x"72",x"6f",x"70"),
  1034 => (x"70",x"20",x"64",x"65"),
  1035 => (x"69",x"74",x"72",x"61"),
  1036 => (x"6e",x"6f",x"69",x"74"),
  1037 => (x"70",x"79",x"74",x"20"),
  1038 => (x"00",x"0d",x"21",x"65"),
  1039 => (x"33",x"54",x"41",x"46"),
  1040 => (x"20",x"20",x"20",x"32"),
  1041 => (x"61",x"65",x"52",x"00"),
  1042 => (x"67",x"6e",x"69",x"64"),
  1043 => (x"52",x"42",x"4d",x"20"),
  1044 => (x"42",x"4d",x"00",x"0a"),
  1045 => (x"75",x"73",x"20",x"52"),
  1046 => (x"73",x"65",x"63",x"63"),
  1047 => (x"6c",x"75",x"66",x"73"),
  1048 => (x"72",x"20",x"79",x"6c"),
  1049 => (x"0a",x"64",x"61",x"65"),
  1050 => (x"54",x"41",x"46",x"00"),
  1051 => (x"20",x"20",x"36",x"31"),
  1052 => (x"41",x"46",x"00",x"20"),
  1053 => (x"20",x"32",x"33",x"54"),
  1054 => (x"50",x"00",x"20",x"20"),
  1055 => (x"69",x"74",x"72",x"61"),
  1056 => (x"6e",x"6f",x"69",x"74"),
  1057 => (x"6e",x"75",x"6f",x"63"),
  1058 => (x"64",x"25",x"20",x"74"),
  1059 => (x"75",x"48",x"00",x"0a"),
  1060 => (x"6e",x"69",x"74",x"6e"),
  1061 => (x"6f",x"66",x"20",x"67"),
  1062 => (x"69",x"66",x"20",x"72"),
  1063 => (x"79",x"73",x"65",x"6c"),
  1064 => (x"6d",x"65",x"74",x"73"),
  1065 => (x"41",x"46",x"00",x"0a"),
  1066 => (x"20",x"32",x"33",x"54"),
  1067 => (x"46",x"00",x"20",x"20"),
  1068 => (x"36",x"31",x"54",x"41"),
  1069 => (x"00",x"20",x"20",x"20"),
  1070 => (x"73",x"75",x"6c",x"43"),
  1071 => (x"20",x"72",x"65",x"74"),
  1072 => (x"65",x"7a",x"69",x"73"),
  1073 => (x"64",x"25",x"20",x"3a"),
  1074 => (x"6c",x"43",x"20",x"2c"),
  1075 => (x"65",x"74",x"73",x"75"),
  1076 => (x"61",x"6d",x"20",x"72"),
  1077 => (x"20",x"2c",x"6b",x"73"),
  1078 => (x"00",x"0a",x"64",x"25"),
  1079 => (x"c4",x"0e",x"5e",x"0e"),
  1080 => (x"29",x"d8",x"49",x"66"),
  1081 => (x"c4",x"99",x"ff",x"c3"),
  1082 => (x"2a",x"c8",x"4a",x"66"),
  1083 => (x"9a",x"c0",x"fc",x"cf"),
  1084 => (x"66",x"c4",x"b1",x"72"),
  1085 => (x"c0",x"32",x"c8",x"4a"),
  1086 => (x"c0",x"c0",x"f0",x"ff"),
  1087 => (x"c4",x"b1",x"72",x"9a"),
  1088 => (x"32",x"d8",x"4a",x"66"),
  1089 => (x"c0",x"c0",x"c0",x"ff"),
  1090 => (x"b1",x"72",x"9a",x"c0"),
  1091 => (x"87",x"c6",x"48",x"71"),
  1092 => (x"4c",x"26",x"4d",x"26"),
  1093 => (x"4f",x"26",x"4b",x"26"),
  1094 => (x"c4",x"0e",x"5e",x"0e"),
  1095 => (x"2a",x"c8",x"4a",x"66"),
  1096 => (x"cf",x"9a",x"ff",x"c3"),
  1097 => (x"c4",x"9a",x"ff",x"ff"),
  1098 => (x"31",x"c8",x"49",x"66"),
  1099 => (x"99",x"c0",x"fc",x"cf"),
  1100 => (x"ff",x"cf",x"b1",x"72"),
  1101 => (x"48",x"71",x"99",x"ff"),
  1102 => (x"0e",x"87",x"db",x"ff"),
  1103 => (x"66",x"c4",x"0e",x"5e"),
  1104 => (x"cf",x"29",x"d0",x"49"),
  1105 => (x"c4",x"99",x"ff",x"ff"),
  1106 => (x"32",x"d0",x"4a",x"66"),
  1107 => (x"9a",x"c0",x"c0",x"f0"),
  1108 => (x"48",x"71",x"b1",x"72"),
  1109 => (x"1e",x"87",x"ff",x"fe"),
  1110 => (x"c0",x"d0",x"1e",x"73"),
  1111 => (x"4b",x"c0",x"c0",x"c0"),
  1112 => (x"87",x"fe",x"0f",x"73"),
  1113 => (x"4d",x"26",x"87",x"c4"),
  1114 => (x"4b",x"26",x"4c",x"26"),
  1115 => (x"c8",x"1e",x"4f",x"26"),
  1116 => (x"df",x"c3",x"49",x"66"),
  1117 => (x"89",x"f7",x"c0",x"99"),
  1118 => (x"03",x"a9",x"b7",x"c0"),
  1119 => (x"e7",x"c0",x"87",x"c3"),
  1120 => (x"48",x"66",x"c4",x"81"),
  1121 => (x"a6",x"c8",x"30",x"c4"),
  1122 => (x"48",x"66",x"c4",x"58"),
  1123 => (x"a6",x"c8",x"b0",x"71"),
  1124 => (x"48",x"66",x"c4",x"58"),
  1125 => (x"0e",x"87",x"d5",x"ff"),
  1126 => (x"0e",x"5c",x"5b",x"5e"),
  1127 => (x"c0",x"c0",x"c0",x"d0"),
  1128 => (x"dd",x"c1",x"4c",x"c0"),
  1129 => (x"c1",x"48",x"bf",x"f8"),
  1130 => (x"fc",x"dd",x"c1",x"80"),
  1131 => (x"66",x"cc",x"97",x"58"),
  1132 => (x"81",x"c0",x"fe",x"49"),
  1133 => (x"a9",x"d3",x"c1",x"b9"),
  1134 => (x"87",x"e1",x"c0",x"05"),
  1135 => (x"48",x"f8",x"dd",x"c1"),
  1136 => (x"dd",x"c1",x"78",x"c0"),
  1137 => (x"78",x"c0",x"48",x"fc"),
  1138 => (x"48",x"c4",x"de",x"c1"),
  1139 => (x"de",x"c1",x"78",x"c0"),
  1140 => (x"78",x"c0",x"48",x"c8"),
  1141 => (x"c1",x"48",x"c0",x"ff"),
  1142 => (x"ee",x"c7",x"78",x"d3"),
  1143 => (x"f8",x"dd",x"c1",x"87"),
  1144 => (x"a8",x"c1",x"48",x"bf"),
  1145 => (x"87",x"c8",x"c1",x"05"),
  1146 => (x"c1",x"48",x"c0",x"ff"),
  1147 => (x"cc",x"97",x"78",x"f4"),
  1148 => (x"c0",x"fe",x"49",x"66"),
  1149 => (x"1e",x"71",x"b9",x"81"),
  1150 => (x"bf",x"c8",x"de",x"c1"),
  1151 => (x"87",x"ee",x"fd",x"1e"),
  1152 => (x"de",x"c1",x"86",x"c8"),
  1153 => (x"de",x"c1",x"58",x"cc"),
  1154 => (x"c3",x"4a",x"bf",x"c8"),
  1155 => (x"c6",x"06",x"aa",x"b7"),
  1156 => (x"72",x"48",x"ca",x"87"),
  1157 => (x"72",x"4a",x"70",x"88"),
  1158 => (x"71",x"81",x"c1",x"49"),
  1159 => (x"c1",x"30",x"c1",x"48"),
  1160 => (x"72",x"58",x"c4",x"de"),
  1161 => (x"80",x"f0",x"c0",x"48"),
  1162 => (x"78",x"08",x"c0",x"ff"),
  1163 => (x"87",x"db",x"c6",x"08"),
  1164 => (x"bf",x"c8",x"de",x"c1"),
  1165 => (x"a8",x"b7",x"c9",x"48"),
  1166 => (x"87",x"cf",x"c6",x"01"),
  1167 => (x"bf",x"c8",x"de",x"c1"),
  1168 => (x"a8",x"b7",x"c0",x"48"),
  1169 => (x"87",x"c3",x"c6",x"06"),
  1170 => (x"bf",x"c8",x"de",x"c1"),
  1171 => (x"80",x"f0",x"c0",x"48"),
  1172 => (x"78",x"08",x"c0",x"ff"),
  1173 => (x"f8",x"dd",x"c1",x"08"),
  1174 => (x"b7",x"c3",x"48",x"bf"),
  1175 => (x"87",x"db",x"01",x"a8"),
  1176 => (x"49",x"66",x"cc",x"97"),
  1177 => (x"b9",x"81",x"c0",x"fe"),
  1178 => (x"de",x"c1",x"1e",x"71"),
  1179 => (x"fb",x"1e",x"bf",x"c4"),
  1180 => (x"86",x"c8",x"87",x"fc"),
  1181 => (x"58",x"c8",x"de",x"c1"),
  1182 => (x"c1",x"87",x"d0",x"c5"),
  1183 => (x"49",x"bf",x"c0",x"de"),
  1184 => (x"dd",x"c1",x"81",x"c3"),
  1185 => (x"a9",x"b7",x"bf",x"f8"),
  1186 => (x"87",x"e1",x"c0",x"04"),
  1187 => (x"49",x"66",x"cc",x"97"),
  1188 => (x"b9",x"81",x"c0",x"fe"),
  1189 => (x"dd",x"c1",x"1e",x"71"),
  1190 => (x"fb",x"1e",x"bf",x"fc"),
  1191 => (x"86",x"c8",x"87",x"d0"),
  1192 => (x"58",x"c0",x"de",x"c1"),
  1193 => (x"48",x"cc",x"de",x"c1"),
  1194 => (x"de",x"c4",x"78",x"c1"),
  1195 => (x"c8",x"de",x"c1",x"87"),
  1196 => (x"b7",x"c0",x"48",x"bf"),
  1197 => (x"db",x"c2",x"06",x"a8"),
  1198 => (x"c8",x"de",x"c1",x"87"),
  1199 => (x"b7",x"c3",x"48",x"bf"),
  1200 => (x"cf",x"c2",x"01",x"a8"),
  1201 => (x"c4",x"de",x"c1",x"87"),
  1202 => (x"31",x"c1",x"49",x"bf"),
  1203 => (x"f8",x"dd",x"c1",x"81"),
  1204 => (x"04",x"a9",x"b7",x"bf"),
  1205 => (x"97",x"87",x"df",x"c1"),
  1206 => (x"fe",x"49",x"66",x"cc"),
  1207 => (x"71",x"b9",x"81",x"c0"),
  1208 => (x"d0",x"de",x"c1",x"1e"),
  1209 => (x"c5",x"fa",x"1e",x"bf"),
  1210 => (x"c1",x"86",x"c8",x"87"),
  1211 => (x"c1",x"58",x"d4",x"de"),
  1212 => (x"49",x"bf",x"cc",x"de"),
  1213 => (x"de",x"c1",x"89",x"c1"),
  1214 => (x"b7",x"c0",x"59",x"d0"),
  1215 => (x"ca",x"c3",x"03",x"a9"),
  1216 => (x"fc",x"dd",x"c1",x"87"),
  1217 => (x"de",x"c1",x"49",x"bf"),
  1218 => (x"51",x"bf",x"97",x"d0"),
  1219 => (x"c1",x"98",x"ff",x"c3"),
  1220 => (x"49",x"bf",x"fc",x"dd"),
  1221 => (x"de",x"c1",x"81",x"c1"),
  1222 => (x"de",x"c1",x"59",x"c0"),
  1223 => (x"a9",x"b7",x"bf",x"d4"),
  1224 => (x"87",x"c9",x"c0",x"06"),
  1225 => (x"48",x"d4",x"de",x"c1"),
  1226 => (x"bf",x"fc",x"dd",x"c1"),
  1227 => (x"cc",x"de",x"c1",x"78"),
  1228 => (x"c2",x"78",x"c1",x"48"),
  1229 => (x"de",x"c1",x"87",x"d5"),
  1230 => (x"c2",x"05",x"bf",x"cc"),
  1231 => (x"de",x"c1",x"87",x"cd"),
  1232 => (x"c4",x"49",x"bf",x"d0"),
  1233 => (x"d4",x"de",x"c1",x"31"),
  1234 => (x"fc",x"dd",x"c1",x"59"),
  1235 => (x"79",x"97",x"09",x"bf"),
  1236 => (x"87",x"f7",x"c1",x"09"),
  1237 => (x"bf",x"c8",x"de",x"c1"),
  1238 => (x"a8",x"b7",x"c7",x"48"),
  1239 => (x"87",x"de",x"c1",x"04"),
  1240 => (x"f4",x"fe",x"4b",x"c0"),
  1241 => (x"c1",x"78",x"c1",x"48"),
  1242 => (x"1e",x"bf",x"d4",x"de"),
  1243 => (x"d3",x"c1",x"1e",x"74"),
  1244 => (x"f4",x"fe",x"1e",x"ea"),
  1245 => (x"86",x"cc",x"87",x"dc"),
  1246 => (x"5c",x"c0",x"de",x"c1"),
  1247 => (x"bf",x"fc",x"dd",x"c1"),
  1248 => (x"d4",x"de",x"c1",x"48"),
  1249 => (x"03",x"a8",x"b7",x"bf"),
  1250 => (x"c1",x"87",x"db",x"c0"),
  1251 => (x"bf",x"bf",x"fc",x"dd"),
  1252 => (x"fc",x"dd",x"c1",x"83"),
  1253 => (x"81",x"c4",x"49",x"bf"),
  1254 => (x"59",x"c0",x"de",x"c1"),
  1255 => (x"bf",x"d4",x"de",x"c1"),
  1256 => (x"ff",x"04",x"a9",x"b7"),
  1257 => (x"1e",x"73",x"87",x"e5"),
  1258 => (x"1e",x"c9",x"d4",x"c1"),
  1259 => (x"87",x"e2",x"f3",x"fe"),
  1260 => (x"c0",x"ff",x"86",x"c8"),
  1261 => (x"78",x"c2",x"c1",x"48"),
  1262 => (x"c0",x"87",x"dc",x"f6"),
  1263 => (x"de",x"c1",x"87",x"cd"),
  1264 => (x"c0",x"48",x"bf",x"c8"),
  1265 => (x"c0",x"ff",x"80",x"f0"),
  1266 => (x"f6",x"08",x"78",x"08"),
  1267 => (x"5e",x"0e",x"87",x"da"),
  1268 => (x"0e",x"5d",x"5c",x"5b"),
  1269 => (x"1e",x"ec",x"d2",x"c1"),
  1270 => (x"87",x"fa",x"f1",x"fe"),
  1271 => (x"c3",x"ff",x"86",x"c4"),
  1272 => (x"98",x"70",x"87",x"c9"),
  1273 => (x"87",x"cf",x"c0",x"02"),
  1274 => (x"87",x"ff",x"d6",x"ff"),
  1275 => (x"c0",x"02",x"98",x"70"),
  1276 => (x"49",x"c1",x"87",x"c5"),
  1277 => (x"c0",x"87",x"c2",x"c0"),
  1278 => (x"c1",x"4d",x"71",x"49"),
  1279 => (x"fe",x"1e",x"c2",x"d3"),
  1280 => (x"c4",x"87",x"d3",x"f1"),
  1281 => (x"d4",x"de",x"c1",x"86"),
  1282 => (x"c0",x"78",x"c0",x"48"),
  1283 => (x"f0",x"fe",x"1e",x"ee"),
  1284 => (x"86",x"c4",x"87",x"ea"),
  1285 => (x"ff",x"c8",x"f4",x"c3"),
  1286 => (x"bf",x"c0",x"ff",x"4a"),
  1287 => (x"c8",x"49",x"74",x"4c"),
  1288 => (x"99",x"71",x"99",x"c0"),
  1289 => (x"87",x"cc",x"c1",x"02"),
  1290 => (x"ff",x"c3",x"4b",x"74"),
  1291 => (x"05",x"ab",x"db",x"9b"),
  1292 => (x"75",x"87",x"f5",x"c0"),
  1293 => (x"e5",x"c0",x"02",x"9d"),
  1294 => (x"c0",x"c0",x"d0",x"87"),
  1295 => (x"c1",x"1e",x"c0",x"c0"),
  1296 => (x"ea",x"1e",x"d0",x"d2"),
  1297 => (x"86",x"c8",x"87",x"c1"),
  1298 => (x"c0",x"02",x"98",x"70"),
  1299 => (x"d2",x"c1",x"87",x"d0"),
  1300 => (x"f0",x"fe",x"1e",x"c4"),
  1301 => (x"86",x"c4",x"87",x"c0"),
  1302 => (x"c0",x"87",x"fc",x"f3"),
  1303 => (x"d2",x"c1",x"87",x"ca"),
  1304 => (x"ef",x"fe",x"1e",x"dc"),
  1305 => (x"86",x"c4",x"87",x"f0"),
  1306 => (x"ea",x"f4",x"1e",x"73"),
  1307 => (x"c3",x"86",x"c4",x"87"),
  1308 => (x"4a",x"c0",x"c9",x"f4"),
  1309 => (x"8a",x"c1",x"49",x"72"),
  1310 => (x"fe",x"05",x"99",x"71"),
  1311 => (x"ca",x"fe",x"87",x"db"),
  1312 => (x"87",x"e2",x"f3",x"87"),
  1313 => (x"74",x"6f",x"6f",x"42"),
  1314 => (x"2e",x"67",x"6e",x"69"),
  1315 => (x"00",x"0a",x"2e",x"2e"),
  1316 => (x"54",x"4f",x"4f",x"42"),
  1317 => (x"20",x"32",x"33",x"38"),
  1318 => (x"00",x"4e",x"49",x"42"),
  1319 => (x"62",x"20",x"44",x"53"),
  1320 => (x"20",x"74",x"6f",x"6f"),
  1321 => (x"6c",x"69",x"61",x"66"),
  1322 => (x"00",x"0a",x"64",x"65"),
  1323 => (x"74",x"69",x"6e",x"49"),
  1324 => (x"69",x"6c",x"61",x"69"),
  1325 => (x"67",x"6e",x"69",x"7a"),
  1326 => (x"20",x"44",x"53",x"20"),
  1327 => (x"64",x"72",x"61",x"63"),
  1328 => (x"53",x"52",x"00",x"0a"),
  1329 => (x"20",x"32",x"33",x"32"),
  1330 => (x"74",x"6f",x"6f",x"62"),
  1331 => (x"70",x"20",x"2d",x"20"),
  1332 => (x"73",x"73",x"65",x"72"),
  1333 => (x"43",x"53",x"45",x"20"),
  1334 => (x"20",x"6f",x"74",x"20"),
  1335 => (x"74",x"6f",x"6f",x"62"),
  1336 => (x"6f",x"72",x"66",x"20"),
  1337 => (x"44",x"53",x"20",x"6d"),
  1338 => (x"68",x"43",x"00",x"2e"),
  1339 => (x"73",x"6b",x"63",x"65"),
  1340 => (x"69",x"6d",x"6d",x"75"),
  1341 => (x"66",x"20",x"67",x"6e"),
  1342 => (x"20",x"6d",x"6f",x"72"),
  1343 => (x"74",x"20",x"64",x"25"),
  1344 => (x"64",x"25",x"20",x"6f"),
  1345 => (x"20",x"2e",x"2e",x"2e"),
  1346 => (x"0a",x"64",x"25",x"00"),
  1347 => (x"0a",x"64",x"25",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
