
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"2c",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"29"),
    10 => (x"87",x"fd",x"00",x"4f"),
    11 => (x"d0",x"de",x"c1",x"4f"),
    12 => (x"c0",x"c0",x"c1",x"4e"),
    13 => (x"d0",x"de",x"c1",x"86"),
    14 => (x"f8",x"d3",x"c1",x"49"),
    15 => (x"89",x"d0",x"89",x"48"),
    16 => (x"40",x"40",x"c0",x"03"),
    17 => (x"87",x"f6",x"40",x"40"),
    18 => (x"c0",x"05",x"81",x"d0"),
    19 => (x"05",x"89",x"c1",x"50"),
    20 => (x"d3",x"c1",x"87",x"f9"),
    21 => (x"d3",x"c1",x"4d",x"f8"),
    22 => (x"ad",x"74",x"4c",x"f8"),
    23 => (x"24",x"87",x"c4",x"02"),
    24 => (x"d6",x"87",x"f7",x"0f"),
    25 => (x"d3",x"c1",x"87",x"f9"),
    26 => (x"d3",x"c1",x"4d",x"f8"),
    27 => (x"ad",x"74",x"4c",x"f8"),
    28 => (x"c4",x"87",x"c6",x"02"),
    29 => (x"f5",x"0f",x"6c",x"8c"),
    30 => (x"87",x"fd",x"00",x"87"),
    31 => (x"74",x"1e",x"73",x"1e"),
    32 => (x"d0",x"1e",x"75",x"1e"),
    33 => (x"d3",x"c1",x"4a",x"66"),
    34 => (x"f0",x"c3",x"4b",x"f8"),
    35 => (x"72",x"4c",x"c0",x"4d"),
    36 => (x"87",x"c6",x"05",x"9a"),
    37 => (x"c0",x"53",x"f0",x"c0"),
    38 => (x"9a",x"72",x"87",x"eb"),
    39 => (x"87",x"e5",x"c0",x"02"),
    40 => (x"49",x"72",x"1e",x"72"),
    41 => (x"c9",x"4a",x"66",x"d8"),
    42 => (x"4a",x"26",x"87",x"d1"),
    43 => (x"11",x"49",x"a1",x"75"),
    44 => (x"72",x"1e",x"71",x"53"),
    45 => (x"4a",x"66",x"d8",x"49"),
    46 => (x"70",x"87",x"c0",x"c9"),
    47 => (x"72",x"49",x"26",x"4a"),
    48 => (x"db",x"ff",x"05",x"9a"),
    49 => (x"f8",x"d3",x"c1",x"87"),
    50 => (x"87",x"da",x"02",x"ab"),
    51 => (x"dc",x"4d",x"66",x"d8"),
    52 => (x"8b",x"c1",x"1e",x"66"),
    53 => (x"71",x"49",x"6b",x"97"),
    54 => (x"c8",x"0f",x"75",x"1e"),
    55 => (x"c1",x"84",x"c1",x"86"),
    56 => (x"05",x"ab",x"f8",x"d3"),
    57 => (x"48",x"74",x"87",x"e9"),
    58 => (x"4c",x"26",x"4d",x"26"),
    59 => (x"4f",x"26",x"4b",x"26"),
    60 => (x"33",x"32",x"31",x"30"),
    61 => (x"37",x"36",x"35",x"34"),
    62 => (x"42",x"41",x"39",x"38"),
    63 => (x"46",x"45",x"44",x"43"),
    64 => (x"1e",x"73",x"1e",x"00"),
    65 => (x"1e",x"75",x"1e",x"74"),
    66 => (x"ff",x"4c",x"66",x"d0"),
    67 => (x"73",x"4b",x"14",x"4d"),
    68 => (x"87",x"d8",x"02",x"9b"),
    69 => (x"66",x"d8",x"85",x"c1"),
    70 => (x"dc",x"1e",x"73",x"1e"),
    71 => (x"86",x"c8",x"0f",x"66"),
    72 => (x"c7",x"05",x"a8",x"73"),
    73 => (x"73",x"4b",x"14",x"87"),
    74 => (x"87",x"e8",x"05",x"9b"),
    75 => (x"4d",x"26",x"48",x"75"),
    76 => (x"4b",x"26",x"4c",x"26"),
    77 => (x"73",x"1e",x"4f",x"26"),
    78 => (x"75",x"1e",x"74",x"1e"),
    79 => (x"c0",x"86",x"f4",x"1e"),
    80 => (x"c0",x"4c",x"66",x"e4"),
    81 => (x"48",x"a6",x"c4",x"4d"),
    82 => (x"66",x"dc",x"78",x"c0"),
    83 => (x"dc",x"4b",x"bf",x"97"),
    84 => (x"80",x"c1",x"48",x"66"),
    85 => (x"58",x"a6",x"e0",x"c0"),
    86 => (x"c4",x"02",x"9b",x"73"),
    87 => (x"66",x"c4",x"87",x"f9"),
    88 => (x"87",x"c8",x"c4",x"02"),
    89 => (x"c0",x"48",x"a6",x"c8"),
    90 => (x"c0",x"80",x"fc",x"78"),
    91 => (x"c0",x"49",x"73",x"78"),
    92 => (x"c1",x"02",x"ab",x"f0"),
    93 => (x"e3",x"c1",x"87",x"e5"),
    94 => (x"e6",x"c1",x"02",x"a9"),
    95 => (x"a9",x"e4",x"c1",x"87"),
    96 => (x"87",x"e2",x"c0",x"02"),
    97 => (x"02",x"a9",x"ec",x"c1"),
    98 => (x"c1",x"87",x"d0",x"c1"),
    99 => (x"dd",x"02",x"a9",x"f0"),
   100 => (x"a9",x"f3",x"c1",x"87"),
   101 => (x"c1",x"87",x"df",x"02"),
   102 => (x"c9",x"02",x"a9",x"f5"),
   103 => (x"a9",x"f8",x"c1",x"87"),
   104 => (x"c1",x"87",x"cb",x"02"),
   105 => (x"a6",x"c8",x"87",x"db"),
   106 => (x"c1",x"78",x"ca",x"48"),
   107 => (x"a6",x"c8",x"87",x"f0"),
   108 => (x"c1",x"78",x"d0",x"48"),
   109 => (x"e8",x"c0",x"87",x"e8"),
   110 => (x"1e",x"74",x"1e",x"66"),
   111 => (x"48",x"66",x"e8",x"c0"),
   112 => (x"ec",x"c0",x"80",x"c4"),
   113 => (x"e8",x"c0",x"58",x"a6"),
   114 => (x"89",x"c4",x"49",x"66"),
   115 => (x"f0",x"fc",x"1e",x"69"),
   116 => (x"70",x"86",x"cc",x"87"),
   117 => (x"4d",x"a5",x"71",x"49"),
   118 => (x"c4",x"87",x"c3",x"c1"),
   119 => (x"78",x"c1",x"48",x"a6"),
   120 => (x"c0",x"87",x"fb",x"c0"),
   121 => (x"c0",x"1e",x"66",x"e8"),
   122 => (x"c4",x"48",x"66",x"e4"),
   123 => (x"a6",x"e8",x"c0",x"80"),
   124 => (x"66",x"e4",x"c0",x"58"),
   125 => (x"69",x"89",x"c4",x"49"),
   126 => (x"c8",x"0f",x"74",x"1e"),
   127 => (x"dd",x"85",x"c1",x"86"),
   128 => (x"ab",x"e5",x"c0",x"87"),
   129 => (x"c0",x"87",x"cb",x"02"),
   130 => (x"c0",x"1e",x"66",x"e8"),
   131 => (x"0f",x"74",x"1e",x"e5"),
   132 => (x"e8",x"c0",x"86",x"c8"),
   133 => (x"1e",x"73",x"1e",x"66"),
   134 => (x"86",x"c8",x"0f",x"74"),
   135 => (x"66",x"c8",x"85",x"c1"),
   136 => (x"87",x"df",x"c1",x"02"),
   137 => (x"48",x"66",x"e0",x"c0"),
   138 => (x"e4",x"c0",x"80",x"c4"),
   139 => (x"e0",x"c0",x"58",x"a6"),
   140 => (x"89",x"c4",x"49",x"66"),
   141 => (x"e4",x"c1",x"7e",x"69"),
   142 => (x"87",x"d8",x"05",x"ab"),
   143 => (x"b7",x"c0",x"48",x"6e"),
   144 => (x"87",x"d0",x"03",x"a8"),
   145 => (x"c1",x"1e",x"ed",x"c0"),
   146 => (x"86",x"c4",x"87",x"ec"),
   147 => (x"08",x"c0",x"48",x"6e"),
   148 => (x"58",x"a6",x"c4",x"88"),
   149 => (x"1e",x"66",x"e8",x"c0"),
   150 => (x"66",x"d0",x"1e",x"74"),
   151 => (x"1e",x"66",x"cc",x"1e"),
   152 => (x"d0",x"87",x"d9",x"f8"),
   153 => (x"71",x"49",x"70",x"86"),
   154 => (x"87",x"d7",x"4d",x"a5"),
   155 => (x"05",x"ab",x"e5",x"c0"),
   156 => (x"a6",x"c4",x"87",x"c7"),
   157 => (x"ca",x"78",x"c1",x"48"),
   158 => (x"66",x"e8",x"c0",x"87"),
   159 => (x"74",x"1e",x"73",x"1e"),
   160 => (x"dc",x"86",x"c8",x"0f"),
   161 => (x"4b",x"bf",x"97",x"66"),
   162 => (x"c1",x"48",x"66",x"dc"),
   163 => (x"a6",x"e0",x"c0",x"80"),
   164 => (x"05",x"9b",x"73",x"58"),
   165 => (x"75",x"87",x"c7",x"fb"),
   166 => (x"26",x"8e",x"f4",x"48"),
   167 => (x"26",x"4c",x"26",x"4d"),
   168 => (x"1e",x"4f",x"26",x"4b"),
   169 => (x"f6",x"ca",x"1e",x"c0"),
   170 => (x"1e",x"a6",x"d0",x"1e"),
   171 => (x"fa",x"1e",x"66",x"d0"),
   172 => (x"86",x"d0",x"87",x"c4"),
   173 => (x"fc",x"1e",x"4f",x"26"),
   174 => (x"49",x"c0",x"ff",x"86"),
   175 => (x"c0",x"c4",x"48",x"69"),
   176 => (x"58",x"a6",x"c4",x"98"),
   177 => (x"87",x"f4",x"02",x"6e"),
   178 => (x"48",x"79",x"66",x"c8"),
   179 => (x"4f",x"26",x"8e",x"fc"),
   180 => (x"74",x"1e",x"73",x"1e"),
   181 => (x"4b",x"66",x"cc",x"1e"),
   182 => (x"4a",x"13",x"4c",x"c0"),
   183 => (x"d2",x"02",x"9a",x"72"),
   184 => (x"71",x"49",x"72",x"87"),
   185 => (x"87",x"ce",x"ff",x"1e"),
   186 => (x"84",x"c1",x"86",x"c4"),
   187 => (x"9a",x"72",x"4a",x"13"),
   188 => (x"74",x"87",x"ee",x"05"),
   189 => (x"26",x"4c",x"26",x"48"),
   190 => (x"1e",x"4f",x"26",x"4b"),
   191 => (x"9a",x"72",x"1e",x"73"),
   192 => (x"87",x"e7",x"c0",x"02"),
   193 => (x"4b",x"c1",x"48",x"c0"),
   194 => (x"d1",x"06",x"a9",x"72"),
   195 => (x"06",x"82",x"72",x"87"),
   196 => (x"83",x"73",x"87",x"c9"),
   197 => (x"f4",x"01",x"a9",x"72"),
   198 => (x"c1",x"87",x"c3",x"87"),
   199 => (x"a9",x"72",x"3a",x"b2"),
   200 => (x"80",x"73",x"89",x"03"),
   201 => (x"2b",x"2a",x"c1",x"07"),
   202 => (x"26",x"87",x"f3",x"05"),
   203 => (x"1e",x"4f",x"26",x"4b"),
   204 => (x"4d",x"c4",x"1e",x"75"),
   205 => (x"04",x"a1",x"b7",x"71"),
   206 => (x"81",x"c1",x"b9",x"ff"),
   207 => (x"72",x"07",x"bd",x"c3"),
   208 => (x"ff",x"04",x"a2",x"b7"),
   209 => (x"c1",x"82",x"c1",x"ba"),
   210 => (x"ee",x"fe",x"07",x"bd"),
   211 => (x"04",x"2d",x"c1",x"87"),
   212 => (x"80",x"c1",x"b8",x"ff"),
   213 => (x"ff",x"04",x"2d",x"07"),
   214 => (x"07",x"81",x"c1",x"b9"),
   215 => (x"4f",x"26",x"4d",x"26"),
   216 => (x"d0",x"1e",x"73",x"1e"),
   217 => (x"c0",x"c0",x"c0",x"c0"),
   218 => (x"fe",x"0f",x"73",x"4b"),
   219 => (x"26",x"87",x"c4",x"87"),
   220 => (x"26",x"4c",x"26",x"4d"),
   221 => (x"1e",x"4f",x"26",x"4b"),
   222 => (x"c3",x"49",x"66",x"c8"),
   223 => (x"f7",x"c0",x"99",x"df"),
   224 => (x"a9",x"b7",x"c0",x"89"),
   225 => (x"c0",x"87",x"c3",x"03"),
   226 => (x"66",x"c4",x"81",x"e7"),
   227 => (x"c8",x"30",x"c4",x"48"),
   228 => (x"66",x"c4",x"58",x"a6"),
   229 => (x"c8",x"b0",x"71",x"48"),
   230 => (x"66",x"c4",x"58",x"a6"),
   231 => (x"87",x"d5",x"ff",x"48"),
   232 => (x"74",x"1e",x"73",x"1e"),
   233 => (x"c0",x"c0",x"d0",x"1e"),
   234 => (x"c1",x"4c",x"c0",x"c0"),
   235 => (x"48",x"bf",x"c8",x"d4"),
   236 => (x"d4",x"c1",x"80",x"c1"),
   237 => (x"cc",x"97",x"58",x"cc"),
   238 => (x"c0",x"fe",x"49",x"66"),
   239 => (x"d3",x"c1",x"b9",x"81"),
   240 => (x"87",x"db",x"05",x"a9"),
   241 => (x"48",x"c8",x"d4",x"c1"),
   242 => (x"d4",x"c1",x"78",x"c0"),
   243 => (x"78",x"c0",x"48",x"cc"),
   244 => (x"48",x"d4",x"d4",x"c1"),
   245 => (x"d4",x"c1",x"78",x"c0"),
   246 => (x"78",x"c0",x"48",x"d8"),
   247 => (x"c1",x"87",x"f4",x"c6"),
   248 => (x"48",x"bf",x"c8",x"d4"),
   249 => (x"c0",x"05",x"a8",x"c1"),
   250 => (x"cc",x"97",x"87",x"f8"),
   251 => (x"c0",x"fe",x"49",x"66"),
   252 => (x"1e",x"71",x"b9",x"81"),
   253 => (x"bf",x"d8",x"d4",x"c1"),
   254 => (x"87",x"fb",x"fd",x"1e"),
   255 => (x"d4",x"c1",x"86",x"c8"),
   256 => (x"d4",x"c1",x"58",x"dc"),
   257 => (x"c3",x"4a",x"bf",x"d8"),
   258 => (x"c6",x"06",x"aa",x"b7"),
   259 => (x"72",x"48",x"ca",x"87"),
   260 => (x"72",x"4a",x"70",x"88"),
   261 => (x"71",x"81",x"c1",x"49"),
   262 => (x"c1",x"30",x"c1",x"48"),
   263 => (x"c5",x"58",x"d4",x"d4"),
   264 => (x"d4",x"c1",x"87",x"f1"),
   265 => (x"c9",x"48",x"bf",x"d8"),
   266 => (x"c5",x"01",x"a8",x"b7"),
   267 => (x"d4",x"c1",x"87",x"e5"),
   268 => (x"c0",x"48",x"bf",x"d8"),
   269 => (x"c5",x"06",x"a8",x"b7"),
   270 => (x"d4",x"c1",x"87",x"d9"),
   271 => (x"c3",x"48",x"bf",x"c8"),
   272 => (x"db",x"01",x"a8",x"b7"),
   273 => (x"66",x"cc",x"97",x"87"),
   274 => (x"81",x"c0",x"fe",x"49"),
   275 => (x"c1",x"1e",x"71",x"b9"),
   276 => (x"1e",x"bf",x"d4",x"d4"),
   277 => (x"c8",x"87",x"e0",x"fc"),
   278 => (x"d8",x"d4",x"c1",x"86"),
   279 => (x"87",x"f3",x"c4",x"58"),
   280 => (x"bf",x"d0",x"d4",x"c1"),
   281 => (x"c1",x"81",x"c3",x"49"),
   282 => (x"b7",x"bf",x"c8",x"d4"),
   283 => (x"e1",x"c0",x"04",x"a9"),
   284 => (x"66",x"cc",x"97",x"87"),
   285 => (x"81",x"c0",x"fe",x"49"),
   286 => (x"c1",x"1e",x"71",x"b9"),
   287 => (x"1e",x"bf",x"cc",x"d4"),
   288 => (x"c8",x"87",x"f4",x"fb"),
   289 => (x"d0",x"d4",x"c1",x"86"),
   290 => (x"dc",x"d4",x"c1",x"58"),
   291 => (x"c4",x"78",x"c1",x"48"),
   292 => (x"d4",x"c1",x"87",x"c1"),
   293 => (x"c0",x"48",x"bf",x"d8"),
   294 => (x"c2",x"06",x"a8",x"b7"),
   295 => (x"d4",x"c1",x"87",x"d8"),
   296 => (x"c3",x"48",x"bf",x"d8"),
   297 => (x"c2",x"01",x"a8",x"b7"),
   298 => (x"d4",x"c1",x"87",x"cc"),
   299 => (x"c1",x"49",x"bf",x"d4"),
   300 => (x"d4",x"c1",x"81",x"31"),
   301 => (x"a9",x"b7",x"bf",x"c8"),
   302 => (x"87",x"dc",x"c1",x"04"),
   303 => (x"49",x"66",x"cc",x"97"),
   304 => (x"b9",x"81",x"c0",x"fe"),
   305 => (x"d4",x"c1",x"1e",x"71"),
   306 => (x"fa",x"1e",x"bf",x"e0"),
   307 => (x"86",x"c8",x"87",x"e9"),
   308 => (x"58",x"e4",x"d4",x"c1"),
   309 => (x"bf",x"dc",x"d4",x"c1"),
   310 => (x"c1",x"89",x"c1",x"49"),
   311 => (x"c0",x"59",x"e0",x"d4"),
   312 => (x"c2",x"03",x"a9",x"b7"),
   313 => (x"d4",x"c1",x"87",x"ed"),
   314 => (x"c1",x"49",x"bf",x"cc"),
   315 => (x"bf",x"97",x"e0",x"d4"),
   316 => (x"cc",x"d4",x"c1",x"51"),
   317 => (x"81",x"c1",x"49",x"bf"),
   318 => (x"59",x"d0",x"d4",x"c1"),
   319 => (x"bf",x"e4",x"d4",x"c1"),
   320 => (x"c0",x"06",x"a9",x"b7"),
   321 => (x"d4",x"c1",x"87",x"c9"),
   322 => (x"d4",x"c1",x"48",x"e4"),
   323 => (x"c1",x"78",x"bf",x"cc"),
   324 => (x"c1",x"48",x"dc",x"d4"),
   325 => (x"87",x"fb",x"c1",x"78"),
   326 => (x"bf",x"dc",x"d4",x"c1"),
   327 => (x"87",x"f3",x"c1",x"05"),
   328 => (x"bf",x"e0",x"d4",x"c1"),
   329 => (x"c1",x"31",x"c4",x"49"),
   330 => (x"c1",x"59",x"e4",x"d4"),
   331 => (x"09",x"bf",x"cc",x"d4"),
   332 => (x"c1",x"09",x"79",x"97"),
   333 => (x"d4",x"c1",x"87",x"dd"),
   334 => (x"c7",x"48",x"bf",x"d8"),
   335 => (x"c1",x"04",x"a8",x"b7"),
   336 => (x"4b",x"c0",x"87",x"d1"),
   337 => (x"c1",x"48",x"f4",x"fe"),
   338 => (x"e4",x"d4",x"c1",x"78"),
   339 => (x"1e",x"74",x"1e",x"bf"),
   340 => (x"f5",x"1e",x"d6",x"d6"),
   341 => (x"86",x"cc",x"87",x"cd"),
   342 => (x"5c",x"d0",x"d4",x"c1"),
   343 => (x"bf",x"cc",x"d4",x"c1"),
   344 => (x"e4",x"d4",x"c1",x"48"),
   345 => (x"03",x"a8",x"b7",x"bf"),
   346 => (x"c1",x"87",x"db",x"c0"),
   347 => (x"bf",x"bf",x"cc",x"d4"),
   348 => (x"cc",x"d4",x"c1",x"83"),
   349 => (x"81",x"c4",x"49",x"bf"),
   350 => (x"59",x"d0",x"d4",x"c1"),
   351 => (x"bf",x"e4",x"d4",x"c1"),
   352 => (x"ff",x"04",x"a9",x"b7"),
   353 => (x"1e",x"73",x"87",x"e5"),
   354 => (x"f4",x"1e",x"f5",x"d6"),
   355 => (x"86",x"c8",x"87",x"d5"),
   356 => (x"f7",x"87",x"cd",x"f7"),
   357 => (x"68",x"43",x"87",x"db"),
   358 => (x"73",x"6b",x"63",x"65"),
   359 => (x"69",x"6d",x"6d",x"75"),
   360 => (x"66",x"20",x"67",x"6e"),
   361 => (x"20",x"6d",x"6f",x"72"),
   362 => (x"74",x"20",x"64",x"25"),
   363 => (x"64",x"25",x"20",x"6f"),
   364 => (x"20",x"2e",x"2e",x"2e"),
   365 => (x"0a",x"64",x"25",x"00"),
   366 => (x"6f",x"6f",x"42",x"00"),
   367 => (x"67",x"6e",x"69",x"74"),
   368 => (x"0a",x"2e",x"2e",x"2e"),
   369 => (x"4f",x"4f",x"42",x"00"),
   370 => (x"32",x"33",x"38",x"54"),
   371 => (x"4e",x"49",x"42",x"20"),
   372 => (x"20",x"44",x"53",x"00"),
   373 => (x"74",x"6f",x"6f",x"62"),
   374 => (x"69",x"61",x"66",x"20"),
   375 => (x"0a",x"64",x"65",x"6c"),
   376 => (x"69",x"6e",x"49",x"00"),
   377 => (x"6c",x"61",x"69",x"74"),
   378 => (x"6e",x"69",x"7a",x"69"),
   379 => (x"44",x"53",x"20",x"67"),
   380 => (x"72",x"61",x"63",x"20"),
   381 => (x"52",x"00",x"0a",x"64"),
   382 => (x"32",x"33",x"32",x"53"),
   383 => (x"6f",x"6f",x"62",x"20"),
   384 => (x"20",x"2d",x"20",x"74"),
   385 => (x"73",x"65",x"72",x"70"),
   386 => (x"53",x"45",x"20",x"73"),
   387 => (x"6f",x"74",x"20",x"43"),
   388 => (x"6f",x"6f",x"62",x"20"),
   389 => (x"72",x"66",x"20",x"74"),
   390 => (x"53",x"20",x"6d",x"6f"),
   391 => (x"1e",x"00",x"2e",x"44"),
   392 => (x"1e",x"74",x"1e",x"73"),
   393 => (x"e1",x"d7",x"1e",x"75"),
   394 => (x"87",x"e4",x"f2",x"1e"),
   395 => (x"ee",x"c0",x"86",x"c4"),
   396 => (x"98",x"70",x"87",x"c6"),
   397 => (x"c3",x"87",x"cc",x"02"),
   398 => (x"98",x"70",x"87",x"db"),
   399 => (x"c1",x"87",x"c4",x"02"),
   400 => (x"c0",x"87",x"c2",x"49"),
   401 => (x"d7",x"4d",x"71",x"49"),
   402 => (x"c3",x"f2",x"1e",x"f7"),
   403 => (x"c1",x"86",x"c4",x"87"),
   404 => (x"c0",x"48",x"e4",x"d4"),
   405 => (x"1e",x"ee",x"c0",x"78"),
   406 => (x"c4",x"87",x"db",x"f1"),
   407 => (x"c8",x"f4",x"c3",x"86"),
   408 => (x"c0",x"ff",x"4a",x"ff"),
   409 => (x"49",x"74",x"4c",x"bf"),
   410 => (x"02",x"99",x"c0",x"c8"),
   411 => (x"74",x"87",x"c5",x"c1"),
   412 => (x"9b",x"ff",x"c3",x"4b"),
   413 => (x"c0",x"05",x"ab",x"db"),
   414 => (x"9d",x"75",x"87",x"ee"),
   415 => (x"87",x"e0",x"c0",x"02"),
   416 => (x"c0",x"c0",x"c0",x"d0"),
   417 => (x"c5",x"d7",x"1e",x"c0"),
   418 => (x"87",x"d7",x"dc",x"1e"),
   419 => (x"98",x"70",x"86",x"c8"),
   420 => (x"d6",x"87",x"cd",x"02"),
   421 => (x"f7",x"f0",x"1e",x"f9"),
   422 => (x"f3",x"86",x"c4",x"87"),
   423 => (x"87",x"c8",x"87",x"c2"),
   424 => (x"f0",x"1e",x"d1",x"d7"),
   425 => (x"86",x"c4",x"87",x"ea"),
   426 => (x"f3",x"f3",x"1e",x"73"),
   427 => (x"c3",x"86",x"c4",x"87"),
   428 => (x"4a",x"c0",x"c9",x"f4"),
   429 => (x"8a",x"c1",x"49",x"72"),
   430 => (x"fe",x"05",x"99",x"71"),
   431 => (x"d4",x"fe",x"87",x"e4"),
   432 => (x"87",x"eb",x"f2",x"87"),
   433 => (x"c0",x"1e",x"73",x"1e"),
   434 => (x"48",x"66",x"d0",x"4b"),
   435 => (x"06",x"a8",x"b7",x"c0"),
   436 => (x"c8",x"87",x"f6",x"c0"),
   437 => (x"4a",x"bf",x"97",x"66"),
   438 => (x"ba",x"82",x"c0",x"fe"),
   439 => (x"c1",x"48",x"66",x"c8"),
   440 => (x"58",x"a6",x"cc",x"80"),
   441 => (x"bf",x"97",x"66",x"cc"),
   442 => (x"81",x"c0",x"fe",x"49"),
   443 => (x"48",x"66",x"cc",x"b9"),
   444 => (x"a6",x"d0",x"80",x"c1"),
   445 => (x"aa",x"b7",x"71",x"58"),
   446 => (x"c1",x"87",x"c4",x"02"),
   447 => (x"c1",x"87",x"cc",x"48"),
   448 => (x"b7",x"66",x"d0",x"83"),
   449 => (x"ca",x"ff",x"04",x"ab"),
   450 => (x"c4",x"48",x"c0",x"87"),
   451 => (x"26",x"4d",x"26",x"87"),
   452 => (x"26",x"4b",x"26",x"4c"),
   453 => (x"1e",x"73",x"1e",x"4f"),
   454 => (x"1e",x"75",x"1e",x"74"),
   455 => (x"48",x"f0",x"dc",x"c1"),
   456 => (x"eb",x"c0",x"78",x"c0"),
   457 => (x"e7",x"ee",x"1e",x"f2"),
   458 => (x"c1",x"86",x"c4",x"87"),
   459 => (x"c0",x"1e",x"e8",x"d4"),
   460 => (x"ec",x"ef",x"c0",x"1e"),
   461 => (x"70",x"86",x"c8",x"87"),
   462 => (x"87",x"ce",x"05",x"98"),
   463 => (x"1e",x"de",x"e8",x"c0"),
   464 => (x"c4",x"87",x"cd",x"ee"),
   465 => (x"cb",x"48",x"c0",x"86"),
   466 => (x"eb",x"c0",x"87",x"d1"),
   467 => (x"ff",x"ed",x"1e",x"ff"),
   468 => (x"c0",x"86",x"c4",x"87"),
   469 => (x"dc",x"dd",x"c1",x"4b"),
   470 => (x"c8",x"78",x"c1",x"48"),
   471 => (x"d6",x"ec",x"c0",x"1e"),
   472 => (x"de",x"d5",x"c1",x"1e"),
   473 => (x"87",x"dc",x"fd",x"1e"),
   474 => (x"98",x"70",x"86",x"cc"),
   475 => (x"c1",x"87",x"c6",x"05"),
   476 => (x"c0",x"48",x"dc",x"dd"),
   477 => (x"c0",x"1e",x"c8",x"78"),
   478 => (x"c1",x"1e",x"df",x"ec"),
   479 => (x"fd",x"1e",x"fa",x"d5"),
   480 => (x"86",x"cc",x"87",x"c2"),
   481 => (x"c6",x"05",x"98",x"70"),
   482 => (x"dc",x"dd",x"c1",x"87"),
   483 => (x"c1",x"78",x"c0",x"48"),
   484 => (x"1e",x"bf",x"dc",x"dd"),
   485 => (x"1e",x"e8",x"ec",x"c0"),
   486 => (x"c8",x"87",x"c8",x"ec"),
   487 => (x"dc",x"dd",x"c1",x"86"),
   488 => (x"d3",x"c2",x"02",x"bf"),
   489 => (x"e8",x"d4",x"c1",x"87"),
   490 => (x"e6",x"db",x"c1",x"4d"),
   491 => (x"e6",x"dc",x"c1",x"4c"),
   492 => (x"71",x"49",x"bf",x"9f"),
   493 => (x"e6",x"dc",x"c1",x"1e"),
   494 => (x"e8",x"d4",x"c1",x"49"),
   495 => (x"d0",x"1e",x"71",x"89"),
   496 => (x"1e",x"c0",x"c8",x"1e"),
   497 => (x"1e",x"d0",x"e9",x"c0"),
   498 => (x"d4",x"87",x"d8",x"eb"),
   499 => (x"49",x"a4",x"c8",x"86"),
   500 => (x"dc",x"c1",x"4b",x"69"),
   501 => (x"49",x"bf",x"9f",x"e6"),
   502 => (x"a9",x"ea",x"d6",x"c5"),
   503 => (x"87",x"d0",x"c0",x"05"),
   504 => (x"69",x"49",x"a4",x"c8"),
   505 => (x"dd",x"f3",x"c0",x"1e"),
   506 => (x"70",x"86",x"c4",x"87"),
   507 => (x"87",x"dd",x"c0",x"4b"),
   508 => (x"49",x"a5",x"fe",x"c7"),
   509 => (x"ca",x"49",x"69",x"9f"),
   510 => (x"02",x"a9",x"d5",x"e9"),
   511 => (x"c0",x"87",x"ce",x"c0"),
   512 => (x"eb",x"1e",x"f2",x"e8"),
   513 => (x"86",x"c4",x"87",x"ca"),
   514 => (x"ce",x"c8",x"48",x"c0"),
   515 => (x"c0",x"1e",x"73",x"87"),
   516 => (x"ea",x"1e",x"cd",x"ea"),
   517 => (x"86",x"c8",x"87",x"cd"),
   518 => (x"1e",x"e8",x"d4",x"c1"),
   519 => (x"eb",x"c0",x"1e",x"73"),
   520 => (x"86",x"c8",x"87",x"ff"),
   521 => (x"c0",x"05",x"98",x"70"),
   522 => (x"48",x"c0",x"87",x"c5"),
   523 => (x"c0",x"87",x"ec",x"c7"),
   524 => (x"ea",x"1e",x"e5",x"ea"),
   525 => (x"86",x"c4",x"87",x"da"),
   526 => (x"1e",x"fb",x"ec",x"c0"),
   527 => (x"c4",x"87",x"e4",x"e9"),
   528 => (x"c0",x"1e",x"c8",x"86"),
   529 => (x"c1",x"1e",x"d3",x"ed"),
   530 => (x"f9",x"1e",x"fa",x"d5"),
   531 => (x"86",x"cc",x"87",x"f6"),
   532 => (x"c0",x"05",x"98",x"70"),
   533 => (x"dc",x"c1",x"87",x"c9"),
   534 => (x"78",x"c1",x"48",x"f0"),
   535 => (x"c8",x"87",x"e3",x"c0"),
   536 => (x"dc",x"ed",x"c0",x"1e"),
   537 => (x"de",x"d5",x"c1",x"1e"),
   538 => (x"87",x"d8",x"f9",x"1e"),
   539 => (x"98",x"70",x"86",x"cc"),
   540 => (x"87",x"ce",x"c0",x"02"),
   541 => (x"1e",x"cc",x"eb",x"c0"),
   542 => (x"c4",x"87",x"e8",x"e8"),
   543 => (x"c6",x"48",x"c0",x"86"),
   544 => (x"dc",x"c1",x"87",x"d9"),
   545 => (x"49",x"bf",x"97",x"e6"),
   546 => (x"05",x"a9",x"d5",x"c1"),
   547 => (x"c1",x"87",x"cd",x"c0"),
   548 => (x"bf",x"97",x"e7",x"dc"),
   549 => (x"a9",x"ea",x"c2",x"49"),
   550 => (x"87",x"c5",x"c0",x"02"),
   551 => (x"fa",x"c5",x"48",x"c0"),
   552 => (x"e8",x"d4",x"c1",x"87"),
   553 => (x"c3",x"49",x"bf",x"97"),
   554 => (x"c0",x"02",x"a9",x"e9"),
   555 => (x"d4",x"c1",x"87",x"d2"),
   556 => (x"49",x"bf",x"97",x"e8"),
   557 => (x"02",x"a9",x"eb",x"c3"),
   558 => (x"c0",x"87",x"c5",x"c0"),
   559 => (x"87",x"db",x"c5",x"48"),
   560 => (x"97",x"f3",x"d4",x"c1"),
   561 => (x"99",x"71",x"49",x"bf"),
   562 => (x"87",x"cc",x"c0",x"05"),
   563 => (x"97",x"f4",x"d4",x"c1"),
   564 => (x"a9",x"c2",x"49",x"bf"),
   565 => (x"87",x"c5",x"c0",x"02"),
   566 => (x"fe",x"c4",x"48",x"c0"),
   567 => (x"f5",x"d4",x"c1",x"87"),
   568 => (x"c1",x"48",x"bf",x"97"),
   569 => (x"c1",x"58",x"ec",x"dc"),
   570 => (x"49",x"bf",x"e8",x"dc"),
   571 => (x"8a",x"c1",x"4a",x"71"),
   572 => (x"5a",x"f0",x"dc",x"c1"),
   573 => (x"1e",x"71",x"1e",x"72"),
   574 => (x"1e",x"e5",x"ed",x"c0"),
   575 => (x"cc",x"87",x"e4",x"e6"),
   576 => (x"f6",x"d4",x"c1",x"86"),
   577 => (x"73",x"49",x"bf",x"97"),
   578 => (x"f7",x"d4",x"c1",x"81"),
   579 => (x"c8",x"4a",x"bf",x"97"),
   580 => (x"fc",x"dc",x"c1",x"32"),
   581 => (x"78",x"a1",x"72",x"48"),
   582 => (x"97",x"f8",x"d4",x"c1"),
   583 => (x"dd",x"c1",x"48",x"bf"),
   584 => (x"dc",x"c1",x"58",x"d4"),
   585 => (x"c2",x"02",x"bf",x"f0"),
   586 => (x"1e",x"c8",x"87",x"df"),
   587 => (x"1e",x"e9",x"eb",x"c0"),
   588 => (x"1e",x"fa",x"d5",x"c1"),
   589 => (x"cc",x"87",x"cd",x"f6"),
   590 => (x"02",x"98",x"70",x"86"),
   591 => (x"c0",x"87",x"c5",x"c0"),
   592 => (x"87",x"d7",x"c3",x"48"),
   593 => (x"bf",x"e8",x"dc",x"c1"),
   594 => (x"c4",x"48",x"72",x"4a"),
   595 => (x"d8",x"dd",x"c1",x"30"),
   596 => (x"d0",x"dd",x"c1",x"58"),
   597 => (x"cd",x"d5",x"c1",x"5a"),
   598 => (x"c8",x"49",x"bf",x"97"),
   599 => (x"cc",x"d5",x"c1",x"31"),
   600 => (x"73",x"4b",x"bf",x"97"),
   601 => (x"d5",x"c1",x"49",x"a1"),
   602 => (x"4b",x"bf",x"97",x"ce"),
   603 => (x"a1",x"73",x"33",x"d0"),
   604 => (x"cf",x"d5",x"c1",x"49"),
   605 => (x"d8",x"4b",x"bf",x"97"),
   606 => (x"49",x"a1",x"73",x"33"),
   607 => (x"59",x"dc",x"dd",x"c1"),
   608 => (x"bf",x"d0",x"dd",x"c1"),
   609 => (x"fc",x"dc",x"c1",x"91"),
   610 => (x"dd",x"c1",x"81",x"bf"),
   611 => (x"d5",x"c1",x"59",x"c4"),
   612 => (x"4b",x"bf",x"97",x"d5"),
   613 => (x"d5",x"c1",x"33",x"c8"),
   614 => (x"4c",x"bf",x"97",x"d4"),
   615 => (x"c1",x"4b",x"a3",x"74"),
   616 => (x"bf",x"97",x"d6",x"d5"),
   617 => (x"74",x"34",x"d0",x"4c"),
   618 => (x"d5",x"c1",x"4b",x"a3"),
   619 => (x"4c",x"bf",x"97",x"d7"),
   620 => (x"34",x"d8",x"9c",x"cf"),
   621 => (x"c1",x"4b",x"a3",x"74"),
   622 => (x"c2",x"5b",x"c8",x"dd"),
   623 => (x"c1",x"92",x"73",x"8b"),
   624 => (x"72",x"48",x"c8",x"dd"),
   625 => (x"d0",x"c1",x"78",x"a1"),
   626 => (x"fa",x"d4",x"c1",x"87"),
   627 => (x"c8",x"49",x"bf",x"97"),
   628 => (x"f9",x"d4",x"c1",x"31"),
   629 => (x"72",x"4a",x"bf",x"97"),
   630 => (x"dd",x"c1",x"49",x"a1"),
   631 => (x"31",x"c5",x"59",x"d8"),
   632 => (x"c9",x"81",x"ff",x"c7"),
   633 => (x"d0",x"dd",x"c1",x"29"),
   634 => (x"ff",x"d4",x"c1",x"59"),
   635 => (x"c8",x"4a",x"bf",x"97"),
   636 => (x"fe",x"d4",x"c1",x"32"),
   637 => (x"73",x"4b",x"bf",x"97"),
   638 => (x"dd",x"c1",x"4a",x"a2"),
   639 => (x"dd",x"c1",x"5a",x"dc"),
   640 => (x"c1",x"92",x"bf",x"d0"),
   641 => (x"82",x"bf",x"fc",x"dc"),
   642 => (x"5a",x"cc",x"dd",x"c1"),
   643 => (x"48",x"c4",x"dd",x"c1"),
   644 => (x"dd",x"c1",x"78",x"c0"),
   645 => (x"a1",x"72",x"48",x"c0"),
   646 => (x"f3",x"48",x"c1",x"78"),
   647 => (x"65",x"52",x"87",x"ef"),
   648 => (x"6f",x"20",x"64",x"61"),
   649 => (x"42",x"4d",x"20",x"66"),
   650 => (x"61",x"66",x"20",x"52"),
   651 => (x"64",x"65",x"6c",x"69"),
   652 => (x"6f",x"4e",x"00",x"0a"),
   653 => (x"72",x"61",x"70",x"20"),
   654 => (x"69",x"74",x"69",x"74"),
   655 => (x"73",x"20",x"6e",x"6f"),
   656 => (x"61",x"6e",x"67",x"69"),
   657 => (x"65",x"72",x"75",x"74"),
   658 => (x"75",x"6f",x"66",x"20"),
   659 => (x"00",x"0a",x"64",x"6e"),
   660 => (x"73",x"52",x"42",x"4d"),
   661 => (x"3a",x"65",x"7a",x"69"),
   662 => (x"2c",x"64",x"25",x"20"),
   663 => (x"72",x"61",x"70",x"20"),
   664 => (x"69",x"74",x"69",x"74"),
   665 => (x"69",x"73",x"6e",x"6f"),
   666 => (x"20",x"3a",x"65",x"7a"),
   667 => (x"20",x"2c",x"64",x"25"),
   668 => (x"73",x"66",x"66",x"6f"),
   669 => (x"6f",x"20",x"74",x"65"),
   670 => (x"69",x"73",x"20",x"66"),
   671 => (x"25",x"20",x"3a",x"67"),
   672 => (x"73",x"20",x"2c",x"64"),
   673 => (x"30",x"20",x"67",x"69"),
   674 => (x"0a",x"78",x"25",x"78"),
   675 => (x"61",x"65",x"52",x"00"),
   676 => (x"67",x"6e",x"69",x"64"),
   677 => (x"6f",x"6f",x"62",x"20"),
   678 => (x"65",x"73",x"20",x"74"),
   679 => (x"72",x"6f",x"74",x"63"),
   680 => (x"0a",x"64",x"25",x"20"),
   681 => (x"61",x"65",x"52",x"00"),
   682 => (x"6f",x"62",x"20",x"64"),
   683 => (x"73",x"20",x"74",x"6f"),
   684 => (x"6f",x"74",x"63",x"65"),
   685 => (x"72",x"66",x"20",x"72"),
   686 => (x"66",x"20",x"6d",x"6f"),
   687 => (x"74",x"73",x"72",x"69"),
   688 => (x"72",x"61",x"70",x"20"),
   689 => (x"69",x"74",x"69",x"74"),
   690 => (x"00",x"0a",x"6e",x"6f"),
   691 => (x"75",x"73",x"6e",x"55"),
   692 => (x"72",x"6f",x"70",x"70"),
   693 => (x"20",x"64",x"65",x"74"),
   694 => (x"74",x"72",x"61",x"70"),
   695 => (x"6f",x"69",x"74",x"69"),
   696 => (x"79",x"74",x"20",x"6e"),
   697 => (x"0d",x"21",x"65",x"70"),
   698 => (x"54",x"41",x"46",x"00"),
   699 => (x"20",x"20",x"32",x"33"),
   700 => (x"65",x"52",x"00",x"20"),
   701 => (x"6e",x"69",x"64",x"61"),
   702 => (x"42",x"4d",x"20",x"67"),
   703 => (x"4d",x"00",x"0a",x"52"),
   704 => (x"73",x"20",x"52",x"42"),
   705 => (x"65",x"63",x"63",x"75"),
   706 => (x"75",x"66",x"73",x"73"),
   707 => (x"20",x"79",x"6c",x"6c"),
   708 => (x"64",x"61",x"65",x"72"),
   709 => (x"41",x"46",x"00",x"0a"),
   710 => (x"20",x"36",x"31",x"54"),
   711 => (x"46",x"00",x"20",x"20"),
   712 => (x"32",x"33",x"54",x"41"),
   713 => (x"00",x"20",x"20",x"20"),
   714 => (x"74",x"72",x"61",x"50"),
   715 => (x"6f",x"69",x"74",x"69"),
   716 => (x"75",x"6f",x"63",x"6e"),
   717 => (x"25",x"20",x"74",x"6e"),
   718 => (x"48",x"00",x"0a",x"64"),
   719 => (x"69",x"74",x"6e",x"75"),
   720 => (x"66",x"20",x"67",x"6e"),
   721 => (x"66",x"20",x"72",x"6f"),
   722 => (x"73",x"65",x"6c",x"69"),
   723 => (x"65",x"74",x"73",x"79"),
   724 => (x"46",x"00",x"0a",x"6d"),
   725 => (x"32",x"33",x"54",x"41"),
   726 => (x"00",x"20",x"20",x"20"),
   727 => (x"31",x"54",x"41",x"46"),
   728 => (x"20",x"20",x"20",x"36"),
   729 => (x"75",x"6c",x"43",x"00"),
   730 => (x"72",x"65",x"74",x"73"),
   731 => (x"7a",x"69",x"73",x"20"),
   732 => (x"25",x"20",x"3a",x"65"),
   733 => (x"43",x"20",x"2c",x"64"),
   734 => (x"74",x"73",x"75",x"6c"),
   735 => (x"6d",x"20",x"72",x"65"),
   736 => (x"2c",x"6b",x"73",x"61"),
   737 => (x"0a",x"64",x"25",x"20"),
   738 => (x"65",x"70",x"4f",x"00"),
   739 => (x"20",x"64",x"65",x"6e"),
   740 => (x"65",x"6c",x"69",x"66"),
   741 => (x"6f",x"6c",x"20",x"2c"),
   742 => (x"6e",x"69",x"64",x"61"),
   743 => (x"2e",x"2e",x"2e",x"67"),
   744 => (x"61",x"43",x"00",x"0a"),
   745 => (x"20",x"74",x"27",x"6e"),
   746 => (x"6e",x"65",x"70",x"6f"),
   747 => (x"0a",x"73",x"25",x"20"),
   748 => (x"1e",x"73",x"1e",x"00"),
   749 => (x"dc",x"c1",x"1e",x"74"),
   750 => (x"ce",x"02",x"bf",x"f0"),
   751 => (x"4a",x"66",x"cc",x"87"),
   752 => (x"cc",x"2a",x"b7",x"c7"),
   753 => (x"ff",x"c1",x"4b",x"66"),
   754 => (x"cc",x"87",x"cc",x"9b"),
   755 => (x"b7",x"c8",x"4a",x"66"),
   756 => (x"4b",x"66",x"cc",x"2a"),
   757 => (x"c1",x"9b",x"ff",x"c3"),
   758 => (x"c1",x"1e",x"e8",x"d4"),
   759 => (x"49",x"bf",x"fc",x"dc"),
   760 => (x"1e",x"71",x"81",x"72"),
   761 => (x"c8",x"87",x"fa",x"dc"),
   762 => (x"05",x"98",x"70",x"86"),
   763 => (x"48",x"c0",x"87",x"c5"),
   764 => (x"c1",x"87",x"e6",x"c0"),
   765 => (x"02",x"bf",x"f0",x"dc"),
   766 => (x"49",x"73",x"87",x"d2"),
   767 => (x"d4",x"c1",x"91",x"c4"),
   768 => (x"4c",x"69",x"81",x"e8"),
   769 => (x"ff",x"ff",x"ff",x"cf"),
   770 => (x"87",x"cb",x"9c",x"ff"),
   771 => (x"91",x"c2",x"49",x"73"),
   772 => (x"81",x"e8",x"d4",x"c1"),
   773 => (x"74",x"4c",x"69",x"9f"),
   774 => (x"87",x"f3",x"eb",x"48"),
   775 => (x"74",x"1e",x"73",x"1e"),
   776 => (x"f4",x"1e",x"75",x"1e"),
   777 => (x"c1",x"4b",x"c0",x"86"),
   778 => (x"7e",x"bf",x"c4",x"dd"),
   779 => (x"c1",x"48",x"a6",x"c4"),
   780 => (x"78",x"bf",x"c8",x"dd"),
   781 => (x"bf",x"f0",x"dc",x"c1"),
   782 => (x"c1",x"87",x"c9",x"02"),
   783 => (x"49",x"bf",x"e8",x"dc"),
   784 => (x"87",x"c7",x"31",x"c4"),
   785 => (x"bf",x"cc",x"dd",x"c1"),
   786 => (x"cc",x"31",x"c4",x"49"),
   787 => (x"4d",x"c0",x"59",x"a6"),
   788 => (x"c0",x"48",x"66",x"c8"),
   789 => (x"e9",x"c2",x"06",x"a8"),
   790 => (x"cf",x"49",x"75",x"87"),
   791 => (x"87",x"da",x"05",x"99"),
   792 => (x"1e",x"e8",x"d4",x"c1"),
   793 => (x"48",x"49",x"66",x"c8"),
   794 => (x"a6",x"cc",x"80",x"c1"),
   795 => (x"da",x"1e",x"71",x"58"),
   796 => (x"86",x"c8",x"87",x"ef"),
   797 => (x"4b",x"e8",x"d4",x"c1"),
   798 => (x"e0",x"c0",x"87",x"c3"),
   799 => (x"49",x"6b",x"97",x"83"),
   800 => (x"c1",x"02",x"99",x"71"),
   801 => (x"6b",x"97",x"87",x"f3"),
   802 => (x"a9",x"e5",x"c3",x"49"),
   803 => (x"87",x"e9",x"c1",x"02"),
   804 => (x"97",x"49",x"a3",x"cb"),
   805 => (x"99",x"d8",x"49",x"69"),
   806 => (x"87",x"dd",x"c1",x"05"),
   807 => (x"d8",x"ff",x"1e",x"73"),
   808 => (x"86",x"c4",x"87",x"ee"),
   809 => (x"e4",x"c0",x"1e",x"cb"),
   810 => (x"1e",x"73",x"1e",x"66"),
   811 => (x"cc",x"87",x"d5",x"e8"),
   812 => (x"05",x"98",x"70",x"86"),
   813 => (x"dc",x"87",x"c2",x"c1"),
   814 => (x"66",x"dc",x"4a",x"a3"),
   815 => (x"6a",x"81",x"c4",x"49"),
   816 => (x"4a",x"a3",x"da",x"79"),
   817 => (x"c8",x"49",x"66",x"dc"),
   818 => (x"48",x"6a",x"9f",x"81"),
   819 => (x"4c",x"71",x"79",x"70"),
   820 => (x"bf",x"f0",x"dc",x"c1"),
   821 => (x"d4",x"87",x"d0",x"02"),
   822 => (x"69",x"9f",x"49",x"a3"),
   823 => (x"c0",x"4a",x"71",x"49"),
   824 => (x"d0",x"9a",x"ff",x"ff"),
   825 => (x"c0",x"87",x"c2",x"32"),
   826 => (x"6c",x"48",x"72",x"4a"),
   827 => (x"dc",x"7c",x"70",x"80"),
   828 => (x"78",x"c0",x"48",x"66"),
   829 => (x"ff",x"c0",x"48",x"c1"),
   830 => (x"c8",x"85",x"c1",x"87"),
   831 => (x"fd",x"04",x"ad",x"66"),
   832 => (x"dc",x"c1",x"87",x"d7"),
   833 => (x"c0",x"02",x"bf",x"f0"),
   834 => (x"1e",x"6e",x"87",x"ec"),
   835 => (x"c4",x"87",x"e2",x"fa"),
   836 => (x"58",x"a6",x"c4",x"86"),
   837 => (x"ff",x"cf",x"49",x"6e"),
   838 => (x"99",x"f8",x"ff",x"ff"),
   839 => (x"87",x"d6",x"02",x"a9"),
   840 => (x"89",x"c2",x"49",x"6e"),
   841 => (x"bf",x"e8",x"dc",x"c1"),
   842 => (x"c0",x"dd",x"c1",x"91"),
   843 => (x"80",x"71",x"48",x"bf"),
   844 => (x"fc",x"58",x"a6",x"c8"),
   845 => (x"48",x"c0",x"87",x"d8"),
   846 => (x"d0",x"e7",x"8e",x"f4"),
   847 => (x"1e",x"73",x"1e",x"87"),
   848 => (x"49",x"bf",x"66",x"c8"),
   849 => (x"66",x"c8",x"81",x"c1"),
   850 => (x"c1",x"09",x"79",x"09"),
   851 => (x"99",x"bf",x"ec",x"dc"),
   852 => (x"c8",x"87",x"d0",x"05"),
   853 => (x"83",x"c8",x"4b",x"66"),
   854 => (x"d4",x"f9",x"1e",x"6b"),
   855 => (x"70",x"86",x"c4",x"87"),
   856 => (x"c1",x"7b",x"71",x"49"),
   857 => (x"87",x"e9",x"e6",x"48"),
   858 => (x"c0",x"dd",x"c1",x"1e"),
   859 => (x"66",x"c4",x"49",x"bf"),
   860 => (x"6a",x"82",x"c8",x"4a"),
   861 => (x"c1",x"8a",x"c2",x"4a"),
   862 => (x"92",x"bf",x"e8",x"dc"),
   863 => (x"c1",x"49",x"a1",x"72"),
   864 => (x"4a",x"bf",x"ec",x"dc"),
   865 => (x"9a",x"bf",x"66",x"c4"),
   866 => (x"c8",x"49",x"a1",x"72"),
   867 => (x"1e",x"71",x"1e",x"66"),
   868 => (x"c8",x"87",x"ce",x"d6"),
   869 => (x"05",x"98",x"70",x"86"),
   870 => (x"48",x"c0",x"87",x"c4"),
   871 => (x"48",x"c1",x"87",x"c2"),
   872 => (x"1e",x"87",x"f0",x"e5"),
   873 => (x"1e",x"74",x"1e",x"73"),
   874 => (x"c1",x"1e",x"66",x"cc"),
   875 => (x"f9",x"1e",x"e0",x"dd"),
   876 => (x"86",x"c8",x"87",x"ea"),
   877 => (x"c1",x"02",x"98",x"70"),
   878 => (x"dd",x"c1",x"87",x"d2"),
   879 => (x"c7",x"49",x"bf",x"e4"),
   880 => (x"29",x"c9",x"81",x"ff"),
   881 => (x"4b",x"c0",x"4c",x"71"),
   882 => (x"1e",x"c9",x"ee",x"c0"),
   883 => (x"87",x"c0",x"d4",x"ff"),
   884 => (x"b7",x"c0",x"86",x"c4"),
   885 => (x"c4",x"c1",x"06",x"ac"),
   886 => (x"1e",x"66",x"d0",x"87"),
   887 => (x"1e",x"e0",x"dd",x"c1"),
   888 => (x"c8",x"87",x"c5",x"fe"),
   889 => (x"05",x"98",x"70",x"86"),
   890 => (x"48",x"c0",x"87",x"c5"),
   891 => (x"c1",x"87",x"f0",x"c0"),
   892 => (x"fd",x"1e",x"e0",x"dd"),
   893 => (x"86",x"c4",x"87",x"c7"),
   894 => (x"c8",x"48",x"66",x"d0"),
   895 => (x"a6",x"d4",x"80",x"c0"),
   896 => (x"74",x"83",x"c1",x"58"),
   897 => (x"ff",x"04",x"ab",x"b7"),
   898 => (x"87",x"d1",x"87",x"cf"),
   899 => (x"c0",x"1e",x"66",x"cc"),
   900 => (x"ff",x"1e",x"e2",x"ee"),
   901 => (x"c8",x"87",x"cc",x"d2"),
   902 => (x"c2",x"48",x"c0",x"86"),
   903 => (x"e3",x"48",x"c1",x"87"),
   904 => (x"e8",x"1e",x"87",x"ed"),
   905 => (x"4a",x"d4",x"ff",x"86"),
   906 => (x"6a",x"7a",x"ff",x"c3"),
   907 => (x"7a",x"ff",x"c3",x"49"),
   908 => (x"30",x"c8",x"48",x"6a"),
   909 => (x"c8",x"58",x"a6",x"c4"),
   910 => (x"b1",x"6e",x"59",x"a6"),
   911 => (x"6a",x"7a",x"ff",x"c3"),
   912 => (x"cc",x"30",x"d0",x"48"),
   913 => (x"a6",x"d0",x"58",x"a6"),
   914 => (x"b1",x"66",x"c8",x"59"),
   915 => (x"6a",x"7a",x"ff",x"c3"),
   916 => (x"d4",x"30",x"d8",x"48"),
   917 => (x"a6",x"d8",x"58",x"a6"),
   918 => (x"b1",x"66",x"d0",x"59"),
   919 => (x"8e",x"e8",x"48",x"71"),
   920 => (x"f4",x"1e",x"4f",x"26"),
   921 => (x"4a",x"d4",x"ff",x"86"),
   922 => (x"6a",x"7a",x"ff",x"c3"),
   923 => (x"7a",x"ff",x"c3",x"49"),
   924 => (x"30",x"c8",x"48",x"71"),
   925 => (x"6a",x"58",x"a6",x"c4"),
   926 => (x"c3",x"b1",x"6e",x"49"),
   927 => (x"48",x"71",x"7a",x"ff"),
   928 => (x"a6",x"c8",x"30",x"c8"),
   929 => (x"c4",x"49",x"6a",x"58"),
   930 => (x"ff",x"c3",x"b1",x"66"),
   931 => (x"c8",x"48",x"71",x"7a"),
   932 => (x"58",x"a6",x"cc",x"30"),
   933 => (x"66",x"c8",x"49",x"6a"),
   934 => (x"f4",x"48",x"71",x"b1"),
   935 => (x"1e",x"4f",x"26",x"8e"),
   936 => (x"1e",x"74",x"1e",x"73"),
   937 => (x"ff",x"c3",x"1e",x"75"),
   938 => (x"4c",x"d4",x"ff",x"4d"),
   939 => (x"c3",x"48",x"66",x"d0"),
   940 => (x"7c",x"70",x"98",x"ff"),
   941 => (x"bf",x"f0",x"dd",x"c1"),
   942 => (x"d4",x"87",x"c8",x"05"),
   943 => (x"30",x"c9",x"48",x"66"),
   944 => (x"d4",x"58",x"a6",x"d8"),
   945 => (x"29",x"d8",x"49",x"66"),
   946 => (x"ff",x"c3",x"48",x"71"),
   947 => (x"d4",x"7c",x"70",x"98"),
   948 => (x"29",x"d0",x"49",x"66"),
   949 => (x"ff",x"c3",x"48",x"71"),
   950 => (x"d4",x"7c",x"70",x"98"),
   951 => (x"29",x"c8",x"49",x"66"),
   952 => (x"ff",x"c3",x"48",x"71"),
   953 => (x"d4",x"7c",x"70",x"98"),
   954 => (x"ff",x"c3",x"48",x"66"),
   955 => (x"d0",x"7c",x"70",x"98"),
   956 => (x"29",x"d0",x"49",x"66"),
   957 => (x"ff",x"c3",x"48",x"71"),
   958 => (x"6c",x"7c",x"70",x"98"),
   959 => (x"ff",x"f0",x"c9",x"4b"),
   960 => (x"05",x"ab",x"75",x"4a"),
   961 => (x"7c",x"75",x"87",x"ce"),
   962 => (x"8a",x"c1",x"4b",x"6c"),
   963 => (x"75",x"87",x"c5",x"02"),
   964 => (x"87",x"f2",x"02",x"ab"),
   965 => (x"4d",x"26",x"48",x"73"),
   966 => (x"4b",x"26",x"4c",x"26"),
   967 => (x"c0",x"1e",x"4f",x"26"),
   968 => (x"48",x"d4",x"ff",x"49"),
   969 => (x"c1",x"78",x"ff",x"c3"),
   970 => (x"b7",x"c8",x"c3",x"81"),
   971 => (x"87",x"f1",x"04",x"a9"),
   972 => (x"73",x"1e",x"4f",x"26"),
   973 => (x"75",x"1e",x"74",x"1e"),
   974 => (x"f0",x"ff",x"c0",x"1e"),
   975 => (x"c1",x"4d",x"f7",x"c1"),
   976 => (x"c0",x"c0",x"c0",x"c0"),
   977 => (x"d5",x"ff",x"4b",x"c0"),
   978 => (x"df",x"f8",x"c4",x"87"),
   979 => (x"75",x"1e",x"c0",x"4c"),
   980 => (x"87",x"cb",x"fd",x"1e"),
   981 => (x"a8",x"c1",x"86",x"c8"),
   982 => (x"87",x"e5",x"c0",x"05"),
   983 => (x"c3",x"48",x"d4",x"ff"),
   984 => (x"1e",x"73",x"78",x"ff"),
   985 => (x"c1",x"f0",x"e1",x"c0"),
   986 => (x"f2",x"fc",x"1e",x"e9"),
   987 => (x"70",x"86",x"c8",x"87"),
   988 => (x"87",x"ca",x"05",x"98"),
   989 => (x"c3",x"48",x"d4",x"ff"),
   990 => (x"48",x"c1",x"78",x"ff"),
   991 => (x"dd",x"fe",x"87",x"cb"),
   992 => (x"05",x"8c",x"c1",x"87"),
   993 => (x"c0",x"87",x"c6",x"ff"),
   994 => (x"26",x"4d",x"26",x"48"),
   995 => (x"26",x"4b",x"26",x"4c"),
   996 => (x"1e",x"73",x"1e",x"4f"),
   997 => (x"ff",x"c0",x"1e",x"74"),
   998 => (x"4c",x"c1",x"c1",x"f0"),
   999 => (x"c3",x"48",x"d4",x"ff"),
  1000 => (x"ff",x"c0",x"78",x"ff"),
  1001 => (x"cc",x"ff",x"1e",x"d7"),
  1002 => (x"86",x"c4",x"87",x"e6"),
  1003 => (x"1e",x"c0",x"4b",x"d3"),
  1004 => (x"ea",x"fb",x"1e",x"74"),
  1005 => (x"70",x"86",x"c8",x"87"),
  1006 => (x"87",x"ca",x"05",x"98"),
  1007 => (x"c3",x"48",x"d4",x"ff"),
  1008 => (x"48",x"c1",x"78",x"ff"),
  1009 => (x"d5",x"fd",x"87",x"cb"),
  1010 => (x"05",x"8b",x"c1",x"87"),
  1011 => (x"c0",x"87",x"df",x"ff"),
  1012 => (x"26",x"4c",x"26",x"48"),
  1013 => (x"43",x"4f",x"26",x"4b"),
  1014 => (x"43",x"00",x"44",x"4d"),
  1015 => (x"38",x"35",x"44",x"4d"),
  1016 => (x"0a",x"64",x"25",x"20"),
  1017 => (x"43",x"00",x"20",x"20"),
  1018 => (x"38",x"35",x"44",x"4d"),
  1019 => (x"25",x"20",x"32",x"5f"),
  1020 => (x"20",x"20",x"0a",x"64"),
  1021 => (x"44",x"4d",x"43",x"00"),
  1022 => (x"25",x"20",x"38",x"35"),
  1023 => (x"20",x"20",x"0a",x"64"),
  1024 => (x"48",x"44",x"53",x"00"),
  1025 => (x"6e",x"49",x"20",x"43"),
  1026 => (x"61",x"69",x"74",x"69"),
  1027 => (x"61",x"7a",x"69",x"6c"),
  1028 => (x"6e",x"6f",x"69",x"74"),
  1029 => (x"72",x"72",x"65",x"20"),
  1030 => (x"0a",x"21",x"72",x"6f"),
  1031 => (x"64",x"6d",x"63",x"00"),
  1032 => (x"44",x"4d",x"43",x"5f"),
  1033 => (x"65",x"72",x"20",x"38"),
  1034 => (x"6e",x"6f",x"70",x"73"),
  1035 => (x"20",x"3a",x"65",x"73"),
  1036 => (x"00",x"0a",x"64",x"25"),
  1037 => (x"52",x"52",x"45",x"49"),
  1038 => (x"49",x"50",x"53",x"00"),
  1039 => (x"20",x"44",x"53",x"00"),
  1040 => (x"64",x"72",x"61",x"63"),
  1041 => (x"7a",x"69",x"73",x"20"),
  1042 => (x"73",x"69",x"20",x"65"),
  1043 => (x"0a",x"64",x"25",x"20"),
  1044 => (x"69",x"72",x"57",x"00"),
  1045 => (x"66",x"20",x"65",x"74"),
  1046 => (x"65",x"6c",x"69",x"61"),
  1047 => (x"52",x"00",x"0a",x"64"),
  1048 => (x"20",x"64",x"61",x"65"),
  1049 => (x"6d",x"6d",x"6f",x"63"),
  1050 => (x"20",x"64",x"6e",x"61"),
  1051 => (x"6c",x"69",x"61",x"66"),
  1052 => (x"61",x"20",x"64",x"65"),
  1053 => (x"64",x"25",x"20",x"74"),
  1054 => (x"64",x"25",x"28",x"20"),
  1055 => (x"63",x"00",x"0a",x"29"),
  1056 => (x"7a",x"69",x"73",x"5f"),
  1057 => (x"75",x"6d",x"5f",x"65"),
  1058 => (x"20",x"3a",x"74",x"6c"),
  1059 => (x"20",x"2c",x"64",x"25"),
  1060 => (x"64",x"61",x"65",x"72"),
  1061 => (x"5f",x"6c",x"62",x"5f"),
  1062 => (x"3a",x"6e",x"65",x"6c"),
  1063 => (x"2c",x"64",x"25",x"20"),
  1064 => (x"69",x"73",x"63",x"20"),
  1065 => (x"20",x"3a",x"65",x"7a"),
  1066 => (x"00",x"0a",x"64",x"25"),
  1067 => (x"74",x"6c",x"75",x"4d"),
  1068 => (x"0a",x"64",x"25",x"20"),
  1069 => (x"20",x"64",x"25",x"00"),
  1070 => (x"63",x"6f",x"6c",x"62"),
  1071 => (x"6f",x"20",x"73",x"6b"),
  1072 => (x"69",x"73",x"20",x"66"),
  1073 => (x"25",x"20",x"65",x"7a"),
  1074 => (x"25",x"00",x"0a",x"64"),
  1075 => (x"6c",x"62",x"20",x"64"),
  1076 => (x"73",x"6b",x"63",x"6f"),
  1077 => (x"20",x"66",x"6f",x"20"),
  1078 => (x"20",x"32",x"31",x"35"),
  1079 => (x"65",x"74",x"79",x"62"),
  1080 => (x"1e",x"00",x"0a",x"73"),
  1081 => (x"1e",x"74",x"1e",x"73"),
  1082 => (x"d4",x"ff",x"1e",x"75"),
  1083 => (x"87",x"ee",x"f8",x"4c"),
  1084 => (x"c0",x"1e",x"ea",x"c6"),
  1085 => (x"c8",x"c1",x"f0",x"e1"),
  1086 => (x"87",x"e3",x"f6",x"1e"),
  1087 => (x"4b",x"70",x"86",x"c8"),
  1088 => (x"c0",x"c1",x"1e",x"73"),
  1089 => (x"c6",x"ff",x"1e",x"dd"),
  1090 => (x"86",x"c8",x"87",x"d9"),
  1091 => (x"c8",x"02",x"ab",x"c1"),
  1092 => (x"87",x"fd",x"f9",x"87"),
  1093 => (x"d7",x"c2",x"48",x"c0"),
  1094 => (x"87",x"c6",x"f5",x"87"),
  1095 => (x"ff",x"cf",x"49",x"70"),
  1096 => (x"ea",x"c6",x"99",x"ff"),
  1097 => (x"87",x"c8",x"02",x"a9"),
  1098 => (x"c0",x"87",x"e6",x"f9"),
  1099 => (x"87",x"c0",x"c2",x"48"),
  1100 => (x"c0",x"7c",x"ff",x"c3"),
  1101 => (x"f9",x"f7",x"4d",x"f1"),
  1102 => (x"02",x"98",x"70",x"87"),
  1103 => (x"c0",x"87",x"d6",x"c1"),
  1104 => (x"f0",x"ff",x"c0",x"1e"),
  1105 => (x"f5",x"1e",x"fa",x"c1"),
  1106 => (x"86",x"c8",x"87",x"d5"),
  1107 => (x"9b",x"73",x"4b",x"70"),
  1108 => (x"87",x"f5",x"c0",x"05"),
  1109 => (x"ff",x"c0",x"1e",x"73"),
  1110 => (x"c5",x"ff",x"1e",x"db"),
  1111 => (x"86",x"c8",x"87",x"c5"),
  1112 => (x"6c",x"7c",x"ff",x"c3"),
  1113 => (x"c0",x"1e",x"73",x"4b"),
  1114 => (x"ff",x"1e",x"e7",x"ff"),
  1115 => (x"c8",x"87",x"f4",x"c4"),
  1116 => (x"7c",x"ff",x"c3",x"86"),
  1117 => (x"73",x"7c",x"7c",x"7c"),
  1118 => (x"99",x"c0",x"c1",x"49"),
  1119 => (x"c1",x"87",x"c5",x"02"),
  1120 => (x"87",x"ec",x"c0",x"48"),
  1121 => (x"e7",x"c0",x"48",x"c0"),
  1122 => (x"c0",x"1e",x"73",x"87"),
  1123 => (x"ff",x"1e",x"f5",x"ff"),
  1124 => (x"c8",x"87",x"d0",x"c4"),
  1125 => (x"05",x"ad",x"c2",x"86"),
  1126 => (x"c0",x"c1",x"87",x"ce"),
  1127 => (x"c4",x"ff",x"1e",x"c1"),
  1128 => (x"86",x"c4",x"87",x"c1"),
  1129 => (x"87",x"c8",x"48",x"c0"),
  1130 => (x"fe",x"05",x"8d",x"c1"),
  1131 => (x"48",x"c0",x"87",x"c8"),
  1132 => (x"4c",x"26",x"4d",x"26"),
  1133 => (x"4f",x"26",x"4b",x"26"),
  1134 => (x"74",x"1e",x"73",x"1e"),
  1135 => (x"fc",x"1e",x"75",x"1e"),
  1136 => (x"4c",x"d0",x"ff",x"86"),
  1137 => (x"4b",x"c0",x"c0",x"c8"),
  1138 => (x"48",x"f0",x"dd",x"c1"),
  1139 => (x"c0",x"c1",x"78",x"c1"),
  1140 => (x"c3",x"ff",x"1e",x"f9"),
  1141 => (x"86",x"c4",x"87",x"fa"),
  1142 => (x"48",x"6c",x"4d",x"c7"),
  1143 => (x"a6",x"c4",x"98",x"73"),
  1144 => (x"cb",x"02",x"6e",x"58"),
  1145 => (x"73",x"48",x"6c",x"87"),
  1146 => (x"58",x"a6",x"c4",x"98"),
  1147 => (x"87",x"f5",x"05",x"6e"),
  1148 => (x"e9",x"f4",x"7c",x"c0"),
  1149 => (x"73",x"48",x"6c",x"87"),
  1150 => (x"58",x"a6",x"c4",x"98"),
  1151 => (x"87",x"cb",x"02",x"6e"),
  1152 => (x"98",x"73",x"48",x"6c"),
  1153 => (x"6e",x"58",x"a6",x"c4"),
  1154 => (x"c1",x"87",x"f5",x"05"),
  1155 => (x"c0",x"1e",x"c0",x"7c"),
  1156 => (x"c0",x"c1",x"d0",x"e5"),
  1157 => (x"87",x"c7",x"f2",x"1e"),
  1158 => (x"a8",x"c1",x"86",x"c8"),
  1159 => (x"c1",x"87",x"c2",x"05"),
  1160 => (x"05",x"ad",x"c2",x"4d"),
  1161 => (x"c0",x"c1",x"87",x"cf"),
  1162 => (x"c2",x"ff",x"1e",x"f4"),
  1163 => (x"86",x"c4",x"87",x"e2"),
  1164 => (x"de",x"c1",x"48",x"c0"),
  1165 => (x"05",x"8d",x"c1",x"87"),
  1166 => (x"fa",x"87",x"df",x"fe"),
  1167 => (x"dd",x"c1",x"87",x"e5"),
  1168 => (x"dd",x"c1",x"58",x"f4"),
  1169 => (x"cd",x"05",x"bf",x"f0"),
  1170 => (x"c0",x"1e",x"c1",x"87"),
  1171 => (x"d0",x"c1",x"f0",x"ff"),
  1172 => (x"87",x"cb",x"f1",x"1e"),
  1173 => (x"d4",x"ff",x"86",x"c8"),
  1174 => (x"78",x"ff",x"c3",x"48"),
  1175 => (x"c1",x"87",x"d1",x"c5"),
  1176 => (x"c1",x"58",x"f8",x"dd"),
  1177 => (x"1e",x"bf",x"f4",x"dd"),
  1178 => (x"1e",x"fd",x"c0",x"c1"),
  1179 => (x"87",x"f3",x"c0",x"ff"),
  1180 => (x"48",x"6c",x"86",x"c8"),
  1181 => (x"a6",x"c4",x"98",x"73"),
  1182 => (x"cc",x"02",x"6e",x"58"),
  1183 => (x"73",x"48",x"6c",x"87"),
  1184 => (x"58",x"a6",x"c4",x"98"),
  1185 => (x"f4",x"ff",x"05",x"6e"),
  1186 => (x"ff",x"7c",x"c0",x"87"),
  1187 => (x"ff",x"c3",x"48",x"d4"),
  1188 => (x"fc",x"48",x"c1",x"78"),
  1189 => (x"26",x"4d",x"26",x"8e"),
  1190 => (x"26",x"4b",x"26",x"4c"),
  1191 => (x"1e",x"73",x"1e",x"4f"),
  1192 => (x"1e",x"75",x"1e",x"74"),
  1193 => (x"d4",x"4d",x"d4",x"ff"),
  1194 => (x"66",x"d0",x"4c",x"66"),
  1195 => (x"c5",x"4a",x"c0",x"4b"),
  1196 => (x"49",x"df",x"cd",x"ee"),
  1197 => (x"6d",x"7d",x"ff",x"c3"),
  1198 => (x"a8",x"fe",x"c3",x"48"),
  1199 => (x"87",x"ce",x"c1",x"05"),
  1200 => (x"48",x"ec",x"dd",x"c1"),
  1201 => (x"b7",x"c4",x"78",x"c0"),
  1202 => (x"87",x"db",x"04",x"ac"),
  1203 => (x"70",x"87",x"d3",x"ed"),
  1204 => (x"c4",x"7b",x"71",x"49"),
  1205 => (x"ec",x"dd",x"c1",x"83"),
  1206 => (x"80",x"71",x"48",x"bf"),
  1207 => (x"58",x"f0",x"dd",x"c1"),
  1208 => (x"ac",x"b7",x"8c",x"c4"),
  1209 => (x"c0",x"87",x"e5",x"03"),
  1210 => (x"de",x"06",x"ac",x"b7"),
  1211 => (x"7d",x"ff",x"c3",x"87"),
  1212 => (x"97",x"71",x"49",x"6d"),
  1213 => (x"c1",x"83",x"c1",x"7b"),
  1214 => (x"48",x"bf",x"ec",x"dd"),
  1215 => (x"dd",x"c1",x"80",x"71"),
  1216 => (x"8c",x"c1",x"58",x"f0"),
  1217 => (x"01",x"ac",x"b7",x"c0"),
  1218 => (x"c1",x"87",x"e2",x"ff"),
  1219 => (x"89",x"c1",x"4a",x"49"),
  1220 => (x"87",x"e0",x"fe",x"05"),
  1221 => (x"72",x"7d",x"ff",x"c3"),
  1222 => (x"26",x"4d",x"26",x"48"),
  1223 => (x"26",x"4b",x"26",x"4c"),
  1224 => (x"1e",x"73",x"1e",x"4f"),
  1225 => (x"1e",x"75",x"1e",x"74"),
  1226 => (x"d0",x"ff",x"86",x"fc"),
  1227 => (x"c0",x"c0",x"c8",x"4c"),
  1228 => (x"ff",x"4d",x"c0",x"4b"),
  1229 => (x"ff",x"c3",x"48",x"d4"),
  1230 => (x"73",x"48",x"6c",x"78"),
  1231 => (x"58",x"a6",x"c4",x"98"),
  1232 => (x"87",x"cb",x"02",x"6e"),
  1233 => (x"98",x"73",x"48",x"6c"),
  1234 => (x"6e",x"58",x"a6",x"c4"),
  1235 => (x"c4",x"87",x"f5",x"05"),
  1236 => (x"d4",x"ff",x"7c",x"c1"),
  1237 => (x"78",x"ff",x"c3",x"48"),
  1238 => (x"c0",x"1e",x"66",x"d4"),
  1239 => (x"d1",x"c1",x"f0",x"ff"),
  1240 => (x"87",x"fb",x"ec",x"1e"),
  1241 => (x"49",x"70",x"86",x"c8"),
  1242 => (x"d2",x"02",x"99",x"71"),
  1243 => (x"d8",x"1e",x"71",x"87"),
  1244 => (x"c1",x"c1",x"1e",x"66"),
  1245 => (x"fc",x"fe",x"1e",x"df"),
  1246 => (x"86",x"cc",x"87",x"e9"),
  1247 => (x"c8",x"87",x"e5",x"c0"),
  1248 => (x"66",x"dc",x"1e",x"c0"),
  1249 => (x"87",x"d5",x"fc",x"1e"),
  1250 => (x"4d",x"70",x"86",x"c8"),
  1251 => (x"98",x"73",x"48",x"6c"),
  1252 => (x"6e",x"58",x"a6",x"c4"),
  1253 => (x"6c",x"87",x"cb",x"02"),
  1254 => (x"c4",x"98",x"73",x"48"),
  1255 => (x"05",x"6e",x"58",x"a6"),
  1256 => (x"7c",x"c0",x"87",x"f5"),
  1257 => (x"8e",x"fc",x"48",x"75"),
  1258 => (x"4c",x"26",x"4d",x"26"),
  1259 => (x"4f",x"26",x"4b",x"26"),
  1260 => (x"74",x"1e",x"73",x"1e"),
  1261 => (x"fc",x"1e",x"75",x"1e"),
  1262 => (x"c0",x"1e",x"c0",x"86"),
  1263 => (x"c9",x"c1",x"f0",x"ff"),
  1264 => (x"87",x"db",x"eb",x"1e"),
  1265 => (x"1e",x"d2",x"86",x"c8"),
  1266 => (x"1e",x"fe",x"dd",x"c1"),
  1267 => (x"c8",x"87",x"ce",x"fb"),
  1268 => (x"c1",x"4d",x"c0",x"86"),
  1269 => (x"ad",x"b7",x"d2",x"85"),
  1270 => (x"c1",x"87",x"f8",x"04"),
  1271 => (x"bf",x"97",x"fe",x"dd"),
  1272 => (x"99",x"c0",x"c3",x"49"),
  1273 => (x"05",x"a9",x"c0",x"c1"),
  1274 => (x"c1",x"87",x"e8",x"c0"),
  1275 => (x"bf",x"97",x"c5",x"de"),
  1276 => (x"c1",x"31",x"d0",x"49"),
  1277 => (x"bf",x"97",x"c6",x"de"),
  1278 => (x"72",x"32",x"c8",x"4a"),
  1279 => (x"c7",x"de",x"c1",x"b1"),
  1280 => (x"72",x"4a",x"bf",x"97"),
  1281 => (x"cf",x"4d",x"71",x"b1"),
  1282 => (x"9d",x"ff",x"ff",x"ff"),
  1283 => (x"35",x"ca",x"85",x"c1"),
  1284 => (x"c1",x"87",x"e7",x"c2"),
  1285 => (x"bf",x"97",x"c7",x"de"),
  1286 => (x"c6",x"33",x"c1",x"4b"),
  1287 => (x"c8",x"de",x"c1",x"9b"),
  1288 => (x"c7",x"49",x"bf",x"97"),
  1289 => (x"b3",x"71",x"29",x"b7"),
  1290 => (x"97",x"c3",x"de",x"c1"),
  1291 => (x"48",x"71",x"49",x"bf"),
  1292 => (x"a6",x"c4",x"98",x"cf"),
  1293 => (x"c4",x"de",x"c1",x"58"),
  1294 => (x"c3",x"4c",x"bf",x"97"),
  1295 => (x"c1",x"34",x"ca",x"9c"),
  1296 => (x"bf",x"97",x"c5",x"de"),
  1297 => (x"71",x"31",x"c2",x"49"),
  1298 => (x"c6",x"de",x"c1",x"b4"),
  1299 => (x"c3",x"49",x"bf",x"97"),
  1300 => (x"b7",x"c6",x"99",x"c0"),
  1301 => (x"74",x"b4",x"71",x"29"),
  1302 => (x"1e",x"66",x"c4",x"1e"),
  1303 => (x"c1",x"c1",x"1e",x"73"),
  1304 => (x"f8",x"fe",x"1e",x"ff"),
  1305 => (x"86",x"d0",x"87",x"fd"),
  1306 => (x"48",x"c1",x"83",x"c2"),
  1307 => (x"4b",x"70",x"30",x"73"),
  1308 => (x"c2",x"c1",x"1e",x"73"),
  1309 => (x"f8",x"fe",x"1e",x"ec"),
  1310 => (x"86",x"c8",x"87",x"e9"),
  1311 => (x"30",x"6e",x"48",x"c1"),
  1312 => (x"c1",x"58",x"a6",x"c4"),
  1313 => (x"73",x"4d",x"49",x"a4"),
  1314 => (x"75",x"1e",x"6e",x"95"),
  1315 => (x"f5",x"c2",x"c1",x"1e"),
  1316 => (x"ce",x"f8",x"fe",x"1e"),
  1317 => (x"6e",x"86",x"cc",x"87"),
  1318 => (x"b7",x"c0",x"c8",x"48"),
  1319 => (x"87",x"ce",x"06",x"a8"),
  1320 => (x"35",x"c1",x"4b",x"6e"),
  1321 => (x"c0",x"c8",x"2b",x"b7"),
  1322 => (x"ff",x"01",x"ab",x"b7"),
  1323 => (x"1e",x"75",x"87",x"f4"),
  1324 => (x"1e",x"cb",x"c3",x"c1"),
  1325 => (x"87",x"eb",x"f7",x"fe"),
  1326 => (x"48",x"75",x"86",x"c8"),
  1327 => (x"4d",x"26",x"8e",x"fc"),
  1328 => (x"4b",x"26",x"4c",x"26"),
  1329 => (x"c4",x"1e",x"4f",x"26"),
  1330 => (x"29",x"d8",x"49",x"66"),
  1331 => (x"c4",x"99",x"ff",x"c3"),
  1332 => (x"2a",x"c8",x"4a",x"66"),
  1333 => (x"9a",x"c0",x"fc",x"cf"),
  1334 => (x"66",x"c4",x"b1",x"72"),
  1335 => (x"c0",x"32",x"c8",x"4a"),
  1336 => (x"c0",x"c0",x"f0",x"ff"),
  1337 => (x"c4",x"b1",x"72",x"9a"),
  1338 => (x"32",x"d8",x"4a",x"66"),
  1339 => (x"c0",x"c0",x"c0",x"ff"),
  1340 => (x"b1",x"72",x"9a",x"c0"),
  1341 => (x"4f",x"26",x"48",x"71"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
