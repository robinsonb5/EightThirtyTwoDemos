library ieee;
use ieee.std_logic_1164.all;

package board_pkg is
	constant board_sdram_width : integer := 32;
	constant board_sdram_dqm : integer := 4;
end package;

