
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2a",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"82"),
    10 => (x"e0",x"c1",x"4f",x"4f"),
    11 => (x"c0",x"c1",x"4e",x"c4"),
    12 => (x"e0",x"c1",x"86",x"c0"),
    13 => (x"d5",x"c1",x"49",x"c4"),
    14 => (x"d0",x"89",x"48",x"ec"),
    15 => (x"40",x"c0",x"03",x"89"),
    16 => (x"f6",x"40",x"40",x"40"),
    17 => (x"05",x"81",x"d0",x"87"),
    18 => (x"89",x"c1",x"50",x"c0"),
    19 => (x"c1",x"87",x"f9",x"05"),
    20 => (x"c1",x"4c",x"eb",x"d5"),
    21 => (x"74",x"4d",x"eb",x"d5"),
    22 => (x"87",x"c6",x"02",x"ad"),
    23 => (x"0f",x"6c",x"8c",x"c4"),
    24 => (x"d9",x"af",x"87",x"f5"),
    25 => (x"6b",x"27",x"87",x"e3"),
    26 => (x"4c",x"00",x"00",x"15"),
    27 => (x"00",x"15",x"6b",x"27"),
    28 => (x"ad",x"74",x"4d",x"00"),
    29 => (x"24",x"87",x"c4",x"02"),
    30 => (x"00",x"87",x"f7",x"0f"),
    31 => (x"00",x"00",x"87",x"fd"),
    32 => (x"e0",x"c1",x"00",x"00"),
    33 => (x"c0",x"c1",x"4e",x"c4"),
    34 => (x"00",x"86",x"86",x"c0"),
    35 => (x"87",x"d1",x"db",x"98"),
    36 => (x"87",x"fc",x"98",x"00"),
    37 => (x"00",x"00",x"00",x"00"),
    38 => (x"bf",x"a7",x"f9",x"48"),
    39 => (x"c1",x"48",x"4f",x"08"),
    40 => (x"59",x"a7",x"f5",x"49"),
    41 => (x"70",x"70",x"00",x"af"),
    42 => (x"87",x"ec",x"1e",x"4f"),
    43 => (x"c0",x"05",x"98",x"48"),
    44 => (x"58",x"a7",x"e5",x"48"),
    45 => (x"4f",x"26",x"af",x"07"),
    46 => (x"5c",x"5b",x"5e",x"0e"),
    47 => (x"86",x"fc",x"0e",x"5d"),
    48 => (x"e0",x"c0",x"4a",x"71"),
    49 => (x"d5",x"c1",x"4c",x"66"),
    50 => (x"7e",x"c0",x"4b",x"ec"),
    51 => (x"ce",x"05",x"9a",x"72"),
    52 => (x"ed",x"d5",x"c1",x"87"),
    53 => (x"ec",x"d5",x"c1",x"4b"),
    54 => (x"50",x"f0",x"c0",x"48"),
    55 => (x"72",x"87",x"cd",x"c1"),
    56 => (x"e4",x"c0",x"02",x"9a"),
    57 => (x"4d",x"66",x"d4",x"87"),
    58 => (x"49",x"72",x"1e",x"72"),
    59 => (x"c2",x"cb",x"4a",x"75"),
    60 => (x"c5",x"4a",x"26",x"87"),
    61 => (x"53",x"11",x"81",x"dd"),
    62 => (x"4a",x"75",x"49",x"72"),
    63 => (x"70",x"87",x"f4",x"ca"),
    64 => (x"72",x"8c",x"c1",x"4a"),
    65 => (x"df",x"ff",x"05",x"9a"),
    66 => (x"ac",x"b7",x"c0",x"87"),
    67 => (x"c0",x"87",x"dd",x"06"),
    68 => (x"c5",x"02",x"66",x"e4"),
    69 => (x"4a",x"f0",x"c0",x"87"),
    70 => (x"e0",x"c0",x"87",x"c3"),
    71 => (x"97",x"0a",x"73",x"4a"),
    72 => (x"83",x"c1",x"0a",x"7a"),
    73 => (x"ac",x"b7",x"c0",x"8c"),
    74 => (x"87",x"e3",x"ff",x"01"),
    75 => (x"ab",x"ec",x"d5",x"c1"),
    76 => (x"d8",x"87",x"de",x"02"),
    77 => (x"66",x"dc",x"4c",x"66"),
    78 => (x"97",x"8b",x"c1",x"1e"),
    79 => (x"0f",x"74",x"49",x"6b"),
    80 => (x"48",x"6e",x"86",x"c4"),
    81 => (x"a6",x"c4",x"80",x"c1"),
    82 => (x"ec",x"d5",x"c1",x"58"),
    83 => (x"e5",x"ff",x"05",x"ab"),
    84 => (x"fc",x"48",x"6e",x"87"),
    85 => (x"26",x"4d",x"26",x"8e"),
    86 => (x"26",x"4b",x"26",x"4c"),
    87 => (x"32",x"31",x"30",x"4f"),
    88 => (x"36",x"35",x"34",x"33"),
    89 => (x"41",x"39",x"38",x"37"),
    90 => (x"45",x"44",x"43",x"42"),
    91 => (x"5e",x"0e",x"00",x"46"),
    92 => (x"0e",x"5d",x"5c",x"5b"),
    93 => (x"4d",x"ff",x"4b",x"71"),
    94 => (x"02",x"9c",x"4c",x"13"),
    95 => (x"85",x"c1",x"87",x"d7"),
    96 => (x"74",x"1e",x"66",x"d4"),
    97 => (x"0f",x"66",x"d4",x"49"),
    98 => (x"a8",x"74",x"86",x"c4"),
    99 => (x"13",x"87",x"c6",x"05"),
   100 => (x"e9",x"05",x"9c",x"4c"),
   101 => (x"26",x"48",x"75",x"87"),
   102 => (x"26",x"4c",x"26",x"4d"),
   103 => (x"0e",x"4f",x"26",x"4b"),
   104 => (x"5d",x"5c",x"5b",x"5e"),
   105 => (x"c4",x"86",x"e8",x"0e"),
   106 => (x"e8",x"c0",x"59",x"a6"),
   107 => (x"4c",x"c0",x"4d",x"66"),
   108 => (x"c0",x"48",x"a6",x"c8"),
   109 => (x"bf",x"97",x"6e",x"78"),
   110 => (x"c1",x"48",x"6e",x"4b"),
   111 => (x"58",x"a6",x"c4",x"80"),
   112 => (x"c6",x"02",x"9b",x"73"),
   113 => (x"66",x"c8",x"87",x"ce"),
   114 => (x"87",x"d6",x"c5",x"02"),
   115 => (x"c0",x"48",x"a6",x"cc"),
   116 => (x"c0",x"80",x"fc",x"78"),
   117 => (x"c0",x"4a",x"73",x"78"),
   118 => (x"c3",x"02",x"8a",x"e0"),
   119 => (x"8a",x"c3",x"87",x"c2"),
   120 => (x"87",x"fc",x"c2",x"02"),
   121 => (x"c2",x"02",x"8a",x"c2"),
   122 => (x"02",x"8a",x"87",x"e4"),
   123 => (x"c4",x"87",x"f1",x"c2"),
   124 => (x"eb",x"c2",x"02",x"8a"),
   125 => (x"02",x"8a",x"c2",x"87"),
   126 => (x"c3",x"87",x"e5",x"c2"),
   127 => (x"e7",x"c2",x"02",x"8a"),
   128 => (x"02",x"8a",x"d4",x"87"),
   129 => (x"8a",x"87",x"f4",x"c0"),
   130 => (x"87",x"ff",x"c0",x"02"),
   131 => (x"c0",x"02",x"8a",x"ca"),
   132 => (x"8a",x"c1",x"87",x"f1"),
   133 => (x"87",x"df",x"c1",x"02"),
   134 => (x"87",x"df",x"02",x"8a"),
   135 => (x"c1",x"02",x"8a",x"c8"),
   136 => (x"8a",x"c4",x"87",x"cd"),
   137 => (x"87",x"e3",x"c0",x"02"),
   138 => (x"c0",x"02",x"8a",x"c3"),
   139 => (x"8a",x"c2",x"87",x"e5"),
   140 => (x"c3",x"87",x"c8",x"02"),
   141 => (x"87",x"d3",x"02",x"8a"),
   142 => (x"cc",x"87",x"f9",x"c1"),
   143 => (x"78",x"ca",x"48",x"a6"),
   144 => (x"cc",x"87",x"d1",x"c2"),
   145 => (x"78",x"c2",x"48",x"a6"),
   146 => (x"cc",x"87",x"c9",x"c2"),
   147 => (x"78",x"d0",x"48",x"a6"),
   148 => (x"c0",x"87",x"c1",x"c2"),
   149 => (x"c0",x"1e",x"66",x"f0"),
   150 => (x"c4",x"1e",x"66",x"f0"),
   151 => (x"c4",x"4a",x"75",x"85"),
   152 => (x"fc",x"49",x"6a",x"8a"),
   153 => (x"86",x"c8",x"87",x"c8"),
   154 => (x"4c",x"a4",x"49",x"70"),
   155 => (x"c8",x"87",x"e5",x"c1"),
   156 => (x"78",x"c1",x"48",x"a6"),
   157 => (x"c0",x"87",x"dd",x"c1"),
   158 => (x"c4",x"1e",x"66",x"f0"),
   159 => (x"c4",x"4a",x"75",x"85"),
   160 => (x"c0",x"49",x"6a",x"8a"),
   161 => (x"c4",x"0f",x"66",x"f0"),
   162 => (x"c1",x"84",x"c1",x"86"),
   163 => (x"f0",x"c0",x"87",x"c6"),
   164 => (x"e5",x"c0",x"1e",x"66"),
   165 => (x"66",x"f0",x"c0",x"49"),
   166 => (x"c1",x"86",x"c4",x"0f"),
   167 => (x"87",x"f4",x"c0",x"84"),
   168 => (x"c1",x"48",x"a6",x"c8"),
   169 => (x"87",x"ec",x"c0",x"78"),
   170 => (x"c1",x"48",x"a6",x"d0"),
   171 => (x"c1",x"80",x"f8",x"78"),
   172 => (x"87",x"e0",x"c0",x"78"),
   173 => (x"06",x"ab",x"f0",x"c0"),
   174 => (x"f9",x"c0",x"87",x"da"),
   175 => (x"87",x"d4",x"03",x"ab"),
   176 => (x"ca",x"49",x"66",x"d4"),
   177 => (x"c0",x"4a",x"73",x"91"),
   178 => (x"a6",x"d4",x"8a",x"f0"),
   179 => (x"78",x"a1",x"72",x"48"),
   180 => (x"78",x"c1",x"80",x"f4"),
   181 => (x"c1",x"02",x"66",x"cc"),
   182 => (x"85",x"c4",x"87",x"e9"),
   183 => (x"89",x"c4",x"49",x"75"),
   184 => (x"78",x"69",x"48",x"a6"),
   185 => (x"05",x"ab",x"e4",x"c1"),
   186 => (x"66",x"c4",x"87",x"d8"),
   187 => (x"a8",x"b7",x"c0",x"48"),
   188 => (x"c0",x"87",x"cf",x"03"),
   189 => (x"fa",x"c1",x"49",x"ed"),
   190 => (x"48",x"66",x"c4",x"87"),
   191 => (x"c8",x"88",x"08",x"c0"),
   192 => (x"66",x"d0",x"58",x"a6"),
   193 => (x"1e",x"66",x"d8",x"1e"),
   194 => (x"1e",x"66",x"f8",x"c0"),
   195 => (x"1e",x"66",x"f8",x"c0"),
   196 => (x"d8",x"1e",x"66",x"dc"),
   197 => (x"df",x"f6",x"49",x"66"),
   198 => (x"70",x"86",x"d4",x"87"),
   199 => (x"c0",x"4c",x"a4",x"49"),
   200 => (x"e5",x"c0",x"87",x"e1"),
   201 => (x"87",x"cf",x"05",x"ab"),
   202 => (x"c0",x"48",x"a6",x"d0"),
   203 => (x"c0",x"80",x"c4",x"78"),
   204 => (x"c1",x"80",x"f4",x"78"),
   205 => (x"c0",x"87",x"cc",x"78"),
   206 => (x"73",x"1e",x"66",x"f0"),
   207 => (x"66",x"f0",x"c0",x"49"),
   208 => (x"6e",x"86",x"c4",x"0f"),
   209 => (x"6e",x"4b",x"bf",x"97"),
   210 => (x"c4",x"80",x"c1",x"48"),
   211 => (x"9b",x"73",x"58",x"a6"),
   212 => (x"87",x"f2",x"f9",x"05"),
   213 => (x"8e",x"e8",x"48",x"74"),
   214 => (x"4c",x"26",x"4d",x"26"),
   215 => (x"4f",x"26",x"4b",x"26"),
   216 => (x"cd",x"1e",x"c0",x"1e"),
   217 => (x"a6",x"d0",x"1e",x"f3"),
   218 => (x"49",x"66",x"d0",x"1e"),
   219 => (x"f4",x"87",x"f0",x"f8"),
   220 => (x"1e",x"4f",x"26",x"8e"),
   221 => (x"4a",x"71",x"86",x"fc"),
   222 => (x"69",x"49",x"c0",x"ff"),
   223 => (x"98",x"c0",x"c4",x"48"),
   224 => (x"70",x"58",x"a6",x"c4"),
   225 => (x"87",x"f3",x"02",x"98"),
   226 => (x"fc",x"48",x"79",x"72"),
   227 => (x"0e",x"4f",x"26",x"8e"),
   228 => (x"0e",x"5c",x"5b",x"5e"),
   229 => (x"4c",x"c0",x"4b",x"71"),
   230 => (x"02",x"9a",x"4a",x"13"),
   231 => (x"49",x"72",x"87",x"cd"),
   232 => (x"c1",x"87",x"d0",x"ff"),
   233 => (x"9a",x"4a",x"13",x"84"),
   234 => (x"74",x"87",x"f3",x"05"),
   235 => (x"26",x"4c",x"26",x"48"),
   236 => (x"1e",x"4f",x"26",x"4b"),
   237 => (x"9a",x"72",x"1e",x"73"),
   238 => (x"87",x"e7",x"c0",x"02"),
   239 => (x"4b",x"c1",x"48",x"c0"),
   240 => (x"d1",x"06",x"a9",x"72"),
   241 => (x"06",x"82",x"72",x"87"),
   242 => (x"83",x"73",x"87",x"c9"),
   243 => (x"f4",x"01",x"a9",x"72"),
   244 => (x"c1",x"87",x"c3",x"87"),
   245 => (x"a9",x"72",x"3a",x"b2"),
   246 => (x"80",x"73",x"89",x"03"),
   247 => (x"2b",x"2a",x"c1",x"07"),
   248 => (x"26",x"87",x"f3",x"05"),
   249 => (x"1e",x"4f",x"26",x"4b"),
   250 => (x"4d",x"c4",x"1e",x"75"),
   251 => (x"04",x"a1",x"b7",x"71"),
   252 => (x"81",x"c1",x"b9",x"ff"),
   253 => (x"72",x"07",x"bd",x"c3"),
   254 => (x"ff",x"04",x"a2",x"b7"),
   255 => (x"c1",x"82",x"c1",x"ba"),
   256 => (x"ee",x"fe",x"07",x"bd"),
   257 => (x"04",x"2d",x"c1",x"87"),
   258 => (x"80",x"c1",x"b8",x"ff"),
   259 => (x"ff",x"04",x"2d",x"07"),
   260 => (x"07",x"81",x"c1",x"b9"),
   261 => (x"4f",x"26",x"4d",x"26"),
   262 => (x"c0",x"c0",x"c1",x"1e"),
   263 => (x"b1",x"c0",x"c0",x"c0"),
   264 => (x"4f",x"26",x"0f",x"71"),
   265 => (x"d0",x"1e",x"73",x"1e"),
   266 => (x"c0",x"c0",x"c0",x"c0"),
   267 => (x"87",x"f9",x"f1",x"4b"),
   268 => (x"87",x"fe",x"0f",x"73"),
   269 => (x"4d",x"26",x"87",x"c4"),
   270 => (x"4b",x"26",x"4c",x"26"),
   271 => (x"c4",x"1e",x"4f",x"26"),
   272 => (x"df",x"c3",x"4a",x"66"),
   273 => (x"8a",x"f7",x"c0",x"9a"),
   274 => (x"03",x"aa",x"b7",x"c0"),
   275 => (x"e7",x"c0",x"87",x"c3"),
   276 => (x"72",x"31",x"c4",x"82"),
   277 => (x"26",x"48",x"71",x"b1"),
   278 => (x"5b",x"5e",x"0e",x"4f"),
   279 => (x"71",x"0e",x"5d",x"5c"),
   280 => (x"c0",x"c0",x"d0",x"4a"),
   281 => (x"c1",x"4d",x"c0",x"c0"),
   282 => (x"48",x"bf",x"fc",x"d5"),
   283 => (x"d6",x"c1",x"80",x"c1"),
   284 => (x"49",x"72",x"58",x"c0"),
   285 => (x"b9",x"81",x"c0",x"fe"),
   286 => (x"05",x"a9",x"d3",x"c1"),
   287 => (x"d5",x"c1",x"87",x"db"),
   288 => (x"78",x"c0",x"48",x"fc"),
   289 => (x"48",x"c0",x"d6",x"c1"),
   290 => (x"d6",x"c1",x"78",x"c0"),
   291 => (x"78",x"c0",x"48",x"c8"),
   292 => (x"48",x"cc",x"d6",x"c1"),
   293 => (x"e4",x"c6",x"78",x"c0"),
   294 => (x"fc",x"d5",x"c1",x"87"),
   295 => (x"a8",x"c1",x"48",x"bf"),
   296 => (x"87",x"f3",x"c0",x"05"),
   297 => (x"c0",x"fe",x"49",x"72"),
   298 => (x"1e",x"71",x"b9",x"81"),
   299 => (x"bf",x"cc",x"d6",x"c1"),
   300 => (x"87",x"ca",x"fe",x"49"),
   301 => (x"d6",x"c1",x"86",x"c4"),
   302 => (x"4b",x"70",x"58",x"d0"),
   303 => (x"06",x"ab",x"b7",x"c3"),
   304 => (x"48",x"ca",x"87",x"c6"),
   305 => (x"4b",x"70",x"88",x"73"),
   306 => (x"81",x"c1",x"49",x"73"),
   307 => (x"30",x"c1",x"48",x"71"),
   308 => (x"58",x"c8",x"d6",x"c1"),
   309 => (x"c1",x"87",x"e6",x"c5"),
   310 => (x"48",x"bf",x"cc",x"d6"),
   311 => (x"01",x"a8",x"b7",x"c9"),
   312 => (x"c1",x"87",x"da",x"c5"),
   313 => (x"48",x"bf",x"cc",x"d6"),
   314 => (x"06",x"a8",x"b7",x"c0"),
   315 => (x"c1",x"87",x"ce",x"c5"),
   316 => (x"48",x"bf",x"fc",x"d5"),
   317 => (x"01",x"a8",x"b7",x"c3"),
   318 => (x"49",x"72",x"87",x"d9"),
   319 => (x"b9",x"81",x"c0",x"fe"),
   320 => (x"d6",x"c1",x"1e",x"71"),
   321 => (x"fc",x"49",x"bf",x"c8"),
   322 => (x"86",x"c4",x"87",x"f4"),
   323 => (x"58",x"cc",x"d6",x"c1"),
   324 => (x"c1",x"87",x"ea",x"c4"),
   325 => (x"49",x"bf",x"c4",x"d6"),
   326 => (x"d5",x"c1",x"81",x"c3"),
   327 => (x"a9",x"b7",x"bf",x"fc"),
   328 => (x"72",x"87",x"df",x"04"),
   329 => (x"81",x"c0",x"fe",x"49"),
   330 => (x"c1",x"1e",x"71",x"b9"),
   331 => (x"49",x"bf",x"c0",x"d6"),
   332 => (x"c4",x"87",x"cb",x"fc"),
   333 => (x"c4",x"d6",x"c1",x"86"),
   334 => (x"d0",x"d6",x"c1",x"58"),
   335 => (x"c3",x"78",x"c1",x"48"),
   336 => (x"d6",x"c1",x"87",x"fb"),
   337 => (x"c0",x"48",x"bf",x"cc"),
   338 => (x"c2",x"06",x"a8",x"b7"),
   339 => (x"d6",x"c1",x"87",x"d2"),
   340 => (x"c3",x"48",x"bf",x"cc"),
   341 => (x"c2",x"01",x"a8",x"b7"),
   342 => (x"d6",x"c1",x"87",x"c6"),
   343 => (x"c1",x"49",x"bf",x"c8"),
   344 => (x"d5",x"c1",x"81",x"31"),
   345 => (x"a9",x"b7",x"bf",x"fc"),
   346 => (x"87",x"d6",x"c1",x"04"),
   347 => (x"c0",x"fe",x"49",x"72"),
   348 => (x"1e",x"71",x"b9",x"81"),
   349 => (x"bf",x"d4",x"d6",x"c1"),
   350 => (x"87",x"c2",x"fb",x"49"),
   351 => (x"d6",x"c1",x"86",x"c4"),
   352 => (x"d6",x"c1",x"58",x"d8"),
   353 => (x"c1",x"49",x"bf",x"d0"),
   354 => (x"d4",x"d6",x"c1",x"89"),
   355 => (x"a9",x"b7",x"c0",x"59"),
   356 => (x"87",x"e9",x"c2",x"03"),
   357 => (x"bf",x"c0",x"d6",x"c1"),
   358 => (x"c1",x"51",x"70",x"49"),
   359 => (x"49",x"bf",x"c0",x"d6"),
   360 => (x"d6",x"c1",x"81",x"c1"),
   361 => (x"d6",x"c1",x"59",x"c4"),
   362 => (x"a9",x"b7",x"bf",x"d8"),
   363 => (x"87",x"c9",x"c0",x"06"),
   364 => (x"48",x"d8",x"d6",x"c1"),
   365 => (x"bf",x"c0",x"d6",x"c1"),
   366 => (x"d0",x"d6",x"c1",x"78"),
   367 => (x"c1",x"78",x"c1",x"48"),
   368 => (x"d6",x"c1",x"87",x"fb"),
   369 => (x"c1",x"05",x"bf",x"d0"),
   370 => (x"d6",x"c1",x"87",x"f3"),
   371 => (x"c4",x"49",x"bf",x"d4"),
   372 => (x"d8",x"d6",x"c1",x"31"),
   373 => (x"c0",x"d6",x"c1",x"59"),
   374 => (x"79",x"97",x"09",x"bf"),
   375 => (x"87",x"dd",x"c1",x"09"),
   376 => (x"bf",x"cc",x"d6",x"c1"),
   377 => (x"a8",x"b7",x"c7",x"48"),
   378 => (x"87",x"d1",x"c1",x"04"),
   379 => (x"f4",x"fe",x"4c",x"c0"),
   380 => (x"c1",x"78",x"c1",x"48"),
   381 => (x"1e",x"bf",x"d8",x"d6"),
   382 => (x"c0",x"d9",x"1e",x"75"),
   383 => (x"87",x"e0",x"f5",x"1e"),
   384 => (x"d6",x"c1",x"86",x"cc"),
   385 => (x"d6",x"c1",x"5d",x"c4"),
   386 => (x"c1",x"48",x"bf",x"c0"),
   387 => (x"b7",x"bf",x"d8",x"d6"),
   388 => (x"db",x"c0",x"03",x"a8"),
   389 => (x"c0",x"d6",x"c1",x"87"),
   390 => (x"c1",x"84",x"bf",x"bf"),
   391 => (x"49",x"bf",x"c0",x"d6"),
   392 => (x"d6",x"c1",x"81",x"c4"),
   393 => (x"d6",x"c1",x"59",x"c4"),
   394 => (x"a9",x"b7",x"bf",x"d8"),
   395 => (x"87",x"e5",x"ff",x"04"),
   396 => (x"df",x"d9",x"1e",x"74"),
   397 => (x"87",x"e8",x"f4",x"1e"),
   398 => (x"e7",x"f7",x"86",x"c8"),
   399 => (x"87",x"f6",x"f7",x"87"),
   400 => (x"63",x"65",x"68",x"43"),
   401 => (x"6d",x"75",x"73",x"6b"),
   402 => (x"67",x"6e",x"69",x"6d"),
   403 => (x"6f",x"72",x"66",x"20"),
   404 => (x"64",x"25",x"20",x"6d"),
   405 => (x"20",x"6f",x"74",x"20"),
   406 => (x"2e",x"2e",x"64",x"25"),
   407 => (x"25",x"00",x"20",x"2e"),
   408 => (x"42",x"00",x"0a",x"64"),
   409 => (x"69",x"74",x"6f",x"6f"),
   410 => (x"2e",x"2e",x"67",x"6e"),
   411 => (x"42",x"00",x"0a",x"2e"),
   412 => (x"38",x"54",x"4f",x"4f"),
   413 => (x"42",x"20",x"32",x"33"),
   414 => (x"53",x"00",x"4e",x"49"),
   415 => (x"6f",x"62",x"20",x"44"),
   416 => (x"66",x"20",x"74",x"6f"),
   417 => (x"65",x"6c",x"69",x"61"),
   418 => (x"49",x"00",x"0a",x"64"),
   419 => (x"69",x"74",x"69",x"6e"),
   420 => (x"7a",x"69",x"6c",x"61"),
   421 => (x"20",x"67",x"6e",x"69"),
   422 => (x"63",x"20",x"44",x"53"),
   423 => (x"0a",x"64",x"72",x"61"),
   424 => (x"32",x"53",x"52",x"00"),
   425 => (x"62",x"20",x"32",x"33"),
   426 => (x"20",x"74",x"6f",x"6f"),
   427 => (x"72",x"70",x"20",x"2d"),
   428 => (x"20",x"73",x"73",x"65"),
   429 => (x"20",x"43",x"53",x"45"),
   430 => (x"62",x"20",x"6f",x"74"),
   431 => (x"20",x"74",x"6f",x"6f"),
   432 => (x"6d",x"6f",x"72",x"66"),
   433 => (x"2e",x"44",x"53",x"20"),
   434 => (x"5b",x"5e",x"0e",x"00"),
   435 => (x"1e",x"0e",x"5d",x"5c"),
   436 => (x"f2",x"49",x"cb",x"da"),
   437 => (x"ed",x"c0",x"87",x"f9"),
   438 => (x"98",x"70",x"87",x"d3"),
   439 => (x"c3",x"87",x"cc",x"02"),
   440 => (x"98",x"70",x"87",x"e0"),
   441 => (x"c1",x"87",x"c4",x"02"),
   442 => (x"c0",x"87",x"c2",x"4b"),
   443 => (x"5b",x"a6",x"c4",x"4b"),
   444 => (x"f2",x"49",x"e1",x"da"),
   445 => (x"d6",x"c1",x"87",x"d9"),
   446 => (x"78",x"c0",x"48",x"d8"),
   447 => (x"f1",x"49",x"ee",x"c0"),
   448 => (x"f4",x"c3",x"87",x"f1"),
   449 => (x"ff",x"4a",x"ff",x"c8"),
   450 => (x"49",x"4b",x"bf",x"c0"),
   451 => (x"02",x"99",x"c0",x"c8"),
   452 => (x"73",x"87",x"fd",x"c0"),
   453 => (x"9c",x"ff",x"c3",x"4c"),
   454 => (x"c0",x"05",x"ac",x"db"),
   455 => (x"02",x"6e",x"87",x"e8"),
   456 => (x"c0",x"d0",x"87",x"de"),
   457 => (x"1e",x"c0",x"c0",x"c0"),
   458 => (x"db",x"49",x"ef",x"d9"),
   459 => (x"86",x"c4",x"87",x"f7"),
   460 => (x"cb",x"02",x"98",x"70"),
   461 => (x"49",x"e3",x"d9",x"87"),
   462 => (x"f3",x"87",x"d4",x"f1"),
   463 => (x"87",x"c6",x"87",x"e6"),
   464 => (x"f1",x"49",x"fb",x"d9"),
   465 => (x"49",x"74",x"87",x"c9"),
   466 => (x"c3",x"87",x"ce",x"f4"),
   467 => (x"4a",x"c0",x"c9",x"f4"),
   468 => (x"8a",x"c1",x"49",x"72"),
   469 => (x"fe",x"05",x"99",x"71"),
   470 => (x"df",x"fe",x"87",x"ed"),
   471 => (x"d5",x"f3",x"26",x"87"),
   472 => (x"f9",x"e4",x"1e",x"87"),
   473 => (x"49",x"f2",x"c0",x"87"),
   474 => (x"d0",x"87",x"c8",x"f0"),
   475 => (x"c0",x"c0",x"c0",x"c0"),
   476 => (x"87",x"e4",x"f2",x"49"),
   477 => (x"4f",x"26",x"48",x"c0"),
   478 => (x"5c",x"5b",x"5e",x"0e"),
   479 => (x"c0",x"4b",x"71",x"0e"),
   480 => (x"48",x"66",x"d0",x"4c"),
   481 => (x"06",x"a8",x"b7",x"c0"),
   482 => (x"13",x"87",x"eb",x"c0"),
   483 => (x"82",x"c0",x"fe",x"4a"),
   484 => (x"97",x"66",x"cc",x"ba"),
   485 => (x"c0",x"fe",x"49",x"bf"),
   486 => (x"66",x"cc",x"b9",x"81"),
   487 => (x"d0",x"80",x"c1",x"48"),
   488 => (x"b7",x"71",x"58",x"a6"),
   489 => (x"87",x"c4",x"02",x"aa"),
   490 => (x"87",x"cc",x"48",x"c1"),
   491 => (x"66",x"d0",x"84",x"c1"),
   492 => (x"ff",x"04",x"ac",x"b7"),
   493 => (x"48",x"c0",x"87",x"d5"),
   494 => (x"4d",x"26",x"87",x"c2"),
   495 => (x"4b",x"26",x"4c",x"26"),
   496 => (x"5e",x"0e",x"4f",x"26"),
   497 => (x"0e",x"5d",x"5c",x"5b"),
   498 => (x"48",x"e4",x"de",x"c1"),
   499 => (x"ee",x"c0",x"78",x"c0"),
   500 => (x"fa",x"ee",x"49",x"c4"),
   501 => (x"dc",x"d6",x"c1",x"87"),
   502 => (x"c0",x"49",x"c0",x"1e"),
   503 => (x"c4",x"87",x"f3",x"ee"),
   504 => (x"05",x"98",x"70",x"86"),
   505 => (x"ea",x"c0",x"87",x"cc"),
   506 => (x"e2",x"ee",x"49",x"f0"),
   507 => (x"ca",x"48",x"c0",x"87"),
   508 => (x"ee",x"c0",x"87",x"fb"),
   509 => (x"d6",x"ee",x"49",x"d1"),
   510 => (x"c1",x"4b",x"c0",x"87"),
   511 => (x"c1",x"48",x"d0",x"df"),
   512 => (x"c0",x"1e",x"c8",x"78"),
   513 => (x"c1",x"1e",x"e8",x"ee"),
   514 => (x"fd",x"49",x"d2",x"d7"),
   515 => (x"86",x"c8",x"87",x"ea"),
   516 => (x"c6",x"05",x"98",x"70"),
   517 => (x"d0",x"df",x"c1",x"87"),
   518 => (x"c8",x"78",x"c0",x"48"),
   519 => (x"f1",x"ee",x"c0",x"1e"),
   520 => (x"ee",x"d7",x"c1",x"1e"),
   521 => (x"87",x"d0",x"fd",x"49"),
   522 => (x"98",x"70",x"86",x"c8"),
   523 => (x"c1",x"87",x"c6",x"05"),
   524 => (x"c0",x"48",x"d0",x"df"),
   525 => (x"d0",x"df",x"c1",x"78"),
   526 => (x"ee",x"c0",x"1e",x"bf"),
   527 => (x"df",x"ec",x"1e",x"fa"),
   528 => (x"c1",x"86",x"c8",x"87"),
   529 => (x"02",x"bf",x"d0",x"df"),
   530 => (x"c1",x"87",x"cb",x"c2"),
   531 => (x"48",x"4d",x"dc",x"d6"),
   532 => (x"4c",x"a0",x"fe",x"c6"),
   533 => (x"9f",x"da",x"de",x"c1"),
   534 => (x"c7",x"1e",x"49",x"bf"),
   535 => (x"48",x"49",x"a0",x"fe"),
   536 => (x"89",x"a0",x"c2",x"f8"),
   537 => (x"1e",x"d0",x"1e",x"71"),
   538 => (x"c0",x"1e",x"c0",x"c8"),
   539 => (x"eb",x"1e",x"e2",x"eb"),
   540 => (x"86",x"d4",x"87",x"ee"),
   541 => (x"69",x"49",x"a4",x"c8"),
   542 => (x"da",x"de",x"c1",x"4b"),
   543 => (x"c5",x"49",x"bf",x"9f"),
   544 => (x"05",x"a9",x"ea",x"d6"),
   545 => (x"c8",x"87",x"cd",x"c0"),
   546 => (x"49",x"6a",x"4a",x"a4"),
   547 => (x"87",x"e7",x"f2",x"c0"),
   548 => (x"87",x"db",x"4b",x"70"),
   549 => (x"49",x"a5",x"fe",x"c7"),
   550 => (x"ca",x"49",x"69",x"9f"),
   551 => (x"02",x"a9",x"d5",x"e9"),
   552 => (x"c0",x"87",x"cc",x"c0"),
   553 => (x"eb",x"49",x"c4",x"eb"),
   554 => (x"48",x"c0",x"87",x"e5"),
   555 => (x"73",x"87",x"fe",x"c7"),
   556 => (x"df",x"ec",x"c0",x"1e"),
   557 => (x"87",x"e8",x"ea",x"1e"),
   558 => (x"1e",x"dc",x"d6",x"c1"),
   559 => (x"eb",x"c0",x"49",x"73"),
   560 => (x"86",x"cc",x"87",x"d0"),
   561 => (x"c0",x"05",x"98",x"70"),
   562 => (x"48",x"c0",x"87",x"c5"),
   563 => (x"c0",x"87",x"de",x"c7"),
   564 => (x"ea",x"49",x"f7",x"ec"),
   565 => (x"ef",x"c0",x"87",x"f9"),
   566 => (x"c3",x"ea",x"1e",x"cd"),
   567 => (x"c0",x"1e",x"c8",x"87"),
   568 => (x"c1",x"1e",x"e5",x"ef"),
   569 => (x"fa",x"49",x"ee",x"d7"),
   570 => (x"86",x"cc",x"87",x"ce"),
   571 => (x"c0",x"05",x"98",x"70"),
   572 => (x"de",x"c1",x"87",x"c9"),
   573 => (x"78",x"c1",x"48",x"e4"),
   574 => (x"c8",x"87",x"e3",x"c0"),
   575 => (x"ee",x"ef",x"c0",x"1e"),
   576 => (x"d2",x"d7",x"c1",x"1e"),
   577 => (x"87",x"f0",x"f9",x"49"),
   578 => (x"98",x"70",x"86",x"c8"),
   579 => (x"87",x"ce",x"c0",x"02"),
   580 => (x"1e",x"de",x"ed",x"c0"),
   581 => (x"c4",x"87",x"c9",x"e9"),
   582 => (x"c6",x"48",x"c0",x"86"),
   583 => (x"de",x"c1",x"87",x"cf"),
   584 => (x"49",x"bf",x"97",x"da"),
   585 => (x"05",x"a9",x"d5",x"c1"),
   586 => (x"c1",x"87",x"cd",x"c0"),
   587 => (x"bf",x"97",x"db",x"de"),
   588 => (x"a9",x"ea",x"c2",x"49"),
   589 => (x"87",x"c5",x"c0",x"02"),
   590 => (x"f0",x"c5",x"48",x"c0"),
   591 => (x"dc",x"d6",x"c1",x"87"),
   592 => (x"c3",x"49",x"bf",x"97"),
   593 => (x"c0",x"02",x"a9",x"e9"),
   594 => (x"d6",x"c1",x"87",x"d2"),
   595 => (x"49",x"bf",x"97",x"dc"),
   596 => (x"02",x"a9",x"eb",x"c3"),
   597 => (x"c0",x"87",x"c5",x"c0"),
   598 => (x"87",x"d1",x"c5",x"48"),
   599 => (x"97",x"e7",x"d6",x"c1"),
   600 => (x"05",x"99",x"49",x"bf"),
   601 => (x"c1",x"87",x"cc",x"c0"),
   602 => (x"bf",x"97",x"e8",x"d6"),
   603 => (x"02",x"a9",x"c2",x"49"),
   604 => (x"c0",x"87",x"c5",x"c0"),
   605 => (x"87",x"f5",x"c4",x"48"),
   606 => (x"97",x"e9",x"d6",x"c1"),
   607 => (x"de",x"c1",x"48",x"bf"),
   608 => (x"49",x"70",x"58",x"e0"),
   609 => (x"c1",x"8a",x"c1",x"4a"),
   610 => (x"72",x"5a",x"e4",x"de"),
   611 => (x"c0",x"1e",x"71",x"1e"),
   612 => (x"e7",x"1e",x"f7",x"ef"),
   613 => (x"86",x"cc",x"87",x"ca"),
   614 => (x"97",x"ea",x"d6",x"c1"),
   615 => (x"81",x"73",x"49",x"bf"),
   616 => (x"97",x"eb",x"d6",x"c1"),
   617 => (x"32",x"c8",x"4a",x"bf"),
   618 => (x"48",x"f0",x"de",x"c1"),
   619 => (x"c1",x"78",x"a1",x"72"),
   620 => (x"bf",x"97",x"ec",x"d6"),
   621 => (x"c8",x"df",x"c1",x"48"),
   622 => (x"e4",x"de",x"c1",x"58"),
   623 => (x"dc",x"c2",x"02",x"bf"),
   624 => (x"c0",x"1e",x"c8",x"87"),
   625 => (x"c1",x"1e",x"fb",x"ed"),
   626 => (x"f6",x"49",x"ee",x"d7"),
   627 => (x"86",x"c8",x"87",x"ea"),
   628 => (x"c0",x"02",x"98",x"70"),
   629 => (x"48",x"c0",x"87",x"c5"),
   630 => (x"c1",x"87",x"d2",x"c3"),
   631 => (x"4a",x"bf",x"dc",x"de"),
   632 => (x"c1",x"30",x"c4",x"48"),
   633 => (x"c1",x"58",x"cc",x"df"),
   634 => (x"c1",x"5a",x"c4",x"df"),
   635 => (x"bf",x"97",x"c1",x"d7"),
   636 => (x"c1",x"31",x"c8",x"49"),
   637 => (x"bf",x"97",x"c0",x"d7"),
   638 => (x"c1",x"49",x"a1",x"4b"),
   639 => (x"bf",x"97",x"c2",x"d7"),
   640 => (x"73",x"33",x"d0",x"4b"),
   641 => (x"d7",x"c1",x"49",x"a1"),
   642 => (x"4b",x"bf",x"97",x"c3"),
   643 => (x"a1",x"73",x"33",x"d8"),
   644 => (x"d0",x"df",x"c1",x"49"),
   645 => (x"c4",x"df",x"c1",x"59"),
   646 => (x"de",x"c1",x"91",x"bf"),
   647 => (x"c1",x"81",x"bf",x"f0"),
   648 => (x"c1",x"59",x"f8",x"de"),
   649 => (x"bf",x"97",x"c9",x"d7"),
   650 => (x"c1",x"33",x"c8",x"4b"),
   651 => (x"bf",x"97",x"c8",x"d7"),
   652 => (x"c1",x"4b",x"a3",x"4c"),
   653 => (x"bf",x"97",x"ca",x"d7"),
   654 => (x"74",x"34",x"d0",x"4c"),
   655 => (x"d7",x"c1",x"4b",x"a3"),
   656 => (x"4c",x"bf",x"97",x"cb"),
   657 => (x"34",x"d8",x"9c",x"cf"),
   658 => (x"c1",x"4b",x"a3",x"74"),
   659 => (x"c2",x"5b",x"fc",x"de"),
   660 => (x"c1",x"92",x"73",x"8b"),
   661 => (x"72",x"48",x"fc",x"de"),
   662 => (x"ce",x"c1",x"78",x"a1"),
   663 => (x"ee",x"d6",x"c1",x"87"),
   664 => (x"c8",x"49",x"bf",x"97"),
   665 => (x"ed",x"d6",x"c1",x"31"),
   666 => (x"a1",x"4a",x"bf",x"97"),
   667 => (x"cc",x"df",x"c1",x"49"),
   668 => (x"c7",x"31",x"c5",x"59"),
   669 => (x"29",x"c9",x"81",x"ff"),
   670 => (x"59",x"c4",x"df",x"c1"),
   671 => (x"97",x"f3",x"d6",x"c1"),
   672 => (x"32",x"c8",x"4a",x"bf"),
   673 => (x"97",x"f2",x"d6",x"c1"),
   674 => (x"4a",x"a2",x"4b",x"bf"),
   675 => (x"5a",x"d0",x"df",x"c1"),
   676 => (x"bf",x"c4",x"df",x"c1"),
   677 => (x"f0",x"de",x"c1",x"92"),
   678 => (x"df",x"c1",x"82",x"bf"),
   679 => (x"de",x"c1",x"5a",x"c0"),
   680 => (x"78",x"c0",x"48",x"f8"),
   681 => (x"48",x"f4",x"de",x"c1"),
   682 => (x"c1",x"78",x"a1",x"72"),
   683 => (x"87",x"ca",x"f4",x"48"),
   684 => (x"64",x"61",x"65",x"52"),
   685 => (x"20",x"66",x"6f",x"20"),
   686 => (x"20",x"52",x"42",x"4d"),
   687 => (x"6c",x"69",x"61",x"66"),
   688 => (x"00",x"0a",x"64",x"65"),
   689 => (x"70",x"20",x"6f",x"4e"),
   690 => (x"69",x"74",x"72",x"61"),
   691 => (x"6e",x"6f",x"69",x"74"),
   692 => (x"67",x"69",x"73",x"20"),
   693 => (x"75",x"74",x"61",x"6e"),
   694 => (x"66",x"20",x"65",x"72"),
   695 => (x"64",x"6e",x"75",x"6f"),
   696 => (x"42",x"4d",x"00",x"0a"),
   697 => (x"7a",x"69",x"73",x"52"),
   698 => (x"25",x"20",x"3a",x"65"),
   699 => (x"70",x"20",x"2c",x"64"),
   700 => (x"69",x"74",x"72",x"61"),
   701 => (x"6e",x"6f",x"69",x"74"),
   702 => (x"65",x"7a",x"69",x"73"),
   703 => (x"64",x"25",x"20",x"3a"),
   704 => (x"66",x"6f",x"20",x"2c"),
   705 => (x"74",x"65",x"73",x"66"),
   706 => (x"20",x"66",x"6f",x"20"),
   707 => (x"3a",x"67",x"69",x"73"),
   708 => (x"2c",x"64",x"25",x"20"),
   709 => (x"67",x"69",x"73",x"20"),
   710 => (x"25",x"78",x"30",x"20"),
   711 => (x"52",x"00",x"0a",x"78"),
   712 => (x"69",x"64",x"61",x"65"),
   713 => (x"62",x"20",x"67",x"6e"),
   714 => (x"20",x"74",x"6f",x"6f"),
   715 => (x"74",x"63",x"65",x"73"),
   716 => (x"25",x"20",x"72",x"6f"),
   717 => (x"52",x"00",x"0a",x"64"),
   718 => (x"20",x"64",x"61",x"65"),
   719 => (x"74",x"6f",x"6f",x"62"),
   720 => (x"63",x"65",x"73",x"20"),
   721 => (x"20",x"72",x"6f",x"74"),
   722 => (x"6d",x"6f",x"72",x"66"),
   723 => (x"72",x"69",x"66",x"20"),
   724 => (x"70",x"20",x"74",x"73"),
   725 => (x"69",x"74",x"72",x"61"),
   726 => (x"6e",x"6f",x"69",x"74"),
   727 => (x"6e",x"55",x"00",x"0a"),
   728 => (x"70",x"70",x"75",x"73"),
   729 => (x"65",x"74",x"72",x"6f"),
   730 => (x"61",x"70",x"20",x"64"),
   731 => (x"74",x"69",x"74",x"72"),
   732 => (x"20",x"6e",x"6f",x"69"),
   733 => (x"65",x"70",x"79",x"74"),
   734 => (x"46",x"00",x"0d",x"21"),
   735 => (x"32",x"33",x"54",x"41"),
   736 => (x"00",x"20",x"20",x"20"),
   737 => (x"64",x"61",x"65",x"52"),
   738 => (x"20",x"67",x"6e",x"69"),
   739 => (x"0a",x"52",x"42",x"4d"),
   740 => (x"52",x"42",x"4d",x"00"),
   741 => (x"63",x"75",x"73",x"20"),
   742 => (x"73",x"73",x"65",x"63"),
   743 => (x"6c",x"6c",x"75",x"66"),
   744 => (x"65",x"72",x"20",x"79"),
   745 => (x"00",x"0a",x"64",x"61"),
   746 => (x"31",x"54",x"41",x"46"),
   747 => (x"20",x"20",x"20",x"36"),
   748 => (x"54",x"41",x"46",x"00"),
   749 => (x"20",x"20",x"32",x"33"),
   750 => (x"61",x"50",x"00",x"20"),
   751 => (x"74",x"69",x"74",x"72"),
   752 => (x"63",x"6e",x"6f",x"69"),
   753 => (x"74",x"6e",x"75",x"6f"),
   754 => (x"0a",x"64",x"25",x"20"),
   755 => (x"6e",x"75",x"48",x"00"),
   756 => (x"67",x"6e",x"69",x"74"),
   757 => (x"72",x"6f",x"66",x"20"),
   758 => (x"6c",x"69",x"66",x"20"),
   759 => (x"73",x"79",x"73",x"65"),
   760 => (x"0a",x"6d",x"65",x"74"),
   761 => (x"54",x"41",x"46",x"00"),
   762 => (x"20",x"20",x"32",x"33"),
   763 => (x"41",x"46",x"00",x"20"),
   764 => (x"20",x"36",x"31",x"54"),
   765 => (x"43",x"00",x"20",x"20"),
   766 => (x"74",x"73",x"75",x"6c"),
   767 => (x"73",x"20",x"72",x"65"),
   768 => (x"3a",x"65",x"7a",x"69"),
   769 => (x"2c",x"64",x"25",x"20"),
   770 => (x"75",x"6c",x"43",x"20"),
   771 => (x"72",x"65",x"74",x"73"),
   772 => (x"73",x"61",x"6d",x"20"),
   773 => (x"25",x"20",x"2c",x"6b"),
   774 => (x"4f",x"00",x"0a",x"64"),
   775 => (x"65",x"6e",x"65",x"70"),
   776 => (x"69",x"66",x"20",x"64"),
   777 => (x"20",x"2c",x"65",x"6c"),
   778 => (x"64",x"61",x"6f",x"6c"),
   779 => (x"2e",x"67",x"6e",x"69"),
   780 => (x"00",x"0a",x"2e",x"2e"),
   781 => (x"27",x"6e",x"61",x"43"),
   782 => (x"70",x"6f",x"20",x"74"),
   783 => (x"25",x"20",x"6e",x"65"),
   784 => (x"0e",x"00",x"0a",x"73"),
   785 => (x"5d",x"5c",x"5b",x"5e"),
   786 => (x"c1",x"4a",x"71",x"0e"),
   787 => (x"02",x"bf",x"e4",x"de"),
   788 => (x"4b",x"72",x"87",x"cc"),
   789 => (x"72",x"2b",x"b7",x"c7"),
   790 => (x"9d",x"ff",x"c1",x"4d"),
   791 => (x"4b",x"72",x"87",x"ca"),
   792 => (x"72",x"2b",x"b7",x"c8"),
   793 => (x"9d",x"ff",x"c3",x"4d"),
   794 => (x"1e",x"dc",x"d6",x"c1"),
   795 => (x"bf",x"f0",x"de",x"c1"),
   796 => (x"71",x"81",x"73",x"49"),
   797 => (x"c4",x"87",x"db",x"dc"),
   798 => (x"05",x"98",x"70",x"86"),
   799 => (x"48",x"c0",x"87",x"c5"),
   800 => (x"c1",x"87",x"e6",x"c0"),
   801 => (x"02",x"bf",x"e4",x"de"),
   802 => (x"49",x"75",x"87",x"d2"),
   803 => (x"d6",x"c1",x"91",x"c4"),
   804 => (x"4c",x"69",x"81",x"dc"),
   805 => (x"ff",x"ff",x"ff",x"cf"),
   806 => (x"87",x"cb",x"9c",x"ff"),
   807 => (x"91",x"c2",x"49",x"75"),
   808 => (x"81",x"dc",x"d6",x"c1"),
   809 => (x"74",x"4c",x"69",x"9f"),
   810 => (x"87",x"ce",x"ec",x"48"),
   811 => (x"5c",x"5b",x"5e",x"0e"),
   812 => (x"86",x"f4",x"0e",x"5d"),
   813 => (x"4b",x"c0",x"4c",x"71"),
   814 => (x"bf",x"f8",x"de",x"c1"),
   815 => (x"fc",x"de",x"c1",x"4d"),
   816 => (x"de",x"c1",x"7e",x"bf"),
   817 => (x"c9",x"02",x"bf",x"e4"),
   818 => (x"dc",x"de",x"c1",x"87"),
   819 => (x"32",x"c4",x"4a",x"bf"),
   820 => (x"df",x"c1",x"87",x"c7"),
   821 => (x"c4",x"4a",x"bf",x"c0"),
   822 => (x"5a",x"a6",x"c8",x"32"),
   823 => (x"c0",x"48",x"a6",x"c8"),
   824 => (x"48",x"66",x"c4",x"78"),
   825 => (x"c2",x"06",x"a8",x"c0"),
   826 => (x"66",x"c8",x"87",x"e7"),
   827 => (x"05",x"99",x"cf",x"49"),
   828 => (x"d6",x"c1",x"87",x"d9"),
   829 => (x"66",x"c4",x"1e",x"dc"),
   830 => (x"80",x"c1",x"48",x"49"),
   831 => (x"71",x"58",x"a6",x"c8"),
   832 => (x"c4",x"87",x"cf",x"da"),
   833 => (x"dc",x"d6",x"c1",x"86"),
   834 => (x"c0",x"87",x"c3",x"4b"),
   835 => (x"6b",x"97",x"83",x"e0"),
   836 => (x"c1",x"02",x"99",x"49"),
   837 => (x"6b",x"97",x"87",x"ec"),
   838 => (x"a9",x"e5",x"c3",x"49"),
   839 => (x"87",x"e2",x"c1",x"02"),
   840 => (x"97",x"49",x"a3",x"cb"),
   841 => (x"99",x"d8",x"49",x"69"),
   842 => (x"87",x"d6",x"c1",x"05"),
   843 => (x"d9",x"ff",x"49",x"73"),
   844 => (x"1e",x"cb",x"87",x"dd"),
   845 => (x"1e",x"66",x"e0",x"c0"),
   846 => (x"fb",x"e8",x"49",x"73"),
   847 => (x"70",x"86",x"c8",x"87"),
   848 => (x"fd",x"c0",x"05",x"98"),
   849 => (x"4a",x"a3",x"dc",x"87"),
   850 => (x"6a",x"49",x"a4",x"c4"),
   851 => (x"4a",x"a3",x"da",x"79"),
   852 => (x"9f",x"49",x"a4",x"c8"),
   853 => (x"c4",x"79",x"48",x"6a"),
   854 => (x"de",x"c1",x"59",x"a6"),
   855 => (x"cf",x"02",x"bf",x"e4"),
   856 => (x"49",x"a3",x"d4",x"87"),
   857 => (x"4a",x"49",x"69",x"9f"),
   858 => (x"9a",x"ff",x"ff",x"c0"),
   859 => (x"87",x"c2",x"32",x"d0"),
   860 => (x"48",x"72",x"4a",x"c0"),
   861 => (x"6e",x"80",x"bf",x"6e"),
   862 => (x"c0",x"08",x"78",x"08"),
   863 => (x"c1",x"48",x"c1",x"7c"),
   864 => (x"66",x"c8",x"87",x"c1"),
   865 => (x"cc",x"80",x"c1",x"48"),
   866 => (x"66",x"c4",x"58",x"a6"),
   867 => (x"d9",x"fd",x"04",x"a8"),
   868 => (x"e4",x"de",x"c1",x"87"),
   869 => (x"e8",x"c0",x"02",x"bf"),
   870 => (x"fa",x"49",x"75",x"87"),
   871 => (x"4d",x"70",x"87",x"e5"),
   872 => (x"ff",x"ff",x"cf",x"49"),
   873 => (x"a9",x"99",x"f8",x"ff"),
   874 => (x"75",x"87",x"d6",x"02"),
   875 => (x"c1",x"89",x"c2",x"49"),
   876 => (x"91",x"bf",x"dc",x"de"),
   877 => (x"bf",x"f4",x"de",x"c1"),
   878 => (x"c4",x"80",x"71",x"48"),
   879 => (x"db",x"fc",x"58",x"a6"),
   880 => (x"f4",x"48",x"c0",x"87"),
   881 => (x"87",x"f2",x"e7",x"8e"),
   882 => (x"71",x"1e",x"73",x"1e"),
   883 => (x"c1",x"49",x"6a",x"4a"),
   884 => (x"c1",x"7a",x"71",x"81"),
   885 => (x"99",x"bf",x"e0",x"de"),
   886 => (x"c8",x"87",x"cb",x"05"),
   887 => (x"49",x"6b",x"4b",x"a2"),
   888 => (x"70",x"87",x"e0",x"f9"),
   889 => (x"48",x"c1",x"7b",x"49"),
   890 => (x"1e",x"87",x"d3",x"e7"),
   891 => (x"4b",x"71",x"1e",x"73"),
   892 => (x"bf",x"f4",x"de",x"c1"),
   893 => (x"4a",x"a3",x"c8",x"49"),
   894 => (x"8a",x"c2",x"4a",x"6a"),
   895 => (x"bf",x"dc",x"de",x"c1"),
   896 => (x"49",x"a1",x"72",x"92"),
   897 => (x"bf",x"e0",x"de",x"c1"),
   898 => (x"72",x"9a",x"6b",x"4a"),
   899 => (x"66",x"c8",x"49",x"a1"),
   900 => (x"fd",x"d5",x"71",x"1e"),
   901 => (x"70",x"86",x"c4",x"87"),
   902 => (x"87",x"c4",x"05",x"98"),
   903 => (x"87",x"c2",x"48",x"c0"),
   904 => (x"d9",x"e6",x"48",x"c1"),
   905 => (x"5b",x"5e",x"0e",x"87"),
   906 => (x"71",x"0e",x"5d",x"5c"),
   907 => (x"df",x"c1",x"1e",x"4b"),
   908 => (x"f7",x"f9",x"49",x"d4"),
   909 => (x"70",x"86",x"c4",x"87"),
   910 => (x"ce",x"c1",x"02",x"98"),
   911 => (x"d8",x"df",x"c1",x"87"),
   912 => (x"ff",x"c7",x"49",x"bf"),
   913 => (x"71",x"29",x"c9",x"81"),
   914 => (x"c0",x"4c",x"c0",x"4d"),
   915 => (x"ff",x"49",x"db",x"f0"),
   916 => (x"c0",x"87",x"fc",x"d4"),
   917 => (x"c1",x"06",x"ad",x"b7"),
   918 => (x"66",x"d0",x"87",x"c1"),
   919 => (x"d4",x"df",x"c1",x"1e"),
   920 => (x"87",x"c7",x"fe",x"49"),
   921 => (x"98",x"70",x"86",x"c4"),
   922 => (x"c0",x"87",x"c5",x"05"),
   923 => (x"87",x"ed",x"c0",x"48"),
   924 => (x"49",x"d4",x"df",x"c1"),
   925 => (x"d0",x"87",x"d1",x"fd"),
   926 => (x"c0",x"c8",x"48",x"66"),
   927 => (x"58",x"a6",x"d4",x"80"),
   928 => (x"b7",x"75",x"84",x"c1"),
   929 => (x"d1",x"ff",x"04",x"ac"),
   930 => (x"73",x"87",x"d0",x"87"),
   931 => (x"f4",x"f0",x"c0",x"1e"),
   932 => (x"cb",x"d3",x"ff",x"1e"),
   933 => (x"c0",x"86",x"c8",x"87"),
   934 => (x"c1",x"87",x"c2",x"48"),
   935 => (x"87",x"da",x"e4",x"48"),
   936 => (x"ff",x"86",x"e8",x"1e"),
   937 => (x"ff",x"c3",x"4a",x"d4"),
   938 => (x"c3",x"49",x"6a",x"7a"),
   939 => (x"48",x"6a",x"7a",x"ff"),
   940 => (x"a6",x"c4",x"30",x"c8"),
   941 => (x"59",x"a6",x"c8",x"58"),
   942 => (x"ff",x"c3",x"b1",x"6e"),
   943 => (x"d0",x"48",x"6a",x"7a"),
   944 => (x"58",x"a6",x"cc",x"30"),
   945 => (x"c8",x"59",x"a6",x"d0"),
   946 => (x"ff",x"c3",x"b1",x"66"),
   947 => (x"d8",x"48",x"6a",x"7a"),
   948 => (x"58",x"a6",x"d4",x"30"),
   949 => (x"d0",x"59",x"a6",x"d8"),
   950 => (x"48",x"71",x"b1",x"66"),
   951 => (x"4f",x"26",x"8e",x"e8"),
   952 => (x"ff",x"86",x"f4",x"1e"),
   953 => (x"ff",x"c3",x"4a",x"d4"),
   954 => (x"c3",x"49",x"6a",x"7a"),
   955 => (x"48",x"71",x"7a",x"ff"),
   956 => (x"a6",x"c4",x"30",x"c8"),
   957 => (x"6e",x"49",x"6a",x"58"),
   958 => (x"7a",x"ff",x"c3",x"b1"),
   959 => (x"30",x"c8",x"48",x"71"),
   960 => (x"49",x"6a",x"58",x"a6"),
   961 => (x"c3",x"b1",x"66",x"c4"),
   962 => (x"48",x"71",x"7a",x"ff"),
   963 => (x"a6",x"cc",x"30",x"c8"),
   964 => (x"c8",x"49",x"6a",x"58"),
   965 => (x"48",x"71",x"b1",x"66"),
   966 => (x"4f",x"26",x"8e",x"f4"),
   967 => (x"5c",x"5b",x"5e",x"0e"),
   968 => (x"4d",x"71",x"0e",x"5d"),
   969 => (x"75",x"4c",x"d4",x"ff"),
   970 => (x"98",x"ff",x"c3",x"48"),
   971 => (x"df",x"c1",x"7c",x"70"),
   972 => (x"c8",x"05",x"bf",x"e4"),
   973 => (x"48",x"66",x"d0",x"87"),
   974 => (x"a6",x"d4",x"30",x"c9"),
   975 => (x"49",x"66",x"d0",x"58"),
   976 => (x"48",x"71",x"29",x"d8"),
   977 => (x"70",x"98",x"ff",x"c3"),
   978 => (x"49",x"66",x"d0",x"7c"),
   979 => (x"48",x"71",x"29",x"d0"),
   980 => (x"70",x"98",x"ff",x"c3"),
   981 => (x"49",x"66",x"d0",x"7c"),
   982 => (x"48",x"71",x"29",x"c8"),
   983 => (x"70",x"98",x"ff",x"c3"),
   984 => (x"48",x"66",x"d0",x"7c"),
   985 => (x"70",x"98",x"ff",x"c3"),
   986 => (x"d0",x"49",x"75",x"7c"),
   987 => (x"c3",x"48",x"71",x"29"),
   988 => (x"7c",x"70",x"98",x"ff"),
   989 => (x"f0",x"c9",x"4b",x"6c"),
   990 => (x"ff",x"c3",x"4a",x"ff"),
   991 => (x"87",x"d1",x"05",x"ab"),
   992 => (x"71",x"49",x"ff",x"c3"),
   993 => (x"c1",x"4b",x"6c",x"7c"),
   994 => (x"87",x"c5",x"02",x"8a"),
   995 => (x"f2",x"02",x"ab",x"71"),
   996 => (x"26",x"48",x"73",x"87"),
   997 => (x"26",x"4c",x"26",x"4d"),
   998 => (x"1e",x"4f",x"26",x"4b"),
   999 => (x"d4",x"ff",x"49",x"c0"),
  1000 => (x"78",x"ff",x"c3",x"48"),
  1001 => (x"c8",x"c3",x"81",x"c1"),
  1002 => (x"f1",x"04",x"a9",x"b7"),
  1003 => (x"0e",x"4f",x"26",x"87"),
  1004 => (x"5d",x"5c",x"5b",x"5e"),
  1005 => (x"f0",x"ff",x"c0",x"0e"),
  1006 => (x"c1",x"4d",x"f7",x"c1"),
  1007 => (x"c0",x"c0",x"c0",x"c0"),
  1008 => (x"d6",x"ff",x"4b",x"c0"),
  1009 => (x"df",x"f8",x"c4",x"87"),
  1010 => (x"75",x"1e",x"c0",x"4c"),
  1011 => (x"87",x"cc",x"fd",x"49"),
  1012 => (x"a8",x"c1",x"86",x"c4"),
  1013 => (x"87",x"e5",x"c0",x"05"),
  1014 => (x"c3",x"48",x"d4",x"ff"),
  1015 => (x"1e",x"73",x"78",x"ff"),
  1016 => (x"c1",x"f0",x"e1",x"c0"),
  1017 => (x"f3",x"fc",x"49",x"e9"),
  1018 => (x"70",x"86",x"c4",x"87"),
  1019 => (x"87",x"ca",x"05",x"98"),
  1020 => (x"c3",x"48",x"d4",x"ff"),
  1021 => (x"48",x"c1",x"78",x"ff"),
  1022 => (x"de",x"fe",x"87",x"cb"),
  1023 => (x"05",x"8c",x"c1",x"87"),
  1024 => (x"c0",x"87",x"c6",x"ff"),
  1025 => (x"26",x"4d",x"26",x"48"),
  1026 => (x"26",x"4b",x"26",x"4c"),
  1027 => (x"5b",x"5e",x"0e",x"4f"),
  1028 => (x"ff",x"c0",x"0e",x"5c"),
  1029 => (x"4c",x"c1",x"c1",x"f0"),
  1030 => (x"c3",x"48",x"d4",x"ff"),
  1031 => (x"c1",x"c1",x"78",x"ff"),
  1032 => (x"cd",x"ff",x"49",x"d1"),
  1033 => (x"4b",x"d3",x"87",x"e9"),
  1034 => (x"49",x"74",x"1e",x"c0"),
  1035 => (x"c4",x"87",x"ed",x"fb"),
  1036 => (x"05",x"98",x"70",x"86"),
  1037 => (x"d4",x"ff",x"87",x"ca"),
  1038 => (x"78",x"ff",x"c3",x"48"),
  1039 => (x"87",x"cb",x"48",x"c1"),
  1040 => (x"c1",x"87",x"d8",x"fd"),
  1041 => (x"df",x"ff",x"05",x"8b"),
  1042 => (x"26",x"48",x"c0",x"87"),
  1043 => (x"26",x"4b",x"26",x"4c"),
  1044 => (x"44",x"4d",x"43",x"4f"),
  1045 => (x"44",x"4d",x"43",x"00"),
  1046 => (x"25",x"20",x"38",x"35"),
  1047 => (x"20",x"20",x"0a",x"64"),
  1048 => (x"44",x"4d",x"43",x"00"),
  1049 => (x"32",x"5f",x"38",x"35"),
  1050 => (x"0a",x"64",x"25",x"20"),
  1051 => (x"43",x"00",x"20",x"20"),
  1052 => (x"38",x"35",x"44",x"4d"),
  1053 => (x"0a",x"64",x"25",x"20"),
  1054 => (x"53",x"00",x"20",x"20"),
  1055 => (x"20",x"43",x"48",x"44"),
  1056 => (x"74",x"69",x"6e",x"49"),
  1057 => (x"69",x"6c",x"61",x"69"),
  1058 => (x"69",x"74",x"61",x"7a"),
  1059 => (x"65",x"20",x"6e",x"6f"),
  1060 => (x"72",x"6f",x"72",x"72"),
  1061 => (x"63",x"00",x"0a",x"21"),
  1062 => (x"43",x"5f",x"64",x"6d"),
  1063 => (x"20",x"38",x"44",x"4d"),
  1064 => (x"70",x"73",x"65",x"72"),
  1065 => (x"65",x"73",x"6e",x"6f"),
  1066 => (x"64",x"25",x"20",x"3a"),
  1067 => (x"45",x"49",x"00",x"0a"),
  1068 => (x"53",x"00",x"52",x"52"),
  1069 => (x"53",x"00",x"49",x"50"),
  1070 => (x"61",x"63",x"20",x"44"),
  1071 => (x"73",x"20",x"64",x"72"),
  1072 => (x"20",x"65",x"7a",x"69"),
  1073 => (x"25",x"20",x"73",x"69"),
  1074 => (x"57",x"00",x"0a",x"64"),
  1075 => (x"65",x"74",x"69",x"72"),
  1076 => (x"69",x"61",x"66",x"20"),
  1077 => (x"0a",x"64",x"65",x"6c"),
  1078 => (x"61",x"65",x"52",x"00"),
  1079 => (x"6f",x"63",x"20",x"64"),
  1080 => (x"6e",x"61",x"6d",x"6d"),
  1081 => (x"61",x"66",x"20",x"64"),
  1082 => (x"64",x"65",x"6c",x"69"),
  1083 => (x"20",x"74",x"61",x"20"),
  1084 => (x"28",x"20",x"64",x"25"),
  1085 => (x"0a",x"29",x"64",x"25"),
  1086 => (x"73",x"5f",x"63",x"00"),
  1087 => (x"5f",x"65",x"7a",x"69"),
  1088 => (x"74",x"6c",x"75",x"6d"),
  1089 => (x"64",x"25",x"20",x"3a"),
  1090 => (x"65",x"72",x"20",x"2c"),
  1091 => (x"62",x"5f",x"64",x"61"),
  1092 => (x"65",x"6c",x"5f",x"6c"),
  1093 => (x"25",x"20",x"3a",x"6e"),
  1094 => (x"63",x"20",x"2c",x"64"),
  1095 => (x"65",x"7a",x"69",x"73"),
  1096 => (x"64",x"25",x"20",x"3a"),
  1097 => (x"75",x"4d",x"00",x"0a"),
  1098 => (x"25",x"20",x"74",x"6c"),
  1099 => (x"25",x"00",x"0a",x"64"),
  1100 => (x"6c",x"62",x"20",x"64"),
  1101 => (x"73",x"6b",x"63",x"6f"),
  1102 => (x"20",x"66",x"6f",x"20"),
  1103 => (x"65",x"7a",x"69",x"73"),
  1104 => (x"0a",x"64",x"25",x"20"),
  1105 => (x"20",x"64",x"25",x"00"),
  1106 => (x"63",x"6f",x"6c",x"62"),
  1107 => (x"6f",x"20",x"73",x"6b"),
  1108 => (x"31",x"35",x"20",x"66"),
  1109 => (x"79",x"62",x"20",x"32"),
  1110 => (x"0a",x"73",x"65",x"74"),
  1111 => (x"5b",x"5e",x"0e",x"00"),
  1112 => (x"ff",x"0e",x"5d",x"5c"),
  1113 => (x"f2",x"f8",x"4c",x"d4"),
  1114 => (x"1e",x"ea",x"c6",x"87"),
  1115 => (x"c1",x"f0",x"e1",x"c0"),
  1116 => (x"e7",x"f6",x"49",x"c8"),
  1117 => (x"73",x"4b",x"70",x"87"),
  1118 => (x"d7",x"c2",x"c1",x"1e"),
  1119 => (x"df",x"c7",x"ff",x"1e"),
  1120 => (x"c1",x"86",x"cc",x"87"),
  1121 => (x"87",x"c8",x"02",x"ab"),
  1122 => (x"c0",x"87",x"c2",x"fa"),
  1123 => (x"87",x"d5",x"c2",x"48"),
  1124 => (x"70",x"87",x"cd",x"f5"),
  1125 => (x"ff",x"ff",x"cf",x"49"),
  1126 => (x"a9",x"ea",x"c6",x"99"),
  1127 => (x"f9",x"87",x"c8",x"02"),
  1128 => (x"48",x"c0",x"87",x"eb"),
  1129 => (x"c3",x"87",x"fe",x"c1"),
  1130 => (x"f1",x"c0",x"7c",x"ff"),
  1131 => (x"87",x"ff",x"f7",x"4d"),
  1132 => (x"c1",x"02",x"98",x"70"),
  1133 => (x"1e",x"c0",x"87",x"d4"),
  1134 => (x"c1",x"f0",x"ff",x"c0"),
  1135 => (x"db",x"f5",x"49",x"fa"),
  1136 => (x"70",x"86",x"c4",x"87"),
  1137 => (x"05",x"9b",x"73",x"4b"),
  1138 => (x"73",x"87",x"f3",x"c0"),
  1139 => (x"d5",x"c1",x"c1",x"1e"),
  1140 => (x"cb",x"c6",x"ff",x"1e"),
  1141 => (x"7c",x"ff",x"c3",x"87"),
  1142 => (x"1e",x"73",x"4b",x"6c"),
  1143 => (x"1e",x"e1",x"c1",x"c1"),
  1144 => (x"87",x"fc",x"c5",x"ff"),
  1145 => (x"ff",x"c3",x"86",x"d0"),
  1146 => (x"7c",x"7c",x"7c",x"7c"),
  1147 => (x"c0",x"c1",x"49",x"73"),
  1148 => (x"87",x"c5",x"02",x"99"),
  1149 => (x"ec",x"c0",x"48",x"c1"),
  1150 => (x"c0",x"48",x"c0",x"87"),
  1151 => (x"1e",x"73",x"87",x"e7"),
  1152 => (x"1e",x"ef",x"c1",x"c1"),
  1153 => (x"87",x"d8",x"c5",x"ff"),
  1154 => (x"ad",x"c2",x"86",x"c8"),
  1155 => (x"c1",x"87",x"ce",x"05"),
  1156 => (x"ff",x"1e",x"fb",x"c1"),
  1157 => (x"c4",x"87",x"c9",x"c5"),
  1158 => (x"c8",x"48",x"c0",x"86"),
  1159 => (x"05",x"8d",x"c1",x"87"),
  1160 => (x"c0",x"87",x"ca",x"fe"),
  1161 => (x"26",x"4d",x"26",x"48"),
  1162 => (x"26",x"4b",x"26",x"4c"),
  1163 => (x"5b",x"5e",x"0e",x"4f"),
  1164 => (x"fc",x"0e",x"5d",x"5c"),
  1165 => (x"4c",x"d0",x"ff",x"86"),
  1166 => (x"4b",x"c0",x"c0",x"c8"),
  1167 => (x"48",x"e4",x"df",x"c1"),
  1168 => (x"c2",x"c1",x"78",x"c1"),
  1169 => (x"c5",x"ff",x"49",x"f3"),
  1170 => (x"4d",x"c7",x"87",x"c5"),
  1171 => (x"98",x"73",x"48",x"6c"),
  1172 => (x"6e",x"58",x"a6",x"c4"),
  1173 => (x"6c",x"87",x"cb",x"02"),
  1174 => (x"c4",x"98",x"73",x"48"),
  1175 => (x"05",x"6e",x"58",x"a6"),
  1176 => (x"7c",x"c0",x"87",x"f5"),
  1177 => (x"6c",x"87",x"f4",x"f4"),
  1178 => (x"c4",x"98",x"73",x"48"),
  1179 => (x"02",x"6e",x"58",x"a6"),
  1180 => (x"48",x"6c",x"87",x"cb"),
  1181 => (x"a6",x"c4",x"98",x"73"),
  1182 => (x"f5",x"05",x"6e",x"58"),
  1183 => (x"c0",x"7c",x"c1",x"87"),
  1184 => (x"d0",x"e5",x"c0",x"1e"),
  1185 => (x"f2",x"49",x"c0",x"c1"),
  1186 => (x"86",x"c4",x"87",x"d2"),
  1187 => (x"c2",x"05",x"a8",x"c1"),
  1188 => (x"c2",x"4d",x"c1",x"87"),
  1189 => (x"87",x"cd",x"05",x"ad"),
  1190 => (x"49",x"ee",x"c2",x"c1"),
  1191 => (x"87",x"ef",x"c3",x"ff"),
  1192 => (x"de",x"c1",x"48",x"c0"),
  1193 => (x"05",x"8d",x"c1",x"87"),
  1194 => (x"fa",x"87",x"e1",x"fe"),
  1195 => (x"df",x"c1",x"87",x"ef"),
  1196 => (x"df",x"c1",x"58",x"e8"),
  1197 => (x"cd",x"05",x"bf",x"e4"),
  1198 => (x"c0",x"1e",x"c1",x"87"),
  1199 => (x"d0",x"c1",x"f0",x"ff"),
  1200 => (x"87",x"d8",x"f1",x"49"),
  1201 => (x"d4",x"ff",x"86",x"c4"),
  1202 => (x"78",x"ff",x"c3",x"48"),
  1203 => (x"c1",x"87",x"d6",x"c5"),
  1204 => (x"c1",x"58",x"ec",x"df"),
  1205 => (x"1e",x"bf",x"e8",x"df"),
  1206 => (x"1e",x"f7",x"c2",x"c1"),
  1207 => (x"87",x"c0",x"c2",x"ff"),
  1208 => (x"48",x"6c",x"86",x"c8"),
  1209 => (x"a6",x"c4",x"98",x"73"),
  1210 => (x"cc",x"02",x"6e",x"58"),
  1211 => (x"73",x"48",x"6c",x"87"),
  1212 => (x"58",x"a6",x"c4",x"98"),
  1213 => (x"f4",x"ff",x"05",x"6e"),
  1214 => (x"ff",x"7c",x"c0",x"87"),
  1215 => (x"ff",x"c3",x"48",x"d4"),
  1216 => (x"fc",x"48",x"c1",x"78"),
  1217 => (x"26",x"4d",x"26",x"8e"),
  1218 => (x"26",x"4b",x"26",x"4c"),
  1219 => (x"5b",x"5e",x"0e",x"4f"),
  1220 => (x"71",x"0e",x"5d",x"5c"),
  1221 => (x"4d",x"d4",x"ff",x"4b"),
  1222 => (x"c0",x"4c",x"66",x"d0"),
  1223 => (x"cd",x"ee",x"c5",x"4a"),
  1224 => (x"ff",x"c3",x"49",x"df"),
  1225 => (x"c3",x"48",x"6d",x"7d"),
  1226 => (x"c1",x"05",x"a8",x"fe"),
  1227 => (x"df",x"c1",x"87",x"d1"),
  1228 => (x"78",x"c0",x"48",x"e0"),
  1229 => (x"04",x"ac",x"b7",x"c4"),
  1230 => (x"e3",x"ed",x"87",x"db"),
  1231 => (x"71",x"49",x"70",x"87"),
  1232 => (x"c1",x"83",x"c4",x"7b"),
  1233 => (x"48",x"bf",x"e0",x"df"),
  1234 => (x"df",x"c1",x"80",x"71"),
  1235 => (x"8c",x"c4",x"58",x"e4"),
  1236 => (x"e5",x"03",x"ac",x"b7"),
  1237 => (x"ac",x"b7",x"c0",x"87"),
  1238 => (x"87",x"e0",x"c0",x"06"),
  1239 => (x"6d",x"7d",x"ff",x"c3"),
  1240 => (x"97",x"09",x"73",x"49"),
  1241 => (x"83",x"c1",x"09",x"79"),
  1242 => (x"bf",x"e0",x"df",x"c1"),
  1243 => (x"c1",x"80",x"71",x"48"),
  1244 => (x"c1",x"58",x"e4",x"df"),
  1245 => (x"ac",x"b7",x"c0",x"8c"),
  1246 => (x"87",x"e0",x"ff",x"01"),
  1247 => (x"c1",x"4a",x"49",x"c1"),
  1248 => (x"dd",x"fe",x"05",x"89"),
  1249 => (x"7d",x"ff",x"c3",x"87"),
  1250 => (x"4d",x"26",x"48",x"72"),
  1251 => (x"4b",x"26",x"4c",x"26"),
  1252 => (x"5e",x"0e",x"4f",x"26"),
  1253 => (x"0e",x"5d",x"5c",x"5b"),
  1254 => (x"4d",x"71",x"86",x"f8"),
  1255 => (x"c8",x"4c",x"d0",x"ff"),
  1256 => (x"c0",x"4b",x"c0",x"c0"),
  1257 => (x"48",x"d4",x"ff",x"7e"),
  1258 => (x"6c",x"78",x"ff",x"c3"),
  1259 => (x"c8",x"98",x"73",x"48"),
  1260 => (x"66",x"c4",x"58",x"a6"),
  1261 => (x"6c",x"87",x"cc",x"02"),
  1262 => (x"c8",x"98",x"73",x"48"),
  1263 => (x"66",x"c4",x"58",x"a6"),
  1264 => (x"c4",x"87",x"f4",x"05"),
  1265 => (x"d4",x"ff",x"7c",x"c1"),
  1266 => (x"78",x"ff",x"c3",x"48"),
  1267 => (x"ff",x"c0",x"1e",x"75"),
  1268 => (x"49",x"d1",x"c1",x"f0"),
  1269 => (x"c4",x"87",x"c5",x"ed"),
  1270 => (x"72",x"4a",x"70",x"86"),
  1271 => (x"87",x"d1",x"02",x"9a"),
  1272 => (x"1e",x"75",x"1e",x"72"),
  1273 => (x"1e",x"d9",x"c3",x"c1"),
  1274 => (x"87",x"f4",x"fd",x"fe"),
  1275 => (x"e8",x"c0",x"86",x"cc"),
  1276 => (x"1e",x"c0",x"c8",x"87"),
  1277 => (x"fc",x"49",x"66",x"dc"),
  1278 => (x"86",x"c4",x"87",x"d3"),
  1279 => (x"6c",x"58",x"a6",x"c4"),
  1280 => (x"c8",x"98",x"73",x"48"),
  1281 => (x"66",x"c4",x"58",x"a6"),
  1282 => (x"6c",x"87",x"cc",x"02"),
  1283 => (x"c8",x"98",x"73",x"48"),
  1284 => (x"66",x"c4",x"58",x"a6"),
  1285 => (x"c0",x"87",x"f4",x"05"),
  1286 => (x"f8",x"48",x"6e",x"7c"),
  1287 => (x"26",x"4d",x"26",x"8e"),
  1288 => (x"26",x"4b",x"26",x"4c"),
  1289 => (x"5b",x"5e",x"0e",x"4f"),
  1290 => (x"fc",x"0e",x"5d",x"5c"),
  1291 => (x"c0",x"1e",x"c0",x"86"),
  1292 => (x"c9",x"c1",x"f0",x"ff"),
  1293 => (x"87",x"e4",x"eb",x"49"),
  1294 => (x"df",x"c1",x"1e",x"d2"),
  1295 => (x"cc",x"fb",x"49",x"f2"),
  1296 => (x"c0",x"86",x"c8",x"87"),
  1297 => (x"d2",x"85",x"c1",x"4d"),
  1298 => (x"f8",x"04",x"ad",x"b7"),
  1299 => (x"f2",x"df",x"c1",x"87"),
  1300 => (x"c3",x"49",x"bf",x"97"),
  1301 => (x"c0",x"c1",x"99",x"c0"),
  1302 => (x"e8",x"c0",x"05",x"a9"),
  1303 => (x"f9",x"df",x"c1",x"87"),
  1304 => (x"d0",x"49",x"bf",x"97"),
  1305 => (x"fa",x"df",x"c1",x"31"),
  1306 => (x"c8",x"4a",x"bf",x"97"),
  1307 => (x"c1",x"b1",x"72",x"32"),
  1308 => (x"bf",x"97",x"fb",x"df"),
  1309 => (x"71",x"b1",x"72",x"4a"),
  1310 => (x"ff",x"ff",x"cf",x"4d"),
  1311 => (x"85",x"c1",x"9d",x"ff"),
  1312 => (x"e6",x"c2",x"35",x"ca"),
  1313 => (x"fb",x"df",x"c1",x"87"),
  1314 => (x"c1",x"4b",x"bf",x"97"),
  1315 => (x"c1",x"9b",x"c6",x"33"),
  1316 => (x"bf",x"97",x"fc",x"df"),
  1317 => (x"29",x"b7",x"c7",x"49"),
  1318 => (x"df",x"c1",x"b3",x"71"),
  1319 => (x"49",x"bf",x"97",x"f7"),
  1320 => (x"98",x"cf",x"48",x"71"),
  1321 => (x"c1",x"58",x"a6",x"c4"),
  1322 => (x"bf",x"97",x"f8",x"df"),
  1323 => (x"ca",x"9c",x"c3",x"4c"),
  1324 => (x"f9",x"df",x"c1",x"34"),
  1325 => (x"c2",x"49",x"bf",x"97"),
  1326 => (x"c1",x"b4",x"71",x"31"),
  1327 => (x"bf",x"97",x"fa",x"df"),
  1328 => (x"99",x"c0",x"c3",x"49"),
  1329 => (x"71",x"29",x"b7",x"c6"),
  1330 => (x"c4",x"1e",x"74",x"b4"),
  1331 => (x"1e",x"73",x"1e",x"66"),
  1332 => (x"1e",x"f9",x"c3",x"c1"),
  1333 => (x"87",x"c8",x"fa",x"fe"),
  1334 => (x"48",x"c1",x"83",x"c2"),
  1335 => (x"4b",x"70",x"30",x"73"),
  1336 => (x"c4",x"c1",x"1e",x"73"),
  1337 => (x"f9",x"fe",x"1e",x"e6"),
  1338 => (x"48",x"c1",x"87",x"f6"),
  1339 => (x"dc",x"30",x"66",x"d8"),
  1340 => (x"a4",x"c1",x"58",x"a6"),
  1341 => (x"95",x"73",x"4d",x"49"),
  1342 => (x"75",x"1e",x"66",x"d8"),
  1343 => (x"ef",x"c4",x"c1",x"1e"),
  1344 => (x"db",x"f9",x"fe",x"1e"),
  1345 => (x"86",x"e4",x"c0",x"87"),
  1346 => (x"c0",x"c8",x"48",x"6e"),
  1347 => (x"ce",x"06",x"a8",x"b7"),
  1348 => (x"c1",x"4b",x"6e",x"87"),
  1349 => (x"c8",x"2b",x"b7",x"35"),
  1350 => (x"01",x"ab",x"b7",x"c0"),
  1351 => (x"75",x"87",x"f4",x"ff"),
  1352 => (x"c5",x"c5",x"c1",x"1e"),
  1353 => (x"f7",x"f8",x"fe",x"1e"),
  1354 => (x"75",x"86",x"c8",x"87"),
  1355 => (x"26",x"8e",x"fc",x"48"),
  1356 => (x"26",x"4c",x"26",x"4d"),
  1357 => (x"1e",x"4f",x"26",x"4b"),
  1358 => (x"4b",x"71",x"1e",x"73"),
  1359 => (x"29",x"d8",x"49",x"73"),
  1360 => (x"73",x"99",x"ff",x"c3"),
  1361 => (x"cf",x"2a",x"c8",x"4a"),
  1362 => (x"72",x"9a",x"c0",x"fc"),
  1363 => (x"c8",x"4a",x"73",x"b1"),
  1364 => (x"f0",x"ff",x"c0",x"32"),
  1365 => (x"72",x"9a",x"c0",x"c0"),
  1366 => (x"d8",x"4a",x"73",x"b1"),
  1367 => (x"c0",x"c0",x"ff",x"32"),
  1368 => (x"72",x"9a",x"c0",x"c0"),
  1369 => (x"26",x"48",x"71",x"b1"),
  1370 => (x"26",x"4f",x"26",x"4b"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
