
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity SoC_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of SoC_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"3b",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"38"),
    10 => (x"20",x"00",x"27",x"4f"),
    11 => (x"27",x"4e",x"00",x"00"),
    12 => (x"00",x"00",x"12",x"29"),
    13 => (x"87",x"fd",x"00",x"0f"),
    14 => (x"4f",x"87",x"fd",x"00"),
    15 => (x"ff",x"86",x"fc",x"1e"),
    16 => (x"48",x"69",x"49",x"c0"),
    17 => (x"c4",x"98",x"c0",x"c4"),
    18 => (x"02",x"6e",x"58",x"a6"),
    19 => (x"66",x"c8",x"87",x"f4"),
    20 => (x"8e",x"fc",x"48",x"79"),
    21 => (x"5e",x"0e",x"4f",x"26"),
    22 => (x"0e",x"5d",x"5c",x"5b"),
    23 => (x"c0",x"4b",x"66",x"d0"),
    24 => (x"71",x"49",x"13",x"4c"),
    25 => (x"87",x"d8",x"02",x"99"),
    26 => (x"c0",x"ff",x"4d",x"71"),
    27 => (x"c4",x"49",x"6a",x"4a"),
    28 => (x"f8",x"02",x"99",x"c0"),
    29 => (x"c1",x"7a",x"75",x"87"),
    30 => (x"71",x"49",x"13",x"84"),
    31 => (x"87",x"e8",x"05",x"99"),
    32 => (x"4d",x"26",x"48",x"74"),
    33 => (x"4b",x"26",x"4c",x"26"),
    34 => (x"5e",x"0e",x"4f",x"26"),
    35 => (x"0e",x"5d",x"5c",x"5b"),
    36 => (x"4b",x"c0",x"86",x"f0"),
    37 => (x"c0",x"48",x"a6",x"c4"),
    38 => (x"a6",x"e4",x"c0",x"78"),
    39 => (x"66",x"e0",x"c0",x"4c"),
    40 => (x"80",x"c1",x"48",x"49"),
    41 => (x"58",x"a6",x"e4",x"c0"),
    42 => (x"c0",x"fe",x"4a",x"11"),
    43 => (x"9a",x"72",x"ba",x"82"),
    44 => (x"87",x"d0",x"c4",x"02"),
    45 => (x"c3",x"02",x"66",x"c4"),
    46 => (x"a6",x"c4",x"87",x"df"),
    47 => (x"72",x"78",x"c0",x"48"),
    48 => (x"aa",x"f0",x"c0",x"49"),
    49 => (x"87",x"ef",x"c2",x"02"),
    50 => (x"02",x"a9",x"e3",x"c1"),
    51 => (x"c1",x"87",x"f0",x"c2"),
    52 => (x"c0",x"02",x"a9",x"e4"),
    53 => (x"ec",x"c1",x"87",x"e1"),
    54 => (x"da",x"c2",x"02",x"a9"),
    55 => (x"a9",x"f0",x"c1",x"87"),
    56 => (x"c1",x"87",x"d4",x"02"),
    57 => (x"c1",x"02",x"a9",x"f3"),
    58 => (x"f5",x"c1",x"87",x"f8"),
    59 => (x"87",x"c7",x"02",x"a9"),
    60 => (x"05",x"a9",x"f8",x"c1"),
    61 => (x"c4",x"87",x"d9",x"c2"),
    62 => (x"c4",x"49",x"74",x"84"),
    63 => (x"6e",x"7e",x"69",x"89"),
    64 => (x"87",x"d1",x"c1",x"02"),
    65 => (x"c0",x"48",x"a6",x"c8"),
    66 => (x"c0",x"80",x"c4",x"78"),
    67 => (x"dc",x"4a",x"6e",x"78"),
    68 => (x"9a",x"cf",x"2a",x"b7"),
    69 => (x"30",x"c4",x"48",x"6e"),
    70 => (x"72",x"58",x"a6",x"c4"),
    71 => (x"87",x"c5",x"02",x"9a"),
    72 => (x"c1",x"48",x"a6",x"c8"),
    73 => (x"06",x"aa",x"c9",x"78"),
    74 => (x"f7",x"c0",x"87",x"c5"),
    75 => (x"c0",x"87",x"c3",x"82"),
    76 => (x"66",x"c8",x"82",x"f0"),
    77 => (x"72",x"87",x"c9",x"02"),
    78 => (x"87",x"c0",x"fc",x"1e"),
    79 => (x"83",x"c1",x"86",x"c4"),
    80 => (x"c1",x"48",x"66",x"cc"),
    81 => (x"58",x"a6",x"d0",x"80"),
    82 => (x"c8",x"48",x"66",x"cc"),
    83 => (x"fe",x"04",x"a8",x"b7"),
    84 => (x"d8",x"c1",x"87",x"fb"),
    85 => (x"1e",x"f0",x"c0",x"87"),
    86 => (x"c4",x"87",x"e1",x"fb"),
    87 => (x"c1",x"83",x"c1",x"86"),
    88 => (x"84",x"c4",x"87",x"cb"),
    89 => (x"89",x"c4",x"49",x"74"),
    90 => (x"e9",x"fb",x"1e",x"69"),
    91 => (x"70",x"86",x"c4",x"87"),
    92 => (x"4b",x"a3",x"71",x"49"),
    93 => (x"c4",x"87",x"f6",x"c0"),
    94 => (x"78",x"c1",x"48",x"a6"),
    95 => (x"c4",x"87",x"ee",x"c0"),
    96 => (x"c4",x"49",x"74",x"84"),
    97 => (x"fa",x"1e",x"69",x"89"),
    98 => (x"86",x"c4",x"87",x"f2"),
    99 => (x"87",x"dd",x"83",x"c1"),
   100 => (x"e7",x"fa",x"1e",x"72"),
   101 => (x"d4",x"86",x"c4",x"87"),
   102 => (x"aa",x"e5",x"c0",x"87"),
   103 => (x"c4",x"87",x"c7",x"05"),
   104 => (x"78",x"c1",x"48",x"a6"),
   105 => (x"1e",x"72",x"87",x"c7"),
   106 => (x"c4",x"87",x"d1",x"fa"),
   107 => (x"66",x"e0",x"c0",x"86"),
   108 => (x"80",x"c1",x"48",x"49"),
   109 => (x"58",x"a6",x"e4",x"c0"),
   110 => (x"c0",x"fe",x"4a",x"11"),
   111 => (x"9a",x"72",x"ba",x"82"),
   112 => (x"87",x"f0",x"fb",x"05"),
   113 => (x"8e",x"f0",x"48",x"73"),
   114 => (x"4c",x"26",x"4d",x"26"),
   115 => (x"4f",x"26",x"4b",x"26"),
   116 => (x"ff",x"86",x"e8",x"1e"),
   117 => (x"ff",x"c3",x"4a",x"d4"),
   118 => (x"c3",x"49",x"6a",x"7a"),
   119 => (x"48",x"6a",x"7a",x"ff"),
   120 => (x"a6",x"c4",x"30",x"c8"),
   121 => (x"59",x"a6",x"c8",x"58"),
   122 => (x"ff",x"c3",x"b1",x"6e"),
   123 => (x"d0",x"48",x"6a",x"7a"),
   124 => (x"58",x"a6",x"cc",x"30"),
   125 => (x"c8",x"59",x"a6",x"d0"),
   126 => (x"ff",x"c3",x"b1",x"66"),
   127 => (x"d8",x"48",x"6a",x"7a"),
   128 => (x"58",x"a6",x"d4",x"30"),
   129 => (x"d0",x"59",x"a6",x"d8"),
   130 => (x"48",x"71",x"b1",x"66"),
   131 => (x"87",x"c6",x"8e",x"e8"),
   132 => (x"4c",x"26",x"4d",x"26"),
   133 => (x"4f",x"26",x"4b",x"26"),
   134 => (x"ff",x"86",x"f4",x"1e"),
   135 => (x"ff",x"c3",x"4a",x"d4"),
   136 => (x"c3",x"49",x"6a",x"7a"),
   137 => (x"48",x"71",x"7a",x"ff"),
   138 => (x"a6",x"c4",x"30",x"c8"),
   139 => (x"6e",x"49",x"6a",x"58"),
   140 => (x"7a",x"ff",x"c3",x"b1"),
   141 => (x"30",x"c8",x"48",x"71"),
   142 => (x"6a",x"58",x"a6",x"c8"),
   143 => (x"b1",x"66",x"c4",x"49"),
   144 => (x"71",x"7a",x"ff",x"c3"),
   145 => (x"cc",x"30",x"c8",x"48"),
   146 => (x"49",x"6a",x"58",x"a6"),
   147 => (x"71",x"b1",x"66",x"c8"),
   148 => (x"ff",x"8e",x"f4",x"48"),
   149 => (x"5e",x"0e",x"87",x"c0"),
   150 => (x"ff",x"0e",x"5c",x"5b"),
   151 => (x"66",x"cc",x"4c",x"d4"),
   152 => (x"98",x"ff",x"c3",x"48"),
   153 => (x"cd",x"c1",x"7c",x"70"),
   154 => (x"c8",x"05",x"bf",x"c4"),
   155 => (x"48",x"66",x"d0",x"87"),
   156 => (x"a6",x"d4",x"30",x"c9"),
   157 => (x"49",x"66",x"d0",x"58"),
   158 => (x"48",x"71",x"29",x"d8"),
   159 => (x"70",x"98",x"ff",x"c3"),
   160 => (x"49",x"66",x"d0",x"7c"),
   161 => (x"48",x"71",x"29",x"d0"),
   162 => (x"70",x"98",x"ff",x"c3"),
   163 => (x"49",x"66",x"d0",x"7c"),
   164 => (x"48",x"71",x"29",x"c8"),
   165 => (x"70",x"98",x"ff",x"c3"),
   166 => (x"48",x"66",x"d0",x"7c"),
   167 => (x"70",x"98",x"ff",x"c3"),
   168 => (x"49",x"66",x"cc",x"7c"),
   169 => (x"48",x"71",x"29",x"d0"),
   170 => (x"70",x"98",x"ff",x"c3"),
   171 => (x"c9",x"4a",x"6c",x"7c"),
   172 => (x"c3",x"4b",x"ff",x"f0"),
   173 => (x"d0",x"05",x"aa",x"ff"),
   174 => (x"7c",x"ff",x"c3",x"87"),
   175 => (x"8b",x"c1",x"4a",x"6c"),
   176 => (x"c3",x"87",x"c6",x"02"),
   177 => (x"f0",x"02",x"aa",x"ff"),
   178 => (x"fd",x"48",x"72",x"87"),
   179 => (x"c0",x"1e",x"87",x"c4"),
   180 => (x"48",x"d4",x"ff",x"49"),
   181 => (x"c1",x"78",x"ff",x"c3"),
   182 => (x"b7",x"c8",x"c3",x"81"),
   183 => (x"87",x"f1",x"04",x"a9"),
   184 => (x"1e",x"87",x"f3",x"fc"),
   185 => (x"87",x"e6",x"1e",x"73"),
   186 => (x"4b",x"df",x"f8",x"c4"),
   187 => (x"ff",x"c0",x"1e",x"c0"),
   188 => (x"1e",x"f7",x"c1",x"f0"),
   189 => (x"c8",x"87",x"df",x"fd"),
   190 => (x"05",x"a8",x"c1",x"86"),
   191 => (x"ff",x"87",x"ea",x"c0"),
   192 => (x"ff",x"c3",x"48",x"d4"),
   193 => (x"c0",x"c0",x"c1",x"78"),
   194 => (x"1e",x"c0",x"c0",x"c0"),
   195 => (x"c1",x"f0",x"e1",x"c0"),
   196 => (x"c1",x"fd",x"1e",x"e9"),
   197 => (x"70",x"86",x"c8",x"87"),
   198 => (x"87",x"ca",x"05",x"98"),
   199 => (x"c3",x"48",x"d4",x"ff"),
   200 => (x"48",x"c1",x"78",x"ff"),
   201 => (x"e5",x"fe",x"87",x"cb"),
   202 => (x"05",x"8b",x"c1",x"87"),
   203 => (x"c0",x"87",x"fd",x"fe"),
   204 => (x"87",x"e0",x"fb",x"48"),
   205 => (x"ff",x"1e",x"73",x"1e"),
   206 => (x"ff",x"c3",x"48",x"d4"),
   207 => (x"1e",x"f1",x"cd",x"78"),
   208 => (x"c4",x"87",x"d3",x"f4"),
   209 => (x"c0",x"4b",x"d3",x"86"),
   210 => (x"f0",x"ff",x"c0",x"1e"),
   211 => (x"fc",x"1e",x"c1",x"c1"),
   212 => (x"86",x"c8",x"87",x"c4"),
   213 => (x"ca",x"05",x"98",x"70"),
   214 => (x"48",x"d4",x"ff",x"87"),
   215 => (x"c1",x"78",x"ff",x"c3"),
   216 => (x"fd",x"87",x"cb",x"48"),
   217 => (x"8b",x"c1",x"87",x"e8"),
   218 => (x"87",x"db",x"ff",x"05"),
   219 => (x"e3",x"fa",x"48",x"c0"),
   220 => (x"44",x"4d",x"43",x"87"),
   221 => (x"5b",x"5e",x"0e",x"00"),
   222 => (x"ff",x"0e",x"5d",x"5c"),
   223 => (x"cd",x"fd",x"4d",x"d4"),
   224 => (x"1e",x"ea",x"c6",x"87"),
   225 => (x"c1",x"f0",x"e1",x"c0"),
   226 => (x"c9",x"fb",x"1e",x"c8"),
   227 => (x"70",x"86",x"c8",x"87"),
   228 => (x"d1",x"1e",x"73",x"4b"),
   229 => (x"f1",x"f3",x"1e",x"fc"),
   230 => (x"c1",x"86",x"c8",x"87"),
   231 => (x"87",x"c8",x"02",x"ab"),
   232 => (x"c0",x"87",x"d1",x"fe"),
   233 => (x"87",x"cf",x"c2",x"48"),
   234 => (x"70",x"87",x"ed",x"f9"),
   235 => (x"ff",x"ff",x"cf",x"49"),
   236 => (x"a9",x"ea",x"c6",x"99"),
   237 => (x"fd",x"87",x"c8",x"02"),
   238 => (x"48",x"c0",x"87",x"fa"),
   239 => (x"c3",x"87",x"f8",x"c1"),
   240 => (x"f1",x"c0",x"7d",x"ff"),
   241 => (x"87",x"db",x"fc",x"4c"),
   242 => (x"c1",x"02",x"98",x"70"),
   243 => (x"1e",x"c0",x"87",x"d0"),
   244 => (x"c1",x"f0",x"ff",x"c0"),
   245 => (x"fd",x"f9",x"1e",x"fa"),
   246 => (x"70",x"86",x"c8",x"87"),
   247 => (x"05",x"9b",x"73",x"4b"),
   248 => (x"73",x"87",x"f1",x"c0"),
   249 => (x"1e",x"fa",x"d0",x"1e"),
   250 => (x"c8",x"87",x"df",x"f2"),
   251 => (x"7d",x"ff",x"c3",x"86"),
   252 => (x"1e",x"73",x"4b",x"6d"),
   253 => (x"f2",x"1e",x"c6",x"d1"),
   254 => (x"86",x"c8",x"87",x"d0"),
   255 => (x"7d",x"7d",x"ff",x"c3"),
   256 => (x"49",x"73",x"7d",x"7d"),
   257 => (x"02",x"99",x"c0",x"c1"),
   258 => (x"48",x"c1",x"87",x"c5"),
   259 => (x"c0",x"87",x"e8",x"c0"),
   260 => (x"87",x"e3",x"c0",x"48"),
   261 => (x"d4",x"d1",x"1e",x"73"),
   262 => (x"87",x"ee",x"f1",x"1e"),
   263 => (x"ac",x"c2",x"86",x"c8"),
   264 => (x"d1",x"87",x"cc",x"05"),
   265 => (x"e1",x"f1",x"1e",x"e0"),
   266 => (x"c0",x"86",x"c4",x"87"),
   267 => (x"c1",x"87",x"c8",x"48"),
   268 => (x"d0",x"fe",x"05",x"8c"),
   269 => (x"f7",x"48",x"c0",x"87"),
   270 => (x"4d",x"43",x"87",x"d6"),
   271 => (x"20",x"38",x"35",x"44"),
   272 => (x"20",x"0a",x"64",x"25"),
   273 => (x"4d",x"43",x"00",x"20"),
   274 => (x"5f",x"38",x"35",x"44"),
   275 => (x"64",x"25",x"20",x"32"),
   276 => (x"00",x"20",x"20",x"0a"),
   277 => (x"35",x"44",x"4d",x"43"),
   278 => (x"64",x"25",x"20",x"38"),
   279 => (x"00",x"20",x"20",x"0a"),
   280 => (x"43",x"48",x"44",x"53"),
   281 => (x"69",x"6e",x"49",x"20"),
   282 => (x"6c",x"61",x"69",x"74"),
   283 => (x"74",x"61",x"7a",x"69"),
   284 => (x"20",x"6e",x"6f",x"69"),
   285 => (x"6f",x"72",x"72",x"65"),
   286 => (x"00",x"0a",x"21",x"72"),
   287 => (x"5f",x"64",x"6d",x"63"),
   288 => (x"38",x"44",x"4d",x"43"),
   289 => (x"73",x"65",x"72",x"20"),
   290 => (x"73",x"6e",x"6f",x"70"),
   291 => (x"25",x"20",x"3a",x"65"),
   292 => (x"0e",x"00",x"0a",x"64"),
   293 => (x"5d",x"5c",x"5b",x"5e"),
   294 => (x"d0",x"ff",x"1e",x"0e"),
   295 => (x"c0",x"c0",x"c8",x"4d"),
   296 => (x"c4",x"cd",x"c1",x"4b"),
   297 => (x"d5",x"78",x"c1",x"48"),
   298 => (x"e9",x"ee",x"1e",x"ef"),
   299 => (x"c7",x"86",x"c4",x"87"),
   300 => (x"73",x"48",x"6d",x"4c"),
   301 => (x"58",x"a6",x"c4",x"98"),
   302 => (x"87",x"cb",x"02",x"6e"),
   303 => (x"98",x"73",x"48",x"6d"),
   304 => (x"6e",x"58",x"a6",x"c4"),
   305 => (x"c0",x"87",x"f5",x"05"),
   306 => (x"87",x"c2",x"f8",x"7d"),
   307 => (x"98",x"73",x"48",x"6d"),
   308 => (x"6e",x"58",x"a6",x"c4"),
   309 => (x"6d",x"87",x"cb",x"02"),
   310 => (x"c4",x"98",x"73",x"48"),
   311 => (x"05",x"6e",x"58",x"a6"),
   312 => (x"7d",x"c1",x"87",x"f5"),
   313 => (x"e5",x"c0",x"1e",x"c0"),
   314 => (x"1e",x"c0",x"c1",x"d0"),
   315 => (x"c8",x"87",x"e7",x"f5"),
   316 => (x"05",x"a8",x"c1",x"86"),
   317 => (x"4c",x"c1",x"87",x"c2"),
   318 => (x"cd",x"05",x"ac",x"c2"),
   319 => (x"1e",x"ea",x"d5",x"87"),
   320 => (x"c4",x"87",x"d3",x"ed"),
   321 => (x"c1",x"48",x"c0",x"86"),
   322 => (x"8c",x"c1",x"87",x"dc"),
   323 => (x"87",x"e1",x"fe",x"05"),
   324 => (x"c1",x"87",x"e2",x"f9"),
   325 => (x"c1",x"58",x"c8",x"cd"),
   326 => (x"05",x"bf",x"c4",x"cd"),
   327 => (x"1e",x"c1",x"87",x"cd"),
   328 => (x"c1",x"f0",x"ff",x"c0"),
   329 => (x"ed",x"f4",x"1e",x"d0"),
   330 => (x"ff",x"86",x"c8",x"87"),
   331 => (x"ff",x"c3",x"48",x"d4"),
   332 => (x"87",x"c8",x"c6",x"78"),
   333 => (x"58",x"cc",x"cd",x"c1"),
   334 => (x"bf",x"c8",x"cd",x"c1"),
   335 => (x"1e",x"f3",x"d5",x"1e"),
   336 => (x"c8",x"87",x"c7",x"ed"),
   337 => (x"73",x"48",x"6d",x"86"),
   338 => (x"58",x"a6",x"c4",x"98"),
   339 => (x"87",x"cc",x"02",x"6e"),
   340 => (x"98",x"73",x"48",x"6d"),
   341 => (x"6e",x"58",x"a6",x"c4"),
   342 => (x"87",x"f4",x"ff",x"05"),
   343 => (x"d4",x"ff",x"7d",x"c0"),
   344 => (x"78",x"ff",x"c3",x"48"),
   345 => (x"f2",x"26",x"48",x"c1"),
   346 => (x"45",x"49",x"87",x"e6"),
   347 => (x"53",x"00",x"52",x"52"),
   348 => (x"53",x"00",x"49",x"50"),
   349 => (x"61",x"63",x"20",x"44"),
   350 => (x"73",x"20",x"64",x"72"),
   351 => (x"20",x"65",x"7a",x"69"),
   352 => (x"25",x"20",x"73",x"69"),
   353 => (x"0e",x"00",x"0a",x"64"),
   354 => (x"0e",x"5c",x"5b",x"5e"),
   355 => (x"cc",x"4c",x"66",x"d0"),
   356 => (x"4a",x"c0",x"4b",x"66"),
   357 => (x"df",x"cd",x"ee",x"c5"),
   358 => (x"48",x"d4",x"ff",x"49"),
   359 => (x"70",x"78",x"ff",x"c3"),
   360 => (x"fe",x"c3",x"48",x"bf"),
   361 => (x"d3",x"c1",x"05",x"a8"),
   362 => (x"c0",x"cd",x"c1",x"87"),
   363 => (x"c4",x"78",x"c0",x"48"),
   364 => (x"db",x"04",x"ac",x"b7"),
   365 => (x"87",x"d8",x"f0",x"87"),
   366 => (x"7b",x"71",x"49",x"70"),
   367 => (x"cd",x"c1",x"83",x"c4"),
   368 => (x"71",x"48",x"bf",x"c0"),
   369 => (x"c4",x"cd",x"c1",x"80"),
   370 => (x"b7",x"8c",x"c4",x"58"),
   371 => (x"87",x"e5",x"03",x"ac"),
   372 => (x"06",x"ac",x"b7",x"c0"),
   373 => (x"ff",x"87",x"e2",x"c0"),
   374 => (x"ff",x"c3",x"48",x"d4"),
   375 => (x"49",x"bf",x"70",x"78"),
   376 => (x"c1",x"7b",x"97",x"71"),
   377 => (x"c0",x"cd",x"c1",x"83"),
   378 => (x"80",x"71",x"48",x"bf"),
   379 => (x"58",x"c4",x"cd",x"c1"),
   380 => (x"b7",x"c0",x"8c",x"c1"),
   381 => (x"de",x"ff",x"01",x"ac"),
   382 => (x"4a",x"49",x"c1",x"87"),
   383 => (x"fe",x"05",x"89",x"c1"),
   384 => (x"d4",x"ff",x"87",x"d7"),
   385 => (x"78",x"ff",x"c3",x"48"),
   386 => (x"c5",x"f0",x"48",x"72"),
   387 => (x"5b",x"5e",x"0e",x"87"),
   388 => (x"c8",x"1e",x"0e",x"5c"),
   389 => (x"c0",x"4c",x"c0",x"c0"),
   390 => (x"48",x"d4",x"ff",x"4b"),
   391 => (x"ff",x"78",x"ff",x"c3"),
   392 => (x"74",x"48",x"bf",x"d0"),
   393 => (x"58",x"a6",x"c4",x"98"),
   394 => (x"87",x"cd",x"02",x"6e"),
   395 => (x"48",x"bf",x"d0",x"ff"),
   396 => (x"a6",x"c4",x"98",x"74"),
   397 => (x"f3",x"05",x"6e",x"58"),
   398 => (x"48",x"d0",x"ff",x"87"),
   399 => (x"ff",x"78",x"c1",x"c4"),
   400 => (x"ff",x"c3",x"48",x"d4"),
   401 => (x"1e",x"66",x"d0",x"78"),
   402 => (x"c1",x"f0",x"ff",x"c0"),
   403 => (x"c5",x"f0",x"1e",x"d1"),
   404 => (x"70",x"86",x"c8",x"87"),
   405 => (x"02",x"99",x"71",x"49"),
   406 => (x"1e",x"71",x"87",x"d0"),
   407 => (x"da",x"1e",x"66",x"d4"),
   408 => (x"e5",x"e8",x"1e",x"dc"),
   409 => (x"c0",x"86",x"cc",x"87"),
   410 => (x"c0",x"c8",x"87",x"ec"),
   411 => (x"1e",x"66",x"d8",x"1e"),
   412 => (x"c8",x"87",x"d4",x"fc"),
   413 => (x"ff",x"4b",x"70",x"86"),
   414 => (x"74",x"48",x"bf",x"d0"),
   415 => (x"58",x"a6",x"c4",x"98"),
   416 => (x"87",x"cd",x"02",x"6e"),
   417 => (x"48",x"bf",x"d0",x"ff"),
   418 => (x"a6",x"c4",x"98",x"74"),
   419 => (x"f3",x"05",x"6e",x"58"),
   420 => (x"48",x"d0",x"ff",x"87"),
   421 => (x"48",x"73",x"78",x"c0"),
   422 => (x"87",x"f6",x"ed",x"26"),
   423 => (x"64",x"61",x"65",x"52"),
   424 => (x"6d",x"6f",x"63",x"20"),
   425 => (x"64",x"6e",x"61",x"6d"),
   426 => (x"69",x"61",x"66",x"20"),
   427 => (x"20",x"64",x"65",x"6c"),
   428 => (x"25",x"20",x"74",x"61"),
   429 => (x"25",x"28",x"20",x"64"),
   430 => (x"00",x"0a",x"29",x"64"),
   431 => (x"5c",x"5b",x"5e",x"0e"),
   432 => (x"c0",x"1e",x"0e",x"5d"),
   433 => (x"f0",x"ff",x"c0",x"1e"),
   434 => (x"ee",x"1e",x"c9",x"c1"),
   435 => (x"86",x"c8",x"87",x"c8"),
   436 => (x"cd",x"c1",x"1e",x"d2"),
   437 => (x"ee",x"fa",x"1e",x"d2"),
   438 => (x"c0",x"86",x"c8",x"87"),
   439 => (x"d2",x"85",x"c1",x"4d"),
   440 => (x"f8",x"04",x"ad",x"b7"),
   441 => (x"d2",x"cd",x"c1",x"87"),
   442 => (x"c3",x"49",x"bf",x"97"),
   443 => (x"c0",x"c1",x"99",x"c0"),
   444 => (x"e8",x"c0",x"05",x"a9"),
   445 => (x"d9",x"cd",x"c1",x"87"),
   446 => (x"d0",x"49",x"bf",x"97"),
   447 => (x"da",x"cd",x"c1",x"31"),
   448 => (x"c8",x"4a",x"bf",x"97"),
   449 => (x"c1",x"b1",x"72",x"32"),
   450 => (x"bf",x"97",x"db",x"cd"),
   451 => (x"71",x"b1",x"72",x"4a"),
   452 => (x"ff",x"ff",x"cf",x"4d"),
   453 => (x"85",x"c1",x"9d",x"ff"),
   454 => (x"e6",x"c2",x"35",x"ca"),
   455 => (x"db",x"cd",x"c1",x"87"),
   456 => (x"c1",x"4b",x"bf",x"97"),
   457 => (x"c1",x"9b",x"c6",x"33"),
   458 => (x"bf",x"97",x"dc",x"cd"),
   459 => (x"29",x"b7",x"c7",x"49"),
   460 => (x"cd",x"c1",x"b3",x"71"),
   461 => (x"49",x"bf",x"97",x"d7"),
   462 => (x"98",x"cf",x"48",x"71"),
   463 => (x"c1",x"58",x"a6",x"c4"),
   464 => (x"bf",x"97",x"d8",x"cd"),
   465 => (x"ca",x"9c",x"c3",x"4c"),
   466 => (x"d9",x"cd",x"c1",x"34"),
   467 => (x"c2",x"49",x"bf",x"97"),
   468 => (x"c1",x"b4",x"71",x"31"),
   469 => (x"bf",x"97",x"da",x"cd"),
   470 => (x"99",x"c0",x"c3",x"49"),
   471 => (x"71",x"29",x"b7",x"c6"),
   472 => (x"c4",x"1e",x"74",x"b4"),
   473 => (x"1e",x"73",x"1e",x"66"),
   474 => (x"e4",x"1e",x"c9",x"df"),
   475 => (x"86",x"d0",x"87",x"dc"),
   476 => (x"48",x"c1",x"83",x"c2"),
   477 => (x"4b",x"70",x"30",x"73"),
   478 => (x"f6",x"df",x"1e",x"73"),
   479 => (x"87",x"ca",x"e4",x"1e"),
   480 => (x"48",x"c1",x"86",x"c8"),
   481 => (x"a6",x"c4",x"30",x"6e"),
   482 => (x"49",x"a4",x"c1",x"58"),
   483 => (x"6e",x"95",x"73",x"4d"),
   484 => (x"df",x"1e",x"75",x"1e"),
   485 => (x"f1",x"e3",x"1e",x"ff"),
   486 => (x"6e",x"86",x"cc",x"87"),
   487 => (x"b7",x"c0",x"c8",x"48"),
   488 => (x"87",x"d4",x"06",x"a8"),
   489 => (x"48",x"6e",x"35",x"c1"),
   490 => (x"c4",x"28",x"b7",x"c1"),
   491 => (x"48",x"6e",x"58",x"a6"),
   492 => (x"a8",x"b7",x"c0",x"c8"),
   493 => (x"87",x"ec",x"ff",x"01"),
   494 => (x"e0",x"c0",x"1e",x"75"),
   495 => (x"c9",x"e3",x"1e",x"d5"),
   496 => (x"75",x"86",x"c8",x"87"),
   497 => (x"c7",x"e9",x"26",x"48"),
   498 => (x"73",x"5f",x"63",x"87"),
   499 => (x"5f",x"65",x"7a",x"69"),
   500 => (x"74",x"6c",x"75",x"6d"),
   501 => (x"64",x"25",x"20",x"3a"),
   502 => (x"65",x"72",x"20",x"2c"),
   503 => (x"62",x"5f",x"64",x"61"),
   504 => (x"65",x"6c",x"5f",x"6c"),
   505 => (x"25",x"20",x"3a",x"6e"),
   506 => (x"63",x"20",x"2c",x"64"),
   507 => (x"65",x"7a",x"69",x"73"),
   508 => (x"64",x"25",x"20",x"3a"),
   509 => (x"75",x"4d",x"00",x"0a"),
   510 => (x"25",x"20",x"74",x"6c"),
   511 => (x"25",x"00",x"0a",x"64"),
   512 => (x"6c",x"62",x"20",x"64"),
   513 => (x"73",x"6b",x"63",x"6f"),
   514 => (x"20",x"66",x"6f",x"20"),
   515 => (x"65",x"7a",x"69",x"73"),
   516 => (x"0a",x"64",x"25",x"20"),
   517 => (x"20",x"64",x"25",x"00"),
   518 => (x"63",x"6f",x"6c",x"62"),
   519 => (x"6f",x"20",x"73",x"6b"),
   520 => (x"31",x"35",x"20",x"66"),
   521 => (x"79",x"62",x"20",x"32"),
   522 => (x"0a",x"73",x"65",x"74"),
   523 => (x"1e",x"73",x"1e",x"00"),
   524 => (x"66",x"d0",x"4b",x"c0"),
   525 => (x"a8",x"b7",x"c0",x"48"),
   526 => (x"87",x"f6",x"c0",x"06"),
   527 => (x"bf",x"97",x"66",x"c8"),
   528 => (x"82",x"c0",x"fe",x"4a"),
   529 => (x"48",x"66",x"c8",x"ba"),
   530 => (x"a6",x"cc",x"80",x"c1"),
   531 => (x"97",x"66",x"cc",x"58"),
   532 => (x"c0",x"fe",x"49",x"bf"),
   533 => (x"66",x"cc",x"b9",x"81"),
   534 => (x"d0",x"80",x"c1",x"48"),
   535 => (x"b7",x"71",x"58",x"a6"),
   536 => (x"87",x"c4",x"02",x"aa"),
   537 => (x"87",x"cc",x"48",x"c1"),
   538 => (x"66",x"d0",x"83",x"c1"),
   539 => (x"ff",x"04",x"ab",x"b7"),
   540 => (x"48",x"c0",x"87",x"ca"),
   541 => (x"4d",x"26",x"87",x"c4"),
   542 => (x"4b",x"26",x"4c",x"26"),
   543 => (x"5e",x"0e",x"4f",x"26"),
   544 => (x"0e",x"5d",x"5c",x"5b"),
   545 => (x"48",x"ec",x"d5",x"c1"),
   546 => (x"f1",x"c0",x"78",x"c0"),
   547 => (x"df",x"ff",x"1e",x"e2"),
   548 => (x"86",x"c4",x"87",x"c4"),
   549 => (x"1e",x"e4",x"cd",x"c1"),
   550 => (x"f0",x"f5",x"1e",x"c0"),
   551 => (x"70",x"86",x"c8",x"87"),
   552 => (x"87",x"cf",x"05",x"98"),
   553 => (x"1e",x"ce",x"ee",x"c0"),
   554 => (x"87",x"ea",x"de",x"ff"),
   555 => (x"48",x"c0",x"86",x"c4"),
   556 => (x"c0",x"87",x"d8",x"cb"),
   557 => (x"ff",x"1e",x"ef",x"f1"),
   558 => (x"c4",x"87",x"db",x"de"),
   559 => (x"c1",x"4b",x"c0",x"86"),
   560 => (x"c1",x"48",x"d8",x"d6"),
   561 => (x"c0",x"1e",x"c8",x"78"),
   562 => (x"c1",x"1e",x"c6",x"f2"),
   563 => (x"fd",x"1e",x"da",x"ce"),
   564 => (x"86",x"cc",x"87",x"db"),
   565 => (x"c6",x"05",x"98",x"70"),
   566 => (x"d8",x"d6",x"c1",x"87"),
   567 => (x"c8",x"78",x"c0",x"48"),
   568 => (x"cf",x"f2",x"c0",x"1e"),
   569 => (x"f6",x"ce",x"c1",x"1e"),
   570 => (x"87",x"c1",x"fd",x"1e"),
   571 => (x"98",x"70",x"86",x"cc"),
   572 => (x"c1",x"87",x"c6",x"05"),
   573 => (x"c0",x"48",x"d8",x"d6"),
   574 => (x"d8",x"d6",x"c1",x"78"),
   575 => (x"f2",x"c0",x"1e",x"bf"),
   576 => (x"de",x"ff",x"1e",x"d8"),
   577 => (x"86",x"c8",x"87",x"c4"),
   578 => (x"bf",x"d8",x"d6",x"c1"),
   579 => (x"87",x"d5",x"c2",x"02"),
   580 => (x"4d",x"e4",x"cd",x"c1"),
   581 => (x"4c",x"e2",x"d4",x"c1"),
   582 => (x"9f",x"e2",x"d5",x"c1"),
   583 => (x"1e",x"71",x"49",x"bf"),
   584 => (x"49",x"e2",x"d5",x"c1"),
   585 => (x"89",x"e4",x"cd",x"c1"),
   586 => (x"1e",x"d0",x"1e",x"71"),
   587 => (x"c0",x"1e",x"c0",x"c8"),
   588 => (x"ff",x"1e",x"c0",x"ef"),
   589 => (x"d4",x"87",x"d3",x"dd"),
   590 => (x"49",x"a4",x"c8",x"86"),
   591 => (x"d5",x"c1",x"4b",x"69"),
   592 => (x"49",x"bf",x"9f",x"e2"),
   593 => (x"a9",x"ea",x"d6",x"c5"),
   594 => (x"87",x"cf",x"c0",x"05"),
   595 => (x"69",x"49",x"a4",x"c8"),
   596 => (x"87",x"fe",x"d8",x"1e"),
   597 => (x"4b",x"70",x"86",x"c4"),
   598 => (x"c7",x"87",x"de",x"c0"),
   599 => (x"9f",x"49",x"a5",x"fe"),
   600 => (x"e9",x"ca",x"49",x"69"),
   601 => (x"c0",x"02",x"a9",x"d5"),
   602 => (x"ee",x"c0",x"87",x"cf"),
   603 => (x"db",x"ff",x"1e",x"e2"),
   604 => (x"86",x"c4",x"87",x"e4"),
   605 => (x"d2",x"c8",x"48",x"c0"),
   606 => (x"c0",x"1e",x"73",x"87"),
   607 => (x"ff",x"1e",x"fd",x"ef"),
   608 => (x"c8",x"87",x"c7",x"dc"),
   609 => (x"e4",x"cd",x"c1",x"86"),
   610 => (x"f1",x"1e",x"73",x"1e"),
   611 => (x"86",x"c8",x"87",x"ff"),
   612 => (x"c0",x"05",x"98",x"70"),
   613 => (x"48",x"c0",x"87",x"c5"),
   614 => (x"c0",x"87",x"f0",x"c7"),
   615 => (x"ff",x"1e",x"d5",x"f0"),
   616 => (x"c4",x"87",x"f3",x"da"),
   617 => (x"eb",x"f2",x"c0",x"86"),
   618 => (x"dd",x"db",x"ff",x"1e"),
   619 => (x"c8",x"86",x"c4",x"87"),
   620 => (x"c3",x"f3",x"c0",x"1e"),
   621 => (x"f6",x"ce",x"c1",x"1e"),
   622 => (x"87",x"f1",x"f9",x"1e"),
   623 => (x"98",x"70",x"86",x"cc"),
   624 => (x"87",x"c9",x"c0",x"05"),
   625 => (x"48",x"ec",x"d5",x"c1"),
   626 => (x"e4",x"c0",x"78",x"c1"),
   627 => (x"c0",x"1e",x"c8",x"87"),
   628 => (x"c1",x"1e",x"cc",x"f3"),
   629 => (x"f9",x"1e",x"da",x"ce"),
   630 => (x"86",x"cc",x"87",x"d3"),
   631 => (x"c0",x"02",x"98",x"70"),
   632 => (x"f0",x"c0",x"87",x"cf"),
   633 => (x"da",x"ff",x"1e",x"fc"),
   634 => (x"86",x"c4",x"87",x"e0"),
   635 => (x"da",x"c6",x"48",x"c0"),
   636 => (x"e2",x"d5",x"c1",x"87"),
   637 => (x"c1",x"49",x"bf",x"97"),
   638 => (x"c0",x"05",x"a9",x"d5"),
   639 => (x"d5",x"c1",x"87",x"cd"),
   640 => (x"49",x"bf",x"97",x"e3"),
   641 => (x"02",x"a9",x"ea",x"c2"),
   642 => (x"c0",x"87",x"c5",x"c0"),
   643 => (x"87",x"fb",x"c5",x"48"),
   644 => (x"97",x"e4",x"cd",x"c1"),
   645 => (x"e9",x"c3",x"49",x"bf"),
   646 => (x"d2",x"c0",x"02",x"a9"),
   647 => (x"e4",x"cd",x"c1",x"87"),
   648 => (x"c3",x"49",x"bf",x"97"),
   649 => (x"c0",x"02",x"a9",x"eb"),
   650 => (x"48",x"c0",x"87",x"c5"),
   651 => (x"c1",x"87",x"dc",x"c5"),
   652 => (x"bf",x"97",x"ef",x"cd"),
   653 => (x"05",x"99",x"71",x"49"),
   654 => (x"c1",x"87",x"cc",x"c0"),
   655 => (x"bf",x"97",x"f0",x"cd"),
   656 => (x"02",x"a9",x"c2",x"49"),
   657 => (x"c0",x"87",x"c5",x"c0"),
   658 => (x"87",x"ff",x"c4",x"48"),
   659 => (x"97",x"f1",x"cd",x"c1"),
   660 => (x"d5",x"c1",x"48",x"bf"),
   661 => (x"d5",x"c1",x"58",x"e8"),
   662 => (x"71",x"49",x"bf",x"e4"),
   663 => (x"c1",x"8a",x"c1",x"4a"),
   664 => (x"72",x"5a",x"ec",x"d5"),
   665 => (x"c0",x"1e",x"71",x"1e"),
   666 => (x"ff",x"1e",x"d5",x"f3"),
   667 => (x"cc",x"87",x"db",x"d8"),
   668 => (x"f2",x"cd",x"c1",x"86"),
   669 => (x"73",x"49",x"bf",x"97"),
   670 => (x"f3",x"cd",x"c1",x"81"),
   671 => (x"c8",x"4a",x"bf",x"97"),
   672 => (x"f8",x"d5",x"c1",x"32"),
   673 => (x"78",x"a1",x"72",x"48"),
   674 => (x"97",x"f4",x"cd",x"c1"),
   675 => (x"d6",x"c1",x"48",x"bf"),
   676 => (x"d5",x"c1",x"58",x"d0"),
   677 => (x"c2",x"02",x"bf",x"ec"),
   678 => (x"1e",x"c8",x"87",x"df"),
   679 => (x"1e",x"d9",x"f1",x"c0"),
   680 => (x"1e",x"f6",x"ce",x"c1"),
   681 => (x"cc",x"87",x"c6",x"f6"),
   682 => (x"02",x"98",x"70",x"86"),
   683 => (x"c0",x"87",x"c5",x"c0"),
   684 => (x"87",x"d7",x"c3",x"48"),
   685 => (x"bf",x"e4",x"d5",x"c1"),
   686 => (x"c4",x"48",x"72",x"4a"),
   687 => (x"d4",x"d6",x"c1",x"30"),
   688 => (x"cc",x"d6",x"c1",x"58"),
   689 => (x"c9",x"ce",x"c1",x"5a"),
   690 => (x"c8",x"49",x"bf",x"97"),
   691 => (x"c8",x"ce",x"c1",x"31"),
   692 => (x"73",x"4b",x"bf",x"97"),
   693 => (x"ce",x"c1",x"49",x"a1"),
   694 => (x"4b",x"bf",x"97",x"ca"),
   695 => (x"a1",x"73",x"33",x"d0"),
   696 => (x"cb",x"ce",x"c1",x"49"),
   697 => (x"d8",x"4b",x"bf",x"97"),
   698 => (x"49",x"a1",x"73",x"33"),
   699 => (x"59",x"d8",x"d6",x"c1"),
   700 => (x"bf",x"cc",x"d6",x"c1"),
   701 => (x"f8",x"d5",x"c1",x"91"),
   702 => (x"d6",x"c1",x"81",x"bf"),
   703 => (x"ce",x"c1",x"59",x"c0"),
   704 => (x"4b",x"bf",x"97",x"d1"),
   705 => (x"ce",x"c1",x"33",x"c8"),
   706 => (x"4c",x"bf",x"97",x"d0"),
   707 => (x"c1",x"4b",x"a3",x"74"),
   708 => (x"bf",x"97",x"d2",x"ce"),
   709 => (x"74",x"34",x"d0",x"4c"),
   710 => (x"ce",x"c1",x"4b",x"a3"),
   711 => (x"4c",x"bf",x"97",x"d3"),
   712 => (x"34",x"d8",x"9c",x"cf"),
   713 => (x"c1",x"4b",x"a3",x"74"),
   714 => (x"c2",x"5b",x"c4",x"d6"),
   715 => (x"c1",x"92",x"73",x"8b"),
   716 => (x"72",x"48",x"c4",x"d6"),
   717 => (x"d0",x"c1",x"78",x"a1"),
   718 => (x"f6",x"cd",x"c1",x"87"),
   719 => (x"c8",x"49",x"bf",x"97"),
   720 => (x"f5",x"cd",x"c1",x"31"),
   721 => (x"72",x"4a",x"bf",x"97"),
   722 => (x"d6",x"c1",x"49",x"a1"),
   723 => (x"31",x"c5",x"59",x"d4"),
   724 => (x"c9",x"81",x"ff",x"c7"),
   725 => (x"cc",x"d6",x"c1",x"29"),
   726 => (x"fb",x"cd",x"c1",x"59"),
   727 => (x"c8",x"4a",x"bf",x"97"),
   728 => (x"fa",x"cd",x"c1",x"32"),
   729 => (x"73",x"4b",x"bf",x"97"),
   730 => (x"d6",x"c1",x"4a",x"a2"),
   731 => (x"d6",x"c1",x"5a",x"d8"),
   732 => (x"c1",x"92",x"bf",x"cc"),
   733 => (x"82",x"bf",x"f8",x"d5"),
   734 => (x"5a",x"c8",x"d6",x"c1"),
   735 => (x"48",x"c0",x"d6",x"c1"),
   736 => (x"d5",x"c1",x"78",x"c0"),
   737 => (x"a1",x"72",x"48",x"fc"),
   738 => (x"f3",x"48",x"c1",x"78"),
   739 => (x"65",x"52",x"87",x"e8"),
   740 => (x"6f",x"20",x"64",x"61"),
   741 => (x"42",x"4d",x"20",x"66"),
   742 => (x"61",x"66",x"20",x"52"),
   743 => (x"64",x"65",x"6c",x"69"),
   744 => (x"6f",x"4e",x"00",x"0a"),
   745 => (x"72",x"61",x"70",x"20"),
   746 => (x"69",x"74",x"69",x"74"),
   747 => (x"73",x"20",x"6e",x"6f"),
   748 => (x"61",x"6e",x"67",x"69"),
   749 => (x"65",x"72",x"75",x"74"),
   750 => (x"75",x"6f",x"66",x"20"),
   751 => (x"00",x"0a",x"64",x"6e"),
   752 => (x"73",x"52",x"42",x"4d"),
   753 => (x"3a",x"65",x"7a",x"69"),
   754 => (x"2c",x"64",x"25",x"20"),
   755 => (x"72",x"61",x"70",x"20"),
   756 => (x"69",x"74",x"69",x"74"),
   757 => (x"69",x"73",x"6e",x"6f"),
   758 => (x"20",x"3a",x"65",x"7a"),
   759 => (x"20",x"2c",x"64",x"25"),
   760 => (x"73",x"66",x"66",x"6f"),
   761 => (x"6f",x"20",x"74",x"65"),
   762 => (x"69",x"73",x"20",x"66"),
   763 => (x"25",x"20",x"3a",x"67"),
   764 => (x"73",x"20",x"2c",x"64"),
   765 => (x"30",x"20",x"67",x"69"),
   766 => (x"0a",x"78",x"25",x"78"),
   767 => (x"61",x"65",x"52",x"00"),
   768 => (x"67",x"6e",x"69",x"64"),
   769 => (x"6f",x"6f",x"62",x"20"),
   770 => (x"65",x"73",x"20",x"74"),
   771 => (x"72",x"6f",x"74",x"63"),
   772 => (x"0a",x"64",x"25",x"20"),
   773 => (x"61",x"65",x"52",x"00"),
   774 => (x"6f",x"62",x"20",x"64"),
   775 => (x"73",x"20",x"74",x"6f"),
   776 => (x"6f",x"74",x"63",x"65"),
   777 => (x"72",x"66",x"20",x"72"),
   778 => (x"66",x"20",x"6d",x"6f"),
   779 => (x"74",x"73",x"72",x"69"),
   780 => (x"72",x"61",x"70",x"20"),
   781 => (x"69",x"74",x"69",x"74"),
   782 => (x"00",x"0a",x"6e",x"6f"),
   783 => (x"75",x"73",x"6e",x"55"),
   784 => (x"72",x"6f",x"70",x"70"),
   785 => (x"20",x"64",x"65",x"74"),
   786 => (x"74",x"72",x"61",x"70"),
   787 => (x"6f",x"69",x"74",x"69"),
   788 => (x"79",x"74",x"20",x"6e"),
   789 => (x"0d",x"21",x"65",x"70"),
   790 => (x"54",x"41",x"46",x"00"),
   791 => (x"20",x"20",x"32",x"33"),
   792 => (x"65",x"52",x"00",x"20"),
   793 => (x"6e",x"69",x"64",x"61"),
   794 => (x"42",x"4d",x"20",x"67"),
   795 => (x"4d",x"00",x"0a",x"52"),
   796 => (x"73",x"20",x"52",x"42"),
   797 => (x"65",x"63",x"63",x"75"),
   798 => (x"75",x"66",x"73",x"73"),
   799 => (x"20",x"79",x"6c",x"6c"),
   800 => (x"64",x"61",x"65",x"72"),
   801 => (x"41",x"46",x"00",x"0a"),
   802 => (x"20",x"36",x"31",x"54"),
   803 => (x"46",x"00",x"20",x"20"),
   804 => (x"32",x"33",x"54",x"41"),
   805 => (x"00",x"20",x"20",x"20"),
   806 => (x"74",x"72",x"61",x"50"),
   807 => (x"6f",x"69",x"74",x"69"),
   808 => (x"75",x"6f",x"63",x"6e"),
   809 => (x"25",x"20",x"74",x"6e"),
   810 => (x"48",x"00",x"0a",x"64"),
   811 => (x"69",x"74",x"6e",x"75"),
   812 => (x"66",x"20",x"67",x"6e"),
   813 => (x"66",x"20",x"72",x"6f"),
   814 => (x"73",x"65",x"6c",x"69"),
   815 => (x"65",x"74",x"73",x"79"),
   816 => (x"46",x"00",x"0a",x"6d"),
   817 => (x"32",x"33",x"54",x"41"),
   818 => (x"00",x"20",x"20",x"20"),
   819 => (x"31",x"54",x"41",x"46"),
   820 => (x"20",x"20",x"20",x"36"),
   821 => (x"75",x"6c",x"43",x"00"),
   822 => (x"72",x"65",x"74",x"73"),
   823 => (x"7a",x"69",x"73",x"20"),
   824 => (x"25",x"20",x"3a",x"65"),
   825 => (x"43",x"20",x"2c",x"64"),
   826 => (x"74",x"73",x"75",x"6c"),
   827 => (x"6d",x"20",x"72",x"65"),
   828 => (x"2c",x"6b",x"73",x"61"),
   829 => (x"0a",x"64",x"25",x"20"),
   830 => (x"5b",x"5e",x"0e",x"00"),
   831 => (x"d5",x"c1",x"0e",x"5c"),
   832 => (x"ce",x"02",x"bf",x"ec"),
   833 => (x"4a",x"66",x"cc",x"87"),
   834 => (x"cc",x"2a",x"b7",x"c7"),
   835 => (x"ff",x"c1",x"4b",x"66"),
   836 => (x"cc",x"87",x"cc",x"9b"),
   837 => (x"b7",x"c8",x"4a",x"66"),
   838 => (x"4b",x"66",x"cc",x"2a"),
   839 => (x"c1",x"9b",x"ff",x"c3"),
   840 => (x"c1",x"1e",x"e4",x"cd"),
   841 => (x"49",x"bf",x"f8",x"d5"),
   842 => (x"1e",x"71",x"81",x"72"),
   843 => (x"c8",x"87",x"de",x"e3"),
   844 => (x"05",x"98",x"70",x"86"),
   845 => (x"48",x"c0",x"87",x"c5"),
   846 => (x"c1",x"87",x"e6",x"c0"),
   847 => (x"02",x"bf",x"ec",x"d5"),
   848 => (x"49",x"73",x"87",x"d2"),
   849 => (x"cd",x"c1",x"91",x"c4"),
   850 => (x"4c",x"69",x"81",x"e4"),
   851 => (x"ff",x"ff",x"ff",x"cf"),
   852 => (x"87",x"cb",x"9c",x"ff"),
   853 => (x"91",x"c2",x"49",x"73"),
   854 => (x"81",x"e4",x"cd",x"c1"),
   855 => (x"74",x"4c",x"69",x"9f"),
   856 => (x"87",x"d4",x"ec",x"48"),
   857 => (x"5c",x"5b",x"5e",x"0e"),
   858 => (x"86",x"f4",x"0e",x"5d"),
   859 => (x"d6",x"c1",x"4b",x"c0"),
   860 => (x"c4",x"7e",x"bf",x"c0"),
   861 => (x"d6",x"c1",x"48",x"a6"),
   862 => (x"c1",x"78",x"bf",x"c4"),
   863 => (x"02",x"bf",x"ec",x"d5"),
   864 => (x"d5",x"c1",x"87",x"c9"),
   865 => (x"c4",x"49",x"bf",x"e4"),
   866 => (x"c1",x"87",x"c7",x"31"),
   867 => (x"49",x"bf",x"c8",x"d6"),
   868 => (x"a6",x"cc",x"31",x"c4"),
   869 => (x"c8",x"4d",x"c0",x"59"),
   870 => (x"a8",x"c0",x"48",x"66"),
   871 => (x"87",x"e9",x"c2",x"06"),
   872 => (x"99",x"cf",x"49",x"75"),
   873 => (x"c1",x"87",x"da",x"05"),
   874 => (x"c8",x"1e",x"e4",x"cd"),
   875 => (x"c1",x"48",x"49",x"66"),
   876 => (x"58",x"a6",x"cc",x"80"),
   877 => (x"d4",x"e1",x"1e",x"71"),
   878 => (x"c1",x"86",x"c8",x"87"),
   879 => (x"c3",x"4b",x"e4",x"cd"),
   880 => (x"83",x"e0",x"c0",x"87"),
   881 => (x"71",x"49",x"6b",x"97"),
   882 => (x"f3",x"c1",x"02",x"99"),
   883 => (x"49",x"6b",x"97",x"87"),
   884 => (x"02",x"a9",x"e5",x"c3"),
   885 => (x"cb",x"87",x"e9",x"c1"),
   886 => (x"69",x"97",x"49",x"a3"),
   887 => (x"05",x"99",x"d8",x"49"),
   888 => (x"73",x"87",x"dd",x"c1"),
   889 => (x"ed",x"c9",x"ff",x"1e"),
   890 => (x"cb",x"86",x"c4",x"87"),
   891 => (x"66",x"e4",x"c0",x"1e"),
   892 => (x"e8",x"1e",x"73",x"1e"),
   893 => (x"86",x"cc",x"87",x"f7"),
   894 => (x"c1",x"05",x"98",x"70"),
   895 => (x"a3",x"dc",x"87",x"c2"),
   896 => (x"49",x"66",x"dc",x"4a"),
   897 => (x"79",x"6a",x"81",x"c4"),
   898 => (x"dc",x"4a",x"a3",x"da"),
   899 => (x"81",x"c8",x"49",x"66"),
   900 => (x"70",x"48",x"6a",x"9f"),
   901 => (x"c1",x"4c",x"71",x"79"),
   902 => (x"02",x"bf",x"ec",x"d5"),
   903 => (x"a3",x"d4",x"87",x"d0"),
   904 => (x"49",x"69",x"9f",x"49"),
   905 => (x"ff",x"c0",x"4a",x"71"),
   906 => (x"32",x"d0",x"9a",x"ff"),
   907 => (x"4a",x"c0",x"87",x"c2"),
   908 => (x"80",x"6c",x"48",x"72"),
   909 => (x"66",x"dc",x"7c",x"70"),
   910 => (x"c1",x"78",x"c0",x"48"),
   911 => (x"87",x"ff",x"c0",x"48"),
   912 => (x"66",x"c8",x"85",x"c1"),
   913 => (x"d7",x"fd",x"04",x"ad"),
   914 => (x"ec",x"d5",x"c1",x"87"),
   915 => (x"ec",x"c0",x"02",x"bf"),
   916 => (x"fa",x"1e",x"6e",x"87"),
   917 => (x"86",x"c4",x"87",x"e3"),
   918 => (x"6e",x"58",x"a6",x"c4"),
   919 => (x"ff",x"ff",x"cf",x"49"),
   920 => (x"a9",x"99",x"f8",x"ff"),
   921 => (x"6e",x"87",x"d6",x"02"),
   922 => (x"c1",x"89",x"c2",x"49"),
   923 => (x"91",x"bf",x"e4",x"d5"),
   924 => (x"bf",x"fc",x"d5",x"c1"),
   925 => (x"c8",x"80",x"71",x"48"),
   926 => (x"d8",x"fc",x"58",x"a6"),
   927 => (x"f4",x"48",x"c0",x"87"),
   928 => (x"87",x"f2",x"e7",x"8e"),
   929 => (x"c8",x"1e",x"73",x"1e"),
   930 => (x"c1",x"49",x"bf",x"66"),
   931 => (x"09",x"66",x"c8",x"81"),
   932 => (x"d5",x"c1",x"09",x"79"),
   933 => (x"05",x"99",x"bf",x"e8"),
   934 => (x"66",x"c8",x"87",x"d0"),
   935 => (x"6b",x"83",x"c8",x"4b"),
   936 => (x"87",x"d5",x"f9",x"1e"),
   937 => (x"49",x"70",x"86",x"c4"),
   938 => (x"48",x"c1",x"7b",x"71"),
   939 => (x"1e",x"87",x"cb",x"e7"),
   940 => (x"bf",x"fc",x"d5",x"c1"),
   941 => (x"4a",x"66",x"c4",x"49"),
   942 => (x"4a",x"6a",x"82",x"c8"),
   943 => (x"d5",x"c1",x"8a",x"c2"),
   944 => (x"72",x"92",x"bf",x"e4"),
   945 => (x"d5",x"c1",x"49",x"a1"),
   946 => (x"c4",x"4a",x"bf",x"e8"),
   947 => (x"72",x"9a",x"bf",x"66"),
   948 => (x"66",x"c8",x"49",x"a1"),
   949 => (x"ff",x"1e",x"71",x"1e"),
   950 => (x"c8",x"87",x"f2",x"dc"),
   951 => (x"05",x"98",x"70",x"86"),
   952 => (x"48",x"c0",x"87",x"c4"),
   953 => (x"48",x"c1",x"87",x"c2"),
   954 => (x"0e",x"87",x"d1",x"e6"),
   955 => (x"0e",x"5c",x"5b",x"5e"),
   956 => (x"c1",x"1e",x"66",x"cc"),
   957 => (x"f9",x"1e",x"dc",x"d6"),
   958 => (x"86",x"c8",x"87",x"ea"),
   959 => (x"c1",x"02",x"98",x"70"),
   960 => (x"d6",x"c1",x"87",x"d2"),
   961 => (x"c7",x"49",x"bf",x"e0"),
   962 => (x"29",x"c9",x"81",x"ff"),
   963 => (x"4b",x"c0",x"4c",x"71"),
   964 => (x"1e",x"ea",x"fd",x"c0"),
   965 => (x"87",x"fe",x"c4",x"ff"),
   966 => (x"b7",x"c0",x"86",x"c4"),
   967 => (x"c4",x"c1",x"06",x"ac"),
   968 => (x"1e",x"66",x"d0",x"87"),
   969 => (x"1e",x"dc",x"d6",x"c1"),
   970 => (x"c8",x"87",x"c4",x"fe"),
   971 => (x"05",x"98",x"70",x"86"),
   972 => (x"48",x"c0",x"87",x"c5"),
   973 => (x"c1",x"87",x"f0",x"c0"),
   974 => (x"fd",x"1e",x"dc",x"d6"),
   975 => (x"86",x"c4",x"87",x"c6"),
   976 => (x"c8",x"48",x"66",x"d0"),
   977 => (x"a6",x"d4",x"80",x"c0"),
   978 => (x"74",x"83",x"c1",x"58"),
   979 => (x"ff",x"04",x"ab",x"b7"),
   980 => (x"87",x"d1",x"87",x"cf"),
   981 => (x"c0",x"1e",x"66",x"cc"),
   982 => (x"ff",x"1e",x"c3",x"fe"),
   983 => (x"c8",x"87",x"eb",x"c4"),
   984 => (x"c2",x"48",x"c0",x"86"),
   985 => (x"e4",x"48",x"c1",x"87"),
   986 => (x"70",x"4f",x"87",x"ce"),
   987 => (x"64",x"65",x"6e",x"65"),
   988 => (x"6c",x"69",x"66",x"20"),
   989 => (x"6c",x"20",x"2c",x"65"),
   990 => (x"69",x"64",x"61",x"6f"),
   991 => (x"2e",x"2e",x"67",x"6e"),
   992 => (x"43",x"00",x"0a",x"2e"),
   993 => (x"74",x"27",x"6e",x"61"),
   994 => (x"65",x"70",x"6f",x"20"),
   995 => (x"73",x"25",x"20",x"6e"),
   996 => (x"c4",x"1e",x"00",x"0a"),
   997 => (x"29",x"d8",x"49",x"66"),
   998 => (x"c4",x"99",x"ff",x"c3"),
   999 => (x"2a",x"c8",x"4a",x"66"),
  1000 => (x"9a",x"c0",x"fc",x"cf"),
  1001 => (x"66",x"c4",x"b1",x"72"),
  1002 => (x"c0",x"32",x"c8",x"4a"),
  1003 => (x"c0",x"c0",x"f0",x"ff"),
  1004 => (x"c4",x"b1",x"72",x"9a"),
  1005 => (x"32",x"d8",x"4a",x"66"),
  1006 => (x"c0",x"c0",x"c0",x"ff"),
  1007 => (x"b1",x"72",x"9a",x"c0"),
  1008 => (x"87",x"c6",x"48",x"71"),
  1009 => (x"4c",x"26",x"4d",x"26"),
  1010 => (x"4f",x"26",x"4b",x"26"),
  1011 => (x"d0",x"1e",x"73",x"1e"),
  1012 => (x"c0",x"c0",x"c0",x"c0"),
  1013 => (x"fe",x"0f",x"73",x"4b"),
  1014 => (x"26",x"87",x"c4",x"87"),
  1015 => (x"26",x"4c",x"26",x"4d"),
  1016 => (x"1e",x"4f",x"26",x"4b"),
  1017 => (x"c3",x"49",x"66",x"c8"),
  1018 => (x"f7",x"c0",x"99",x"df"),
  1019 => (x"a9",x"b7",x"c0",x"89"),
  1020 => (x"c0",x"87",x"c3",x"03"),
  1021 => (x"66",x"c4",x"81",x"e7"),
  1022 => (x"c8",x"30",x"c4",x"48"),
  1023 => (x"66",x"c4",x"58",x"a6"),
  1024 => (x"c8",x"b0",x"71",x"48"),
  1025 => (x"66",x"c4",x"58",x"a6"),
  1026 => (x"87",x"d5",x"ff",x"48"),
  1027 => (x"5c",x"5b",x"5e",x"0e"),
  1028 => (x"c0",x"c0",x"d0",x"0e"),
  1029 => (x"c1",x"4c",x"c0",x"c0"),
  1030 => (x"48",x"bf",x"e8",x"d6"),
  1031 => (x"d6",x"c1",x"80",x"c1"),
  1032 => (x"cc",x"97",x"58",x"ec"),
  1033 => (x"c0",x"fe",x"49",x"66"),
  1034 => (x"d3",x"c1",x"b9",x"81"),
  1035 => (x"87",x"db",x"05",x"a9"),
  1036 => (x"48",x"e8",x"d6",x"c1"),
  1037 => (x"d6",x"c1",x"78",x"c0"),
  1038 => (x"78",x"c0",x"48",x"ec"),
  1039 => (x"48",x"f4",x"d6",x"c1"),
  1040 => (x"d6",x"c1",x"78",x"c0"),
  1041 => (x"78",x"c0",x"48",x"f8"),
  1042 => (x"c1",x"87",x"f8",x"c6"),
  1043 => (x"48",x"bf",x"e8",x"d6"),
  1044 => (x"c0",x"05",x"a8",x"c1"),
  1045 => (x"cc",x"97",x"87",x"f8"),
  1046 => (x"c0",x"fe",x"49",x"66"),
  1047 => (x"1e",x"71",x"b9",x"81"),
  1048 => (x"bf",x"f8",x"d6",x"c1"),
  1049 => (x"87",x"fb",x"fd",x"1e"),
  1050 => (x"d6",x"c1",x"86",x"c8"),
  1051 => (x"d6",x"c1",x"58",x"fc"),
  1052 => (x"c3",x"4a",x"bf",x"f8"),
  1053 => (x"c6",x"06",x"aa",x"b7"),
  1054 => (x"72",x"48",x"ca",x"87"),
  1055 => (x"72",x"4a",x"70",x"88"),
  1056 => (x"71",x"81",x"c1",x"49"),
  1057 => (x"c1",x"30",x"c1",x"48"),
  1058 => (x"c5",x"58",x"f4",x"d6"),
  1059 => (x"d6",x"c1",x"87",x"f5"),
  1060 => (x"c9",x"48",x"bf",x"f8"),
  1061 => (x"c5",x"01",x"a8",x"b7"),
  1062 => (x"d6",x"c1",x"87",x"e9"),
  1063 => (x"c0",x"48",x"bf",x"f8"),
  1064 => (x"c5",x"06",x"a8",x"b7"),
  1065 => (x"d6",x"c1",x"87",x"dd"),
  1066 => (x"c3",x"48",x"bf",x"e8"),
  1067 => (x"db",x"01",x"a8",x"b7"),
  1068 => (x"66",x"cc",x"97",x"87"),
  1069 => (x"81",x"c0",x"fe",x"49"),
  1070 => (x"c1",x"1e",x"71",x"b9"),
  1071 => (x"1e",x"bf",x"f4",x"d6"),
  1072 => (x"c8",x"87",x"e0",x"fc"),
  1073 => (x"f8",x"d6",x"c1",x"86"),
  1074 => (x"87",x"f7",x"c4",x"58"),
  1075 => (x"bf",x"f0",x"d6",x"c1"),
  1076 => (x"c1",x"81",x"c3",x"49"),
  1077 => (x"b7",x"bf",x"e8",x"d6"),
  1078 => (x"e1",x"c0",x"04",x"a9"),
  1079 => (x"66",x"cc",x"97",x"87"),
  1080 => (x"81",x"c0",x"fe",x"49"),
  1081 => (x"c1",x"1e",x"71",x"b9"),
  1082 => (x"1e",x"bf",x"ec",x"d6"),
  1083 => (x"c8",x"87",x"f4",x"fb"),
  1084 => (x"f0",x"d6",x"c1",x"86"),
  1085 => (x"fc",x"d6",x"c1",x"58"),
  1086 => (x"c4",x"78",x"c1",x"48"),
  1087 => (x"d6",x"c1",x"87",x"c5"),
  1088 => (x"c0",x"48",x"bf",x"f8"),
  1089 => (x"c2",x"06",x"a8",x"b7"),
  1090 => (x"d6",x"c1",x"87",x"d8"),
  1091 => (x"c3",x"48",x"bf",x"f8"),
  1092 => (x"c2",x"01",x"a8",x"b7"),
  1093 => (x"d6",x"c1",x"87",x"cc"),
  1094 => (x"c1",x"49",x"bf",x"f4"),
  1095 => (x"d6",x"c1",x"81",x"31"),
  1096 => (x"a9",x"b7",x"bf",x"e8"),
  1097 => (x"87",x"dc",x"c1",x"04"),
  1098 => (x"49",x"66",x"cc",x"97"),
  1099 => (x"b9",x"81",x"c0",x"fe"),
  1100 => (x"d7",x"c1",x"1e",x"71"),
  1101 => (x"fa",x"1e",x"bf",x"c0"),
  1102 => (x"86",x"c8",x"87",x"e9"),
  1103 => (x"58",x"c4",x"d7",x"c1"),
  1104 => (x"bf",x"fc",x"d6",x"c1"),
  1105 => (x"c1",x"89",x"c1",x"49"),
  1106 => (x"c0",x"59",x"c0",x"d7"),
  1107 => (x"c2",x"03",x"a9",x"b7"),
  1108 => (x"d6",x"c1",x"87",x"f1"),
  1109 => (x"c1",x"49",x"bf",x"ec"),
  1110 => (x"bf",x"97",x"c0",x"d7"),
  1111 => (x"ec",x"d6",x"c1",x"51"),
  1112 => (x"81",x"c1",x"49",x"bf"),
  1113 => (x"59",x"f0",x"d6",x"c1"),
  1114 => (x"bf",x"c4",x"d7",x"c1"),
  1115 => (x"c0",x"06",x"a9",x"b7"),
  1116 => (x"d7",x"c1",x"87",x"c9"),
  1117 => (x"d6",x"c1",x"48",x"c4"),
  1118 => (x"c1",x"78",x"bf",x"ec"),
  1119 => (x"c1",x"48",x"fc",x"d6"),
  1120 => (x"87",x"ff",x"c1",x"78"),
  1121 => (x"bf",x"fc",x"d6",x"c1"),
  1122 => (x"87",x"f7",x"c1",x"05"),
  1123 => (x"bf",x"c0",x"d7",x"c1"),
  1124 => (x"c1",x"31",x"c4",x"49"),
  1125 => (x"c1",x"59",x"c4",x"d7"),
  1126 => (x"09",x"bf",x"ec",x"d6"),
  1127 => (x"c1",x"09",x"79",x"97"),
  1128 => (x"d6",x"c1",x"87",x"e1"),
  1129 => (x"c7",x"48",x"bf",x"f8"),
  1130 => (x"c1",x"04",x"a8",x"b7"),
  1131 => (x"4b",x"c0",x"87",x"d5"),
  1132 => (x"c1",x"48",x"f4",x"fe"),
  1133 => (x"c4",x"d7",x"c1",x"78"),
  1134 => (x"1e",x"74",x"1e",x"bf"),
  1135 => (x"1e",x"c6",x"c8",x"c1"),
  1136 => (x"87",x"c6",x"fb",x"fe"),
  1137 => (x"d6",x"c1",x"86",x"cc"),
  1138 => (x"d6",x"c1",x"5c",x"f0"),
  1139 => (x"c1",x"48",x"bf",x"ec"),
  1140 => (x"b7",x"bf",x"c4",x"d7"),
  1141 => (x"db",x"c0",x"03",x"a8"),
  1142 => (x"ec",x"d6",x"c1",x"87"),
  1143 => (x"c1",x"83",x"bf",x"bf"),
  1144 => (x"49",x"bf",x"ec",x"d6"),
  1145 => (x"d6",x"c1",x"81",x"c4"),
  1146 => (x"d7",x"c1",x"59",x"f0"),
  1147 => (x"a9",x"b7",x"bf",x"c4"),
  1148 => (x"87",x"e5",x"ff",x"04"),
  1149 => (x"c8",x"c1",x"1e",x"73"),
  1150 => (x"fa",x"fe",x"1e",x"e5"),
  1151 => (x"86",x"c8",x"87",x"cc"),
  1152 => (x"f7",x"87",x"c9",x"f7"),
  1153 => (x"68",x"43",x"87",x"d7"),
  1154 => (x"73",x"6b",x"63",x"65"),
  1155 => (x"69",x"6d",x"6d",x"75"),
  1156 => (x"66",x"20",x"67",x"6e"),
  1157 => (x"20",x"6d",x"6f",x"72"),
  1158 => (x"74",x"20",x"64",x"25"),
  1159 => (x"64",x"25",x"20",x"6f"),
  1160 => (x"20",x"2e",x"2e",x"2e"),
  1161 => (x"0a",x"64",x"25",x"00"),
  1162 => (x"5b",x"5e",x"0e",x"00"),
  1163 => (x"c1",x"0e",x"5d",x"5c"),
  1164 => (x"fe",x"1e",x"c0",x"cc"),
  1165 => (x"c4",x"87",x"df",x"f8"),
  1166 => (x"d6",x"c9",x"ff",x"86"),
  1167 => (x"02",x"98",x"70",x"87"),
  1168 => (x"d8",x"ff",x"87",x"cd"),
  1169 => (x"98",x"70",x"87",x"f8"),
  1170 => (x"c1",x"87",x"c4",x"02"),
  1171 => (x"c0",x"87",x"c2",x"49"),
  1172 => (x"c1",x"4d",x"71",x"49"),
  1173 => (x"fe",x"1e",x"d6",x"cc"),
  1174 => (x"c4",x"87",x"fb",x"f7"),
  1175 => (x"c4",x"d7",x"c1",x"86"),
  1176 => (x"c0",x"78",x"c0",x"48"),
  1177 => (x"f7",x"fe",x"1e",x"ee"),
  1178 => (x"86",x"c4",x"87",x"d2"),
  1179 => (x"ff",x"c8",x"f4",x"c3"),
  1180 => (x"bf",x"c0",x"ff",x"4a"),
  1181 => (x"c8",x"49",x"74",x"4c"),
  1182 => (x"c1",x"02",x"99",x"c0"),
  1183 => (x"4b",x"74",x"87",x"ca"),
  1184 => (x"db",x"9b",x"ff",x"c3"),
  1185 => (x"f3",x"c0",x"05",x"ab"),
  1186 => (x"02",x"9d",x"75",x"87"),
  1187 => (x"d0",x"87",x"e3",x"c0"),
  1188 => (x"c0",x"c0",x"c0",x"c0"),
  1189 => (x"e4",x"cb",x"c1",x"1e"),
  1190 => (x"87",x"cf",x"f1",x"1e"),
  1191 => (x"98",x"70",x"86",x"c8"),
  1192 => (x"c1",x"87",x"cf",x"02"),
  1193 => (x"fe",x"1e",x"d8",x"cb"),
  1194 => (x"c4",x"87",x"eb",x"f6"),
  1195 => (x"87",x"dc",x"f4",x"86"),
  1196 => (x"cb",x"c1",x"87",x"ca"),
  1197 => (x"f6",x"fe",x"1e",x"f0"),
  1198 => (x"86",x"c4",x"87",x"dc"),
  1199 => (x"cb",x"f5",x"1e",x"73"),
  1200 => (x"c3",x"86",x"c4",x"87"),
  1201 => (x"4a",x"c0",x"c9",x"f4"),
  1202 => (x"8a",x"c1",x"49",x"72"),
  1203 => (x"fe",x"05",x"99",x"71"),
  1204 => (x"ce",x"fe",x"87",x"df"),
  1205 => (x"87",x"c3",x"f4",x"87"),
  1206 => (x"74",x"6f",x"6f",x"42"),
  1207 => (x"2e",x"67",x"6e",x"69"),
  1208 => (x"00",x"0a",x"2e",x"2e"),
  1209 => (x"54",x"4f",x"4f",x"42"),
  1210 => (x"20",x"32",x"33",x"38"),
  1211 => (x"00",x"4e",x"49",x"42"),
  1212 => (x"62",x"20",x"44",x"53"),
  1213 => (x"20",x"74",x"6f",x"6f"),
  1214 => (x"6c",x"69",x"61",x"66"),
  1215 => (x"00",x"0a",x"64",x"65"),
  1216 => (x"74",x"69",x"6e",x"49"),
  1217 => (x"69",x"6c",x"61",x"69"),
  1218 => (x"67",x"6e",x"69",x"7a"),
  1219 => (x"20",x"44",x"53",x"20"),
  1220 => (x"64",x"72",x"61",x"63"),
  1221 => (x"53",x"52",x"00",x"0a"),
  1222 => (x"20",x"32",x"33",x"32"),
  1223 => (x"74",x"6f",x"6f",x"62"),
  1224 => (x"70",x"20",x"2d",x"20"),
  1225 => (x"73",x"73",x"65",x"72"),
  1226 => (x"43",x"53",x"45",x"20"),
  1227 => (x"20",x"6f",x"74",x"20"),
  1228 => (x"74",x"6f",x"6f",x"62"),
  1229 => (x"6f",x"72",x"66",x"20"),
  1230 => (x"44",x"53",x"20",x"6d"),
  1231 => (x"44",x"53",x"00",x"2e"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
