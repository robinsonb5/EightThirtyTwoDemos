
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Dhrystone_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Dhrystone_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**(maxAddrBitBRAM)-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to (2 ** (maxAddrBitBRAM-1)) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"d7",x"01"),
     1 => (x"58",x"0e",x"87",x"da"),
     2 => (x"27",x"0e",x"59",x"5e"),
     3 => (x"00",x"00",x"00",x"41"),
     4 => (x"26",x"49",x"26",x"0f"),
     5 => (x"26",x"80",x"ff",x"48"),
     6 => (x"26",x"27",x"4f",x"08"),
     7 => (x"4f",x"00",x"00",x"00"),
     8 => (x"00",x"00",x"33",x"27"),
     9 => (x"c0",x"c2",x"4f",x"00"),
    10 => (x"f7",x"27",x"4e",x"c0"),
    11 => (x"0f",x"00",x"00",x"06"),
    12 => (x"c1",x"87",x"fd",x"00"),
    13 => (x"27",x"4e",x"c0",x"f0"),
    14 => (x"00",x"00",x"00",x"40"),
    15 => (x"87",x"fd",x"00",x"0f"),
    16 => (x"72",x"1e",x"4f",x"4f"),
    17 => (x"c0",x"ff",x"1e",x"1e"),
    18 => (x"c4",x"48",x"6a",x"4a"),
    19 => (x"a6",x"c4",x"98",x"c0"),
    20 => (x"ff",x"02",x"6e",x"58"),
    21 => (x"66",x"cc",x"87",x"f3"),
    22 => (x"48",x"66",x"cc",x"7a"),
    23 => (x"26",x"4a",x"26",x"26"),
    24 => (x"5a",x"5e",x"0e",x"4f"),
    25 => (x"0e",x"5d",x"5c",x"5b"),
    26 => (x"c0",x"4b",x"66",x"d4"),
    27 => (x"74",x"4c",x"13",x"4d"),
    28 => (x"d9",x"c0",x"02",x"9c"),
    29 => (x"c3",x"4a",x"74",x"87"),
    30 => (x"1e",x"72",x"9a",x"ff"),
    31 => (x"00",x"00",x"42",x"27"),
    32 => (x"86",x"c4",x"0f",x"00"),
    33 => (x"4c",x"13",x"85",x"c1"),
    34 => (x"ff",x"05",x"9c",x"74"),
    35 => (x"48",x"75",x"87",x"e7"),
    36 => (x"4c",x"26",x"4d",x"26"),
    37 => (x"4a",x"26",x"4b",x"26"),
    38 => (x"5e",x"0e",x"4f",x"26"),
    39 => (x"5d",x"5c",x"5b",x"5a"),
    40 => (x"66",x"d8",x"1e",x"0e"),
    41 => (x"18",x"08",x"27",x"4c"),
    42 => (x"76",x"4b",x"00",x"00"),
    43 => (x"10",x"4c",x"27",x"49"),
    44 => (x"c0",x"79",x"00",x"00"),
    45 => (x"05",x"9c",x"74",x"4d"),
    46 => (x"c0",x"87",x"c6",x"c0"),
    47 => (x"f4",x"c0",x"53",x"f0"),
    48 => (x"02",x"9c",x"74",x"87"),
    49 => (x"74",x"87",x"ee",x"c0"),
    50 => (x"c0",x"1e",x"72",x"49"),
    51 => (x"27",x"4a",x"66",x"e0"),
    52 => (x"00",x"00",x"06",x"7b"),
    53 => (x"71",x"4a",x"26",x"0f"),
    54 => (x"12",x"82",x"6e",x"4a"),
    55 => (x"72",x"49",x"74",x"53"),
    56 => (x"66",x"e0",x"c0",x"1e"),
    57 => (x"06",x"7b",x"27",x"4a"),
    58 => (x"26",x"0f",x"00",x"00"),
    59 => (x"74",x"4c",x"70",x"4a"),
    60 => (x"d2",x"ff",x"05",x"9c"),
    61 => (x"18",x"08",x"27",x"87"),
    62 => (x"02",x"ab",x"00",x"00"),
    63 => (x"c0",x"87",x"ea",x"c0"),
    64 => (x"c0",x"4c",x"66",x"e0"),
    65 => (x"c1",x"1e",x"66",x"e4"),
    66 => (x"4a",x"6b",x"97",x"8b"),
    67 => (x"c0",x"c0",x"c0",x"c1"),
    68 => (x"c0",x"c4",x"92",x"c0"),
    69 => (x"72",x"4a",x"92",x"b7"),
    70 => (x"c8",x"0f",x"74",x"1e"),
    71 => (x"27",x"85",x"c1",x"86"),
    72 => (x"00",x"00",x"18",x"08"),
    73 => (x"da",x"ff",x"05",x"ab"),
    74 => (x"26",x"48",x"75",x"87"),
    75 => (x"4c",x"26",x"4d",x"26"),
    76 => (x"4a",x"26",x"4b",x"26"),
    77 => (x"5e",x"0e",x"4f",x"26"),
    78 => (x"5d",x"5c",x"5b",x"5a"),
    79 => (x"4c",x"66",x"d4",x"0e"),
    80 => (x"4b",x"14",x"4d",x"ff"),
    81 => (x"c0",x"c0",x"c0",x"c1"),
    82 => (x"c0",x"c4",x"93",x"c0"),
    83 => (x"73",x"4b",x"93",x"b7"),
    84 => (x"e8",x"c0",x"02",x"9b"),
    85 => (x"dc",x"85",x"c1",x"87"),
    86 => (x"1e",x"73",x"1e",x"66"),
    87 => (x"0f",x"66",x"e0",x"c0"),
    88 => (x"4a",x"70",x"86",x"c8"),
    89 => (x"c0",x"05",x"aa",x"73"),
    90 => (x"4b",x"14",x"87",x"d3"),
    91 => (x"c0",x"c0",x"c0",x"c1"),
    92 => (x"c0",x"c4",x"93",x"c0"),
    93 => (x"73",x"4b",x"93",x"b7"),
    94 => (x"d8",x"ff",x"05",x"9b"),
    95 => (x"26",x"48",x"75",x"87"),
    96 => (x"26",x"4c",x"26",x"4d"),
    97 => (x"26",x"4a",x"26",x"4b"),
    98 => (x"5a",x"5e",x"0e",x"4f"),
    99 => (x"0e",x"5d",x"5c",x"5b"),
   100 => (x"e8",x"c0",x"8e",x"cc"),
   101 => (x"4c",x"c0",x"4b",x"66"),
   102 => (x"c0",x"49",x"a6",x"c4"),
   103 => (x"66",x"e0",x"c0",x"79"),
   104 => (x"c1",x"4d",x"bf",x"97"),
   105 => (x"c0",x"c0",x"c0",x"c0"),
   106 => (x"b7",x"c0",x"c4",x"95"),
   107 => (x"e0",x"c0",x"4d",x"95"),
   108 => (x"80",x"c1",x"48",x"66"),
   109 => (x"58",x"a6",x"e4",x"c0"),
   110 => (x"c5",x"02",x"9d",x"75"),
   111 => (x"66",x"c4",x"87",x"ce"),
   112 => (x"87",x"ce",x"c4",x"02"),
   113 => (x"c0",x"49",x"a6",x"c8"),
   114 => (x"49",x"a6",x"c4",x"79"),
   115 => (x"4a",x"75",x"79",x"c0"),
   116 => (x"02",x"ad",x"f0",x"c0"),
   117 => (x"c1",x"87",x"e8",x"c1"),
   118 => (x"c1",x"02",x"aa",x"e3"),
   119 => (x"e4",x"c1",x"87",x"e9"),
   120 => (x"e6",x"c0",x"02",x"aa"),
   121 => (x"aa",x"ec",x"c1",x"87"),
   122 => (x"87",x"d3",x"c1",x"02"),
   123 => (x"02",x"aa",x"f0",x"c1"),
   124 => (x"c1",x"87",x"e0",x"c0"),
   125 => (x"c0",x"02",x"aa",x"f3"),
   126 => (x"f5",x"c1",x"87",x"e1"),
   127 => (x"ca",x"c0",x"02",x"aa"),
   128 => (x"aa",x"f8",x"c1",x"87"),
   129 => (x"87",x"cb",x"c0",x"02"),
   130 => (x"c8",x"87",x"db",x"c1"),
   131 => (x"79",x"ca",x"49",x"a6"),
   132 => (x"c8",x"87",x"ea",x"c1"),
   133 => (x"79",x"d0",x"49",x"a6"),
   134 => (x"c0",x"87",x"e2",x"c1"),
   135 => (x"73",x"1e",x"66",x"ec"),
   136 => (x"66",x"ec",x"c0",x"1e"),
   137 => (x"c0",x"80",x"c4",x"48"),
   138 => (x"c0",x"58",x"a6",x"f0"),
   139 => (x"c4",x"4a",x"66",x"ec"),
   140 => (x"fc",x"1e",x"6a",x"8a"),
   141 => (x"86",x"cc",x"87",x"c0"),
   142 => (x"84",x"72",x"4a",x"70"),
   143 => (x"c4",x"87",x"fe",x"c0"),
   144 => (x"79",x"c1",x"49",x"a6"),
   145 => (x"c0",x"87",x"f6",x"c0"),
   146 => (x"c0",x"1e",x"66",x"ec"),
   147 => (x"c4",x"48",x"66",x"e8"),
   148 => (x"a6",x"ec",x"c0",x"80"),
   149 => (x"66",x"e8",x"c0",x"58"),
   150 => (x"6a",x"8a",x"c4",x"4a"),
   151 => (x"c8",x"0f",x"73",x"1e"),
   152 => (x"c0",x"84",x"c1",x"86"),
   153 => (x"ec",x"c0",x"87",x"d7"),
   154 => (x"e5",x"c0",x"1e",x"66"),
   155 => (x"c8",x"0f",x"73",x"1e"),
   156 => (x"66",x"ec",x"c0",x"86"),
   157 => (x"73",x"1e",x"75",x"1e"),
   158 => (x"c1",x"86",x"c8",x"0f"),
   159 => (x"02",x"66",x"c8",x"84"),
   160 => (x"c0",x"87",x"e8",x"c1"),
   161 => (x"c4",x"48",x"66",x"e4"),
   162 => (x"a6",x"e8",x"c0",x"80"),
   163 => (x"66",x"e4",x"c0",x"58"),
   164 => (x"76",x"8a",x"c4",x"4a"),
   165 => (x"c1",x"79",x"6a",x"49"),
   166 => (x"c0",x"05",x"ad",x"e4"),
   167 => (x"49",x"6e",x"87",x"dc"),
   168 => (x"03",x"a9",x"b7",x"c0"),
   169 => (x"c0",x"87",x"d3",x"c0"),
   170 => (x"42",x"27",x"1e",x"ed"),
   171 => (x"0f",x"00",x"00",x"00"),
   172 => (x"48",x"6e",x"86",x"c4"),
   173 => (x"c4",x"88",x"08",x"c0"),
   174 => (x"ec",x"c0",x"58",x"a6"),
   175 => (x"1e",x"73",x"1e",x"66"),
   176 => (x"cc",x"1e",x"66",x"d0"),
   177 => (x"d1",x"f7",x"1e",x"66"),
   178 => (x"70",x"86",x"d0",x"87"),
   179 => (x"c0",x"84",x"72",x"4a"),
   180 => (x"e5",x"c0",x"87",x"d9"),
   181 => (x"c8",x"c0",x"05",x"ad"),
   182 => (x"49",x"a6",x"c4",x"87"),
   183 => (x"ca",x"c0",x"79",x"c1"),
   184 => (x"66",x"ec",x"c0",x"87"),
   185 => (x"73",x"1e",x"75",x"1e"),
   186 => (x"c0",x"86",x"c8",x"0f"),
   187 => (x"bf",x"97",x"66",x"e0"),
   188 => (x"c0",x"c0",x"c1",x"4d"),
   189 => (x"c4",x"95",x"c0",x"c0"),
   190 => (x"4d",x"95",x"b7",x"c0"),
   191 => (x"48",x"66",x"e0",x"c0"),
   192 => (x"e4",x"c0",x"80",x"c1"),
   193 => (x"9d",x"75",x"58",x"a6"),
   194 => (x"87",x"f2",x"fa",x"05"),
   195 => (x"86",x"cc",x"48",x"74"),
   196 => (x"4c",x"26",x"4d",x"26"),
   197 => (x"4a",x"26",x"4b",x"26"),
   198 => (x"72",x"1e",x"4f",x"26"),
   199 => (x"27",x"1e",x"c0",x"1e"),
   200 => (x"00",x"00",x"00",x"42"),
   201 => (x"1e",x"66",x"d4",x"1e"),
   202 => (x"27",x"1e",x"66",x"d4"),
   203 => (x"00",x"00",x"01",x"89"),
   204 => (x"70",x"86",x"d0",x"0f"),
   205 => (x"26",x"48",x"72",x"4a"),
   206 => (x"1e",x"4f",x"26",x"4a"),
   207 => (x"a6",x"cc",x"1e",x"72"),
   208 => (x"27",x"1e",x"c0",x"4a"),
   209 => (x"00",x"00",x"00",x"42"),
   210 => (x"d4",x"1e",x"72",x"1e"),
   211 => (x"89",x"27",x"1e",x"66"),
   212 => (x"0f",x"00",x"00",x"01"),
   213 => (x"4a",x"70",x"86",x"d0"),
   214 => (x"4a",x"26",x"48",x"72"),
   215 => (x"5e",x"0e",x"4f",x"26"),
   216 => (x"d0",x"0e",x"5b",x"5a"),
   217 => (x"66",x"d0",x"4b",x"66"),
   218 => (x"6a",x"82",x"c4",x"4a"),
   219 => (x"87",x"dc",x"c0",x"02"),
   220 => (x"82",x"c4",x"4a",x"73"),
   221 => (x"88",x"c1",x"48",x"6a"),
   222 => (x"4a",x"6b",x"7a",x"70"),
   223 => (x"80",x"c1",x"48",x"72"),
   224 => (x"cc",x"97",x"7b",x"70"),
   225 => (x"66",x"cc",x"52",x"66"),
   226 => (x"87",x"c2",x"c0",x"48"),
   227 => (x"4b",x"26",x"48",x"c0"),
   228 => (x"4f",x"26",x"4a",x"26"),
   229 => (x"5b",x"5a",x"5e",x"0e"),
   230 => (x"76",x"8e",x"c8",x"0e"),
   231 => (x"79",x"66",x"d4",x"49"),
   232 => (x"ff",x"49",x"a6",x"c4"),
   233 => (x"4a",x"a6",x"dc",x"79"),
   234 => (x"1e",x"73",x"4b",x"76"),
   235 => (x"00",x"03",x"5e",x"27"),
   236 => (x"1e",x"72",x"1e",x"00"),
   237 => (x"1e",x"66",x"e4",x"c0"),
   238 => (x"00",x"01",x"89",x"27"),
   239 => (x"86",x"d0",x"0f",x"00"),
   240 => (x"48",x"72",x"4a",x"70"),
   241 => (x"4b",x"26",x"86",x"c8"),
   242 => (x"4f",x"26",x"4a",x"26"),
   243 => (x"5b",x"5a",x"5e",x"0e"),
   244 => (x"76",x"8e",x"c8",x"0e"),
   245 => (x"79",x"66",x"d4",x"49"),
   246 => (x"d8",x"49",x"a6",x"c4"),
   247 => (x"e0",x"c0",x"79",x"66"),
   248 => (x"4b",x"76",x"4a",x"a6"),
   249 => (x"5e",x"27",x"1e",x"73"),
   250 => (x"1e",x"00",x"00",x"03"),
   251 => (x"e8",x"c0",x"1e",x"72"),
   252 => (x"89",x"27",x"1e",x"66"),
   253 => (x"0f",x"00",x"00",x"01"),
   254 => (x"4a",x"70",x"86",x"d0"),
   255 => (x"86",x"c8",x"48",x"72"),
   256 => (x"4a",x"26",x"4b",x"26"),
   257 => (x"72",x"1e",x"4f",x"26"),
   258 => (x"76",x"8e",x"c8",x"1e"),
   259 => (x"79",x"66",x"d0",x"49"),
   260 => (x"ff",x"49",x"a6",x"c4"),
   261 => (x"72",x"4a",x"76",x"79"),
   262 => (x"03",x"5e",x"27",x"1e"),
   263 => (x"c0",x"1e",x"00",x"00"),
   264 => (x"c0",x"1e",x"66",x"e0"),
   265 => (x"27",x"1e",x"66",x"e0"),
   266 => (x"00",x"00",x"01",x"89"),
   267 => (x"70",x"86",x"d0",x"0f"),
   268 => (x"c8",x"48",x"72",x"4a"),
   269 => (x"26",x"4a",x"26",x"86"),
   270 => (x"5a",x"5e",x"0e",x"4f"),
   271 => (x"66",x"d0",x"0e",x"5b"),
   272 => (x"7b",x"66",x"cc",x"4b"),
   273 => (x"27",x"1e",x"66",x"cc"),
   274 => (x"00",x"00",x"06",x"68"),
   275 => (x"70",x"86",x"c4",x"0f"),
   276 => (x"05",x"9a",x"72",x"4a"),
   277 => (x"c3",x"87",x"c2",x"c0"),
   278 => (x"4a",x"66",x"cc",x"7b"),
   279 => (x"c0",x"49",x"66",x"cc"),
   280 => (x"db",x"c0",x"02",x"a9"),
   281 => (x"02",x"aa",x"c1",x"87"),
   282 => (x"c2",x"87",x"da",x"c0"),
   283 => (x"ed",x"c0",x"02",x"aa"),
   284 => (x"02",x"aa",x"c3",x"87"),
   285 => (x"c4",x"87",x"ee",x"c0"),
   286 => (x"e6",x"c0",x"02",x"aa"),
   287 => (x"87",x"e5",x"c0",x"87"),
   288 => (x"e0",x"c0",x"7b",x"c0"),
   289 => (x"18",x"20",x"27",x"87"),
   290 => (x"49",x"bf",x"00",x"00"),
   291 => (x"a9",x"b7",x"e4",x"c1"),
   292 => (x"87",x"c5",x"c0",x"06"),
   293 => (x"cc",x"c0",x"7b",x"c0"),
   294 => (x"c0",x"7b",x"c3",x"87"),
   295 => (x"7b",x"c1",x"87",x"c7"),
   296 => (x"c2",x"87",x"c2",x"c0"),
   297 => (x"26",x"4b",x"26",x"7b"),
   298 => (x"1e",x"4f",x"26",x"4a"),
   299 => (x"66",x"c8",x"1e",x"72"),
   300 => (x"cc",x"82",x"c2",x"4a"),
   301 => (x"80",x"72",x"48",x"66"),
   302 => (x"70",x"49",x"66",x"d0"),
   303 => (x"26",x"4a",x"26",x"79"),
   304 => (x"5a",x"5e",x"0e",x"4f"),
   305 => (x"0e",x"5d",x"5c",x"5b"),
   306 => (x"66",x"e0",x"c0",x"1e"),
   307 => (x"75",x"85",x"c5",x"4d"),
   308 => (x"d8",x"94",x"c4",x"4c"),
   309 => (x"e4",x"c0",x"84",x"66"),
   310 => (x"4a",x"75",x"7c",x"66"),
   311 => (x"4b",x"72",x"82",x"c1"),
   312 => (x"66",x"d8",x"93",x"c4"),
   313 => (x"75",x"7b",x"6c",x"83"),
   314 => (x"c4",x"83",x"de",x"4b"),
   315 => (x"83",x"66",x"d8",x"93"),
   316 => (x"49",x"76",x"7b",x"75"),
   317 => (x"b7",x"72",x"79",x"75"),
   318 => (x"df",x"c0",x"01",x"ad"),
   319 => (x"75",x"4c",x"6e",x"87"),
   320 => (x"93",x"c8",x"c3",x"4b"),
   321 => (x"74",x"83",x"66",x"dc"),
   322 => (x"73",x"92",x"c4",x"4a"),
   323 => (x"c1",x"7a",x"75",x"82"),
   324 => (x"c1",x"4a",x"75",x"84"),
   325 => (x"ac",x"b7",x"72",x"82"),
   326 => (x"87",x"e3",x"ff",x"06"),
   327 => (x"c8",x"c3",x"4b",x"75"),
   328 => (x"83",x"66",x"dc",x"93"),
   329 => (x"8a",x"c1",x"4a",x"75"),
   330 => (x"82",x"73",x"92",x"c4"),
   331 => (x"80",x"c1",x"48",x"6a"),
   332 => (x"4a",x"75",x"7a",x"70"),
   333 => (x"66",x"d8",x"92",x"c4"),
   334 => (x"75",x"83",x"72",x"4b"),
   335 => (x"c3",x"84",x"d4",x"4c"),
   336 => (x"66",x"dc",x"94",x"c8"),
   337 => (x"6b",x"82",x"74",x"84"),
   338 => (x"18",x"20",x"27",x"7a"),
   339 => (x"c5",x"49",x"00",x"00"),
   340 => (x"4d",x"26",x"26",x"79"),
   341 => (x"4b",x"26",x"4c",x"26"),
   342 => (x"4f",x"26",x"4a",x"26"),
   343 => (x"5b",x"5a",x"5e",x"0e"),
   344 => (x"d0",x"97",x"0e",x"5c"),
   345 => (x"4b",x"74",x"4c",x"66"),
   346 => (x"c0",x"c0",x"c0",x"c1"),
   347 => (x"c0",x"c4",x"93",x"c0"),
   348 => (x"97",x"4b",x"93",x"b7"),
   349 => (x"c1",x"4a",x"66",x"d4"),
   350 => (x"c0",x"c0",x"c0",x"c0"),
   351 => (x"b7",x"c0",x"c4",x"92"),
   352 => (x"b7",x"72",x"4a",x"92"),
   353 => (x"c5",x"c0",x"02",x"ab"),
   354 => (x"c0",x"48",x"c0",x"87"),
   355 => (x"28",x"27",x"87",x"ca"),
   356 => (x"49",x"00",x"00",x"18"),
   357 => (x"48",x"c1",x"51",x"74"),
   358 => (x"4b",x"26",x"4c",x"26"),
   359 => (x"4f",x"26",x"4a",x"26"),
   360 => (x"5b",x"5a",x"5e",x"0e"),
   361 => (x"97",x"1e",x"0e",x"5c"),
   362 => (x"4b",x"c2",x"4c",x"6e"),
   363 => (x"c1",x"4a",x"66",x"d8"),
   364 => (x"97",x"82",x"73",x"82"),
   365 => (x"c0",x"c1",x"4a",x"6a"),
   366 => (x"92",x"c0",x"c0",x"c0"),
   367 => (x"92",x"b7",x"c0",x"c4"),
   368 => (x"d8",x"1e",x"72",x"4a"),
   369 => (x"82",x"73",x"4a",x"66"),
   370 => (x"c1",x"4a",x"6a",x"97"),
   371 => (x"c0",x"c0",x"c0",x"c0"),
   372 => (x"b7",x"c0",x"c4",x"92"),
   373 => (x"1e",x"72",x"4a",x"92"),
   374 => (x"00",x"05",x"5c",x"27"),
   375 => (x"86",x"c8",x"0f",x"00"),
   376 => (x"9a",x"72",x"4a",x"70"),
   377 => (x"87",x"c5",x"c0",x"05"),
   378 => (x"c1",x"4c",x"c1",x"c1"),
   379 => (x"ab",x"b7",x"c2",x"83"),
   380 => (x"87",x"f8",x"fe",x"06"),
   381 => (x"c0",x"c1",x"4a",x"74"),
   382 => (x"92",x"c0",x"c0",x"c0"),
   383 => (x"92",x"b7",x"c0",x"c4"),
   384 => (x"b7",x"d7",x"c1",x"4a"),
   385 => (x"d7",x"c0",x"04",x"aa"),
   386 => (x"c1",x"4a",x"74",x"87"),
   387 => (x"c0",x"c0",x"c0",x"c0"),
   388 => (x"b7",x"c0",x"c4",x"92"),
   389 => (x"da",x"c1",x"4a",x"92"),
   390 => (x"c0",x"03",x"aa",x"b7"),
   391 => (x"4b",x"c7",x"87",x"c2"),
   392 => (x"c0",x"c1",x"4a",x"74"),
   393 => (x"92",x"c0",x"c0",x"c0"),
   394 => (x"92",x"b7",x"c0",x"c4"),
   395 => (x"aa",x"d2",x"c1",x"4a"),
   396 => (x"87",x"c5",x"c0",x"05"),
   397 => (x"e6",x"c0",x"48",x"c1"),
   398 => (x"4a",x"66",x"d4",x"87"),
   399 => (x"27",x"49",x"66",x"d8"),
   400 => (x"00",x"00",x"06",x"df"),
   401 => (x"c0",x"4a",x"70",x"0f"),
   402 => (x"c0",x"06",x"aa",x"b7"),
   403 => (x"48",x"73",x"87",x"cf"),
   404 => (x"24",x"27",x"80",x"c7"),
   405 => (x"58",x"00",x"00",x"18"),
   406 => (x"c2",x"c0",x"48",x"c1"),
   407 => (x"26",x"48",x"c0",x"87"),
   408 => (x"4b",x"26",x"4c",x"26"),
   409 => (x"4f",x"26",x"4a",x"26"),
   410 => (x"49",x"66",x"c4",x"1e"),
   411 => (x"c0",x"05",x"a9",x"c2"),
   412 => (x"48",x"c1",x"87",x"c5"),
   413 => (x"c0",x"87",x"c2",x"c0"),
   414 => (x"1e",x"4f",x"26",x"48"),
   415 => (x"9a",x"72",x"1e",x"73"),
   416 => (x"c0",x"87",x"e7",x"02"),
   417 => (x"72",x"4b",x"c1",x"48"),
   418 => (x"87",x"d1",x"06",x"a9"),
   419 => (x"c9",x"06",x"82",x"72"),
   420 => (x"72",x"83",x"73",x"87"),
   421 => (x"87",x"f4",x"01",x"a9"),
   422 => (x"b2",x"c1",x"87",x"c3"),
   423 => (x"03",x"a9",x"72",x"3a"),
   424 => (x"07",x"80",x"73",x"89"),
   425 => (x"05",x"2b",x"2a",x"c1"),
   426 => (x"4b",x"26",x"87",x"f3"),
   427 => (x"75",x"1e",x"4f",x"26"),
   428 => (x"71",x"4d",x"c4",x"1e"),
   429 => (x"ff",x"04",x"a1",x"b7"),
   430 => (x"c3",x"81",x"c1",x"b9"),
   431 => (x"b7",x"72",x"07",x"bd"),
   432 => (x"ba",x"ff",x"04",x"a2"),
   433 => (x"bd",x"c1",x"82",x"c1"),
   434 => (x"87",x"ef",x"fe",x"07"),
   435 => (x"ff",x"04",x"2d",x"c1"),
   436 => (x"07",x"80",x"c1",x"b8"),
   437 => (x"b9",x"ff",x"04",x"2d"),
   438 => (x"26",x"07",x"81",x"c1"),
   439 => (x"1e",x"4f",x"26",x"4d"),
   440 => (x"48",x"12",x"1e",x"72"),
   441 => (x"87",x"c4",x"02",x"11"),
   442 => (x"87",x"f6",x"02",x"88"),
   443 => (x"4f",x"26",x"4a",x"26"),
   444 => (x"bf",x"c8",x"ff",x"1e"),
   445 => (x"0e",x"4f",x"26",x"48"),
   446 => (x"5c",x"5b",x"5a",x"5e"),
   447 => (x"8e",x"d0",x"0e",x"5d"),
   448 => (x"27",x"4c",x"66",x"c4"),
   449 => (x"00",x"00",x"18",x"1c"),
   450 => (x"40",x"20",x"27",x"49"),
   451 => (x"27",x"79",x"00",x"00"),
   452 => (x"00",x"00",x"18",x"18"),
   453 => (x"40",x"50",x"27",x"49"),
   454 => (x"27",x"79",x"00",x"00"),
   455 => (x"00",x"00",x"40",x"50"),
   456 => (x"40",x"20",x"27",x"49"),
   457 => (x"27",x"79",x"00",x"00"),
   458 => (x"00",x"00",x"40",x"54"),
   459 => (x"27",x"79",x"c0",x"49"),
   460 => (x"00",x"00",x"40",x"58"),
   461 => (x"27",x"79",x"c2",x"49"),
   462 => (x"00",x"00",x"40",x"5c"),
   463 => (x"79",x"e8",x"c0",x"49"),
   464 => (x"00",x"40",x"60",x"27"),
   465 => (x"d6",x"27",x"49",x"00"),
   466 => (x"48",x"00",x"00",x"11"),
   467 => (x"41",x"20",x"1e",x"72"),
   468 => (x"41",x"20",x"41",x"20"),
   469 => (x"41",x"20",x"41",x"20"),
   470 => (x"41",x"20",x"41",x"20"),
   471 => (x"51",x"10",x"51",x"10"),
   472 => (x"4a",x"26",x"51",x"10"),
   473 => (x"00",x"40",x"80",x"27"),
   474 => (x"f5",x"27",x"49",x"00"),
   475 => (x"48",x"00",x"00",x"11"),
   476 => (x"41",x"20",x"1e",x"72"),
   477 => (x"41",x"20",x"41",x"20"),
   478 => (x"41",x"20",x"41",x"20"),
   479 => (x"41",x"20",x"41",x"20"),
   480 => (x"51",x"10",x"51",x"10"),
   481 => (x"4a",x"26",x"51",x"10"),
   482 => (x"00",x"1f",x"54",x"27"),
   483 => (x"79",x"ca",x"49",x"00"),
   484 => (x"00",x"12",x"14",x"27"),
   485 => (x"3b",x"27",x"1e",x"00"),
   486 => (x"0f",x"00",x"00",x"03"),
   487 => (x"16",x"27",x"86",x"c4"),
   488 => (x"1e",x"00",x"00",x"12"),
   489 => (x"00",x"03",x"3b",x"27"),
   490 => (x"86",x"c4",x"0f",x"00"),
   491 => (x"00",x"12",x"46",x"27"),
   492 => (x"3b",x"27",x"1e",x"00"),
   493 => (x"0f",x"00",x"00",x"03"),
   494 => (x"fc",x"27",x"86",x"c4"),
   495 => (x"bf",x"00",x"00",x"17"),
   496 => (x"87",x"df",x"c0",x"02"),
   497 => (x"00",x"10",x"5d",x"27"),
   498 => (x"3b",x"27",x"1e",x"00"),
   499 => (x"0f",x"00",x"00",x"03"),
   500 => (x"89",x"27",x"86",x"c4"),
   501 => (x"1e",x"00",x"00",x"10"),
   502 => (x"00",x"03",x"3b",x"27"),
   503 => (x"86",x"c4",x"0f",x"00"),
   504 => (x"27",x"87",x"dc",x"c0"),
   505 => (x"00",x"00",x"10",x"8b"),
   506 => (x"03",x"3b",x"27",x"1e"),
   507 => (x"c4",x"0f",x"00",x"00"),
   508 => (x"10",x"ba",x"27",x"86"),
   509 => (x"27",x"1e",x"00",x"00"),
   510 => (x"00",x"00",x"03",x"3b"),
   511 => (x"27",x"86",x"c4",x"0f"),
   512 => (x"00",x"00",x"18",x"00"),
   513 => (x"48",x"27",x"1e",x"bf"),
   514 => (x"1e",x"00",x"00",x"12"),
   515 => (x"00",x"03",x"3b",x"27"),
   516 => (x"86",x"c8",x"0f",x"00"),
   517 => (x"00",x"06",x"f0",x"27"),
   518 => (x"0c",x"27",x"0f",x"00"),
   519 => (x"58",x"00",x"00",x"40"),
   520 => (x"00",x"27",x"4d",x"c1"),
   521 => (x"bf",x"00",x"00",x"18"),
   522 => (x"a9",x"b7",x"c0",x"49"),
   523 => (x"87",x"f8",x"c6",x"06"),
   524 => (x"00",x"10",x"37",x"27"),
   525 => (x"f7",x"27",x"0f",x"00"),
   526 => (x"0f",x"00",x"00",x"0f"),
   527 => (x"79",x"c2",x"49",x"76"),
   528 => (x"a0",x"27",x"4c",x"c3"),
   529 => (x"49",x"00",x"00",x"40"),
   530 => (x"00",x"10",x"db",x"27"),
   531 => (x"1e",x"72",x"48",x"00"),
   532 => (x"41",x"20",x"41",x"20"),
   533 => (x"41",x"20",x"41",x"20"),
   534 => (x"41",x"20",x"41",x"20"),
   535 => (x"51",x"10",x"41",x"20"),
   536 => (x"51",x"10",x"51",x"10"),
   537 => (x"a6",x"c8",x"4a",x"26"),
   538 => (x"27",x"79",x"c1",x"49"),
   539 => (x"00",x"00",x"40",x"a0"),
   540 => (x"40",x"80",x"27",x"1e"),
   541 => (x"27",x"1e",x"00",x"00"),
   542 => (x"00",x"00",x"05",x"a0"),
   543 => (x"70",x"86",x"c8",x"0f"),
   544 => (x"05",x"9a",x"72",x"4a"),
   545 => (x"c1",x"87",x"c5",x"c0"),
   546 => (x"87",x"c2",x"c0",x"4a"),
   547 => (x"24",x"27",x"4a",x"c0"),
   548 => (x"49",x"00",x"00",x"18"),
   549 => (x"49",x"6e",x"79",x"72"),
   550 => (x"03",x"a9",x"b7",x"74"),
   551 => (x"6e",x"87",x"ed",x"c0"),
   552 => (x"72",x"92",x"c5",x"4a"),
   553 => (x"d0",x"88",x"74",x"48"),
   554 => (x"a6",x"cc",x"58",x"a6"),
   555 => (x"74",x"1e",x"72",x"4a"),
   556 => (x"1e",x"66",x"c8",x"1e"),
   557 => (x"00",x"04",x"ab",x"27"),
   558 => (x"86",x"cc",x"0f",x"00"),
   559 => (x"80",x"c1",x"48",x"6e"),
   560 => (x"6e",x"58",x"a6",x"c4"),
   561 => (x"a9",x"b7",x"74",x"49"),
   562 => (x"87",x"d3",x"ff",x"04"),
   563 => (x"c4",x"1e",x"66",x"cc"),
   564 => (x"f8",x"27",x"1e",x"66"),
   565 => (x"1e",x"00",x"00",x"18"),
   566 => (x"00",x"18",x"30",x"27"),
   567 => (x"c1",x"27",x"1e",x"00"),
   568 => (x"0f",x"00",x"00",x"04"),
   569 => (x"18",x"27",x"86",x"d0"),
   570 => (x"bf",x"00",x"00",x"18"),
   571 => (x"0e",x"da",x"27",x"1e"),
   572 => (x"c4",x"0f",x"00",x"00"),
   573 => (x"49",x"a6",x"c4",x"86"),
   574 => (x"27",x"51",x"c1",x"c1"),
   575 => (x"00",x"00",x"18",x"29"),
   576 => (x"c1",x"4a",x"bf",x"97"),
   577 => (x"c0",x"c0",x"c0",x"c0"),
   578 => (x"b7",x"c0",x"c4",x"92"),
   579 => (x"c1",x"c1",x"4a",x"92"),
   580 => (x"c2",x"04",x"aa",x"b7"),
   581 => (x"c3",x"c1",x"87",x"d7"),
   582 => (x"66",x"c8",x"97",x"1e"),
   583 => (x"c0",x"c0",x"c1",x"4a"),
   584 => (x"c4",x"92",x"c0",x"c0"),
   585 => (x"4a",x"92",x"b7",x"c0"),
   586 => (x"5c",x"27",x"1e",x"72"),
   587 => (x"0f",x"00",x"00",x"05"),
   588 => (x"4a",x"70",x"86",x"c8"),
   589 => (x"72",x"49",x"66",x"c8"),
   590 => (x"fd",x"c0",x"05",x"a9"),
   591 => (x"4a",x"a6",x"c8",x"87"),
   592 => (x"1e",x"c0",x"1e",x"72"),
   593 => (x"00",x"04",x"39",x"27"),
   594 => (x"86",x"c8",x"0f",x"00"),
   595 => (x"00",x"40",x"a0",x"27"),
   596 => (x"bc",x"27",x"49",x"00"),
   597 => (x"48",x"00",x"00",x"10"),
   598 => (x"41",x"20",x"1e",x"72"),
   599 => (x"41",x"20",x"41",x"20"),
   600 => (x"41",x"20",x"41",x"20"),
   601 => (x"41",x"20",x"41",x"20"),
   602 => (x"51",x"10",x"51",x"10"),
   603 => (x"4a",x"26",x"51",x"10"),
   604 => (x"20",x"27",x"4c",x"75"),
   605 => (x"49",x"00",x"00",x"18"),
   606 => (x"c4",x"97",x"79",x"75"),
   607 => (x"80",x"c1",x"48",x"66"),
   608 => (x"50",x"08",x"a6",x"c4"),
   609 => (x"4b",x"66",x"c4",x"97"),
   610 => (x"c0",x"c0",x"c0",x"c1"),
   611 => (x"c0",x"c4",x"93",x"c0"),
   612 => (x"27",x"4b",x"93",x"b7"),
   613 => (x"00",x"00",x"18",x"29"),
   614 => (x"c1",x"4a",x"bf",x"97"),
   615 => (x"c0",x"c0",x"c0",x"c0"),
   616 => (x"b7",x"c0",x"c4",x"92"),
   617 => (x"b7",x"72",x"4a",x"92"),
   618 => (x"e9",x"fd",x"06",x"ab"),
   619 => (x"74",x"94",x"6e",x"87"),
   620 => (x"d0",x"1e",x"72",x"49"),
   621 => (x"ae",x"27",x"4a",x"66"),
   622 => (x"0f",x"00",x"00",x"06"),
   623 => (x"48",x"70",x"4a",x"26"),
   624 => (x"74",x"58",x"a6",x"c4"),
   625 => (x"8a",x"66",x"cc",x"4a"),
   626 => (x"4c",x"72",x"92",x"c7"),
   627 => (x"4a",x"76",x"8c",x"6e"),
   628 => (x"74",x"27",x"1e",x"72"),
   629 => (x"0f",x"00",x"00",x"0f"),
   630 => (x"85",x"c1",x"86",x"c4"),
   631 => (x"00",x"18",x"00",x"27"),
   632 => (x"ad",x"b7",x"bf",x"00"),
   633 => (x"87",x"c8",x"f9",x"06"),
   634 => (x"00",x"06",x"f0",x"27"),
   635 => (x"10",x"27",x"0f",x"00"),
   636 => (x"58",x"00",x"00",x"40"),
   637 => (x"00",x"12",x"75",x"27"),
   638 => (x"3b",x"27",x"1e",x"00"),
   639 => (x"0f",x"00",x"00",x"03"),
   640 => (x"85",x"27",x"86",x"c4"),
   641 => (x"1e",x"00",x"00",x"12"),
   642 => (x"00",x"03",x"3b",x"27"),
   643 => (x"86",x"c4",x"0f",x"00"),
   644 => (x"00",x"12",x"87",x"27"),
   645 => (x"3b",x"27",x"1e",x"00"),
   646 => (x"0f",x"00",x"00",x"03"),
   647 => (x"bd",x"27",x"86",x"c4"),
   648 => (x"1e",x"00",x"00",x"12"),
   649 => (x"00",x"03",x"3b",x"27"),
   650 => (x"86",x"c4",x"0f",x"00"),
   651 => (x"00",x"18",x"20",x"27"),
   652 => (x"27",x"1e",x"bf",x"00"),
   653 => (x"00",x"00",x"12",x"bf"),
   654 => (x"03",x"3b",x"27",x"1e"),
   655 => (x"c8",x"0f",x"00",x"00"),
   656 => (x"27",x"1e",x"c5",x"86"),
   657 => (x"00",x"00",x"12",x"d8"),
   658 => (x"03",x"3b",x"27",x"1e"),
   659 => (x"c8",x"0f",x"00",x"00"),
   660 => (x"18",x"24",x"27",x"86"),
   661 => (x"1e",x"bf",x"00",x"00"),
   662 => (x"00",x"12",x"f1",x"27"),
   663 => (x"3b",x"27",x"1e",x"00"),
   664 => (x"0f",x"00",x"00",x"03"),
   665 => (x"1e",x"c1",x"86",x"c8"),
   666 => (x"00",x"13",x"0a",x"27"),
   667 => (x"3b",x"27",x"1e",x"00"),
   668 => (x"0f",x"00",x"00",x"03"),
   669 => (x"28",x"27",x"86",x"c8"),
   670 => (x"97",x"00",x"00",x"18"),
   671 => (x"c0",x"c1",x"4a",x"bf"),
   672 => (x"92",x"c0",x"c0",x"c0"),
   673 => (x"92",x"b7",x"c0",x"c4"),
   674 => (x"27",x"1e",x"72",x"4a"),
   675 => (x"00",x"00",x"13",x"23"),
   676 => (x"03",x"3b",x"27",x"1e"),
   677 => (x"c8",x"0f",x"00",x"00"),
   678 => (x"1e",x"c1",x"c1",x"86"),
   679 => (x"00",x"13",x"3c",x"27"),
   680 => (x"3b",x"27",x"1e",x"00"),
   681 => (x"0f",x"00",x"00",x"03"),
   682 => (x"29",x"27",x"86",x"c8"),
   683 => (x"97",x"00",x"00",x"18"),
   684 => (x"c0",x"c1",x"4a",x"bf"),
   685 => (x"92",x"c0",x"c0",x"c0"),
   686 => (x"92",x"b7",x"c0",x"c4"),
   687 => (x"27",x"1e",x"72",x"4a"),
   688 => (x"00",x"00",x"13",x"55"),
   689 => (x"03",x"3b",x"27",x"1e"),
   690 => (x"c8",x"0f",x"00",x"00"),
   691 => (x"1e",x"c2",x"c1",x"86"),
   692 => (x"00",x"13",x"6e",x"27"),
   693 => (x"3b",x"27",x"1e",x"00"),
   694 => (x"0f",x"00",x"00",x"03"),
   695 => (x"50",x"27",x"86",x"c8"),
   696 => (x"bf",x"00",x"00",x"18"),
   697 => (x"13",x"87",x"27",x"1e"),
   698 => (x"27",x"1e",x"00",x"00"),
   699 => (x"00",x"00",x"03",x"3b"),
   700 => (x"c7",x"86",x"c8",x"0f"),
   701 => (x"13",x"a0",x"27",x"1e"),
   702 => (x"27",x"1e",x"00",x"00"),
   703 => (x"00",x"00",x"03",x"3b"),
   704 => (x"27",x"86",x"c8",x"0f"),
   705 => (x"00",x"00",x"1f",x"54"),
   706 => (x"b9",x"27",x"1e",x"bf"),
   707 => (x"1e",x"00",x"00",x"13"),
   708 => (x"00",x"03",x"3b",x"27"),
   709 => (x"86",x"c8",x"0f",x"00"),
   710 => (x"00",x"13",x"d2",x"27"),
   711 => (x"3b",x"27",x"1e",x"00"),
   712 => (x"0f",x"00",x"00",x"03"),
   713 => (x"fc",x"27",x"86",x"c4"),
   714 => (x"1e",x"00",x"00",x"13"),
   715 => (x"00",x"03",x"3b",x"27"),
   716 => (x"86",x"c4",x"0f",x"00"),
   717 => (x"00",x"18",x"18",x"27"),
   718 => (x"1e",x"bf",x"bf",x"00"),
   719 => (x"00",x"14",x"08",x"27"),
   720 => (x"3b",x"27",x"1e",x"00"),
   721 => (x"0f",x"00",x"00",x"03"),
   722 => (x"21",x"27",x"86",x"c8"),
   723 => (x"1e",x"00",x"00",x"14"),
   724 => (x"00",x"03",x"3b",x"27"),
   725 => (x"86",x"c4",x"0f",x"00"),
   726 => (x"00",x"18",x"18",x"27"),
   727 => (x"c4",x"4a",x"bf",x"00"),
   728 => (x"27",x"1e",x"6a",x"82"),
   729 => (x"00",x"00",x"14",x"52"),
   730 => (x"03",x"3b",x"27",x"1e"),
   731 => (x"c8",x"0f",x"00",x"00"),
   732 => (x"27",x"1e",x"c0",x"86"),
   733 => (x"00",x"00",x"14",x"6b"),
   734 => (x"03",x"3b",x"27",x"1e"),
   735 => (x"c8",x"0f",x"00",x"00"),
   736 => (x"18",x"18",x"27",x"86"),
   737 => (x"4a",x"bf",x"00",x"00"),
   738 => (x"1e",x"6a",x"82",x"c8"),
   739 => (x"00",x"14",x"84",x"27"),
   740 => (x"3b",x"27",x"1e",x"00"),
   741 => (x"0f",x"00",x"00",x"03"),
   742 => (x"1e",x"c2",x"86",x"c8"),
   743 => (x"00",x"14",x"9d",x"27"),
   744 => (x"3b",x"27",x"1e",x"00"),
   745 => (x"0f",x"00",x"00",x"03"),
   746 => (x"18",x"27",x"86",x"c8"),
   747 => (x"bf",x"00",x"00",x"18"),
   748 => (x"6a",x"82",x"cc",x"4a"),
   749 => (x"14",x"b6",x"27",x"1e"),
   750 => (x"27",x"1e",x"00",x"00"),
   751 => (x"00",x"00",x"03",x"3b"),
   752 => (x"d1",x"86",x"c8",x"0f"),
   753 => (x"14",x"cf",x"27",x"1e"),
   754 => (x"27",x"1e",x"00",x"00"),
   755 => (x"00",x"00",x"03",x"3b"),
   756 => (x"27",x"86",x"c8",x"0f"),
   757 => (x"00",x"00",x"18",x"18"),
   758 => (x"82",x"d0",x"4a",x"bf"),
   759 => (x"e8",x"27",x"1e",x"72"),
   760 => (x"1e",x"00",x"00",x"14"),
   761 => (x"00",x"03",x"3b",x"27"),
   762 => (x"86",x"c8",x"0f",x"00"),
   763 => (x"00",x"15",x"01",x"27"),
   764 => (x"3b",x"27",x"1e",x"00"),
   765 => (x"0f",x"00",x"00",x"03"),
   766 => (x"36",x"27",x"86",x"c4"),
   767 => (x"1e",x"00",x"00",x"15"),
   768 => (x"00",x"03",x"3b",x"27"),
   769 => (x"86",x"c4",x"0f",x"00"),
   770 => (x"00",x"18",x"1c",x"27"),
   771 => (x"1e",x"bf",x"bf",x"00"),
   772 => (x"00",x"15",x"47",x"27"),
   773 => (x"3b",x"27",x"1e",x"00"),
   774 => (x"0f",x"00",x"00",x"03"),
   775 => (x"60",x"27",x"86",x"c8"),
   776 => (x"1e",x"00",x"00",x"15"),
   777 => (x"00",x"03",x"3b",x"27"),
   778 => (x"86",x"c4",x"0f",x"00"),
   779 => (x"00",x"18",x"1c",x"27"),
   780 => (x"c4",x"4a",x"bf",x"00"),
   781 => (x"27",x"1e",x"6a",x"82"),
   782 => (x"00",x"00",x"15",x"a0"),
   783 => (x"03",x"3b",x"27",x"1e"),
   784 => (x"c8",x"0f",x"00",x"00"),
   785 => (x"27",x"1e",x"c0",x"86"),
   786 => (x"00",x"00",x"15",x"b9"),
   787 => (x"03",x"3b",x"27",x"1e"),
   788 => (x"c8",x"0f",x"00",x"00"),
   789 => (x"18",x"1c",x"27",x"86"),
   790 => (x"4a",x"bf",x"00",x"00"),
   791 => (x"1e",x"6a",x"82",x"c8"),
   792 => (x"00",x"15",x"d2",x"27"),
   793 => (x"3b",x"27",x"1e",x"00"),
   794 => (x"0f",x"00",x"00",x"03"),
   795 => (x"1e",x"c1",x"86",x"c8"),
   796 => (x"00",x"15",x"eb",x"27"),
   797 => (x"3b",x"27",x"1e",x"00"),
   798 => (x"0f",x"00",x"00",x"03"),
   799 => (x"1c",x"27",x"86",x"c8"),
   800 => (x"bf",x"00",x"00",x"18"),
   801 => (x"6a",x"82",x"cc",x"4a"),
   802 => (x"16",x"04",x"27",x"1e"),
   803 => (x"27",x"1e",x"00",x"00"),
   804 => (x"00",x"00",x"03",x"3b"),
   805 => (x"d2",x"86",x"c8",x"0f"),
   806 => (x"16",x"1d",x"27",x"1e"),
   807 => (x"27",x"1e",x"00",x"00"),
   808 => (x"00",x"00",x"03",x"3b"),
   809 => (x"27",x"86",x"c8",x"0f"),
   810 => (x"00",x"00",x"18",x"1c"),
   811 => (x"82",x"d0",x"4a",x"bf"),
   812 => (x"36",x"27",x"1e",x"72"),
   813 => (x"1e",x"00",x"00",x"16"),
   814 => (x"00",x"03",x"3b",x"27"),
   815 => (x"86",x"c8",x"0f",x"00"),
   816 => (x"00",x"16",x"4f",x"27"),
   817 => (x"3b",x"27",x"1e",x"00"),
   818 => (x"0f",x"00",x"00",x"03"),
   819 => (x"1e",x"6e",x"86",x"c4"),
   820 => (x"00",x"16",x"84",x"27"),
   821 => (x"3b",x"27",x"1e",x"00"),
   822 => (x"0f",x"00",x"00",x"03"),
   823 => (x"1e",x"c5",x"86",x"c8"),
   824 => (x"00",x"16",x"9d",x"27"),
   825 => (x"3b",x"27",x"1e",x"00"),
   826 => (x"0f",x"00",x"00",x"03"),
   827 => (x"1e",x"74",x"86",x"c8"),
   828 => (x"00",x"16",x"b6",x"27"),
   829 => (x"3b",x"27",x"1e",x"00"),
   830 => (x"0f",x"00",x"00",x"03"),
   831 => (x"1e",x"cd",x"86",x"c8"),
   832 => (x"00",x"16",x"cf",x"27"),
   833 => (x"3b",x"27",x"1e",x"00"),
   834 => (x"0f",x"00",x"00",x"03"),
   835 => (x"66",x"cc",x"86",x"c8"),
   836 => (x"16",x"e8",x"27",x"1e"),
   837 => (x"27",x"1e",x"00",x"00"),
   838 => (x"00",x"00",x"03",x"3b"),
   839 => (x"c7",x"86",x"c8",x"0f"),
   840 => (x"17",x"01",x"27",x"1e"),
   841 => (x"27",x"1e",x"00",x"00"),
   842 => (x"00",x"00",x"03",x"3b"),
   843 => (x"c8",x"86",x"c8",x"0f"),
   844 => (x"1a",x"27",x"1e",x"66"),
   845 => (x"1e",x"00",x"00",x"17"),
   846 => (x"00",x"03",x"3b",x"27"),
   847 => (x"86",x"c8",x"0f",x"00"),
   848 => (x"33",x"27",x"1e",x"c1"),
   849 => (x"1e",x"00",x"00",x"17"),
   850 => (x"00",x"03",x"3b",x"27"),
   851 => (x"86",x"c8",x"0f",x"00"),
   852 => (x"00",x"40",x"80",x"27"),
   853 => (x"4c",x"27",x"1e",x"00"),
   854 => (x"1e",x"00",x"00",x"17"),
   855 => (x"00",x"03",x"3b",x"27"),
   856 => (x"86",x"c8",x"0f",x"00"),
   857 => (x"00",x"17",x"65",x"27"),
   858 => (x"3b",x"27",x"1e",x"00"),
   859 => (x"0f",x"00",x"00",x"03"),
   860 => (x"a0",x"27",x"86",x"c4"),
   861 => (x"1e",x"00",x"00",x"40"),
   862 => (x"00",x"17",x"9a",x"27"),
   863 => (x"3b",x"27",x"1e",x"00"),
   864 => (x"0f",x"00",x"00",x"03"),
   865 => (x"b3",x"27",x"86",x"c8"),
   866 => (x"1e",x"00",x"00",x"17"),
   867 => (x"00",x"03",x"3b",x"27"),
   868 => (x"86",x"c4",x"0f",x"00"),
   869 => (x"00",x"17",x"e8",x"27"),
   870 => (x"3b",x"27",x"1e",x"00"),
   871 => (x"0f",x"00",x"00",x"03"),
   872 => (x"0c",x"27",x"86",x"c4"),
   873 => (x"bf",x"00",x"00",x"40"),
   874 => (x"40",x"08",x"27",x"4a"),
   875 => (x"8a",x"bf",x"00",x"00"),
   876 => (x"00",x"40",x"10",x"27"),
   877 => (x"79",x"72",x"49",x"00"),
   878 => (x"ea",x"27",x"1e",x"72"),
   879 => (x"1e",x"00",x"00",x"17"),
   880 => (x"00",x"03",x"3b",x"27"),
   881 => (x"86",x"c8",x"0f",x"00"),
   882 => (x"00",x"40",x"10",x"27"),
   883 => (x"c1",x"49",x"bf",x"00"),
   884 => (x"03",x"a9",x"b7",x"f8"),
   885 => (x"27",x"87",x"ea",x"c0"),
   886 => (x"00",x"00",x"10",x"fa"),
   887 => (x"03",x"3b",x"27",x"1e"),
   888 => (x"c4",x"0f",x"00",x"00"),
   889 => (x"11",x"30",x"27",x"86"),
   890 => (x"27",x"1e",x"00",x"00"),
   891 => (x"00",x"00",x"03",x"3b"),
   892 => (x"27",x"86",x"c4",x"0f"),
   893 => (x"00",x"00",x"11",x"50"),
   894 => (x"03",x"3b",x"27",x"1e"),
   895 => (x"c4",x"0f",x"00",x"00"),
   896 => (x"40",x"10",x"27",x"86"),
   897 => (x"4a",x"bf",x"00",x"00"),
   898 => (x"e8",x"cf",x"4b",x"72"),
   899 => (x"72",x"49",x"73",x"93"),
   900 => (x"18",x"00",x"27",x"1e"),
   901 => (x"4a",x"bf",x"00",x"00"),
   902 => (x"00",x"06",x"ae",x"27"),
   903 => (x"4a",x"26",x"0f",x"00"),
   904 => (x"18",x"27",x"48",x"70"),
   905 => (x"58",x"00",x"00",x"40"),
   906 => (x"00",x"18",x"00",x"27"),
   907 => (x"73",x"4b",x"bf",x"00"),
   908 => (x"94",x"e8",x"cf",x"4c"),
   909 => (x"1e",x"72",x"49",x"74"),
   910 => (x"ae",x"27",x"4a",x"72"),
   911 => (x"0f",x"00",x"00",x"06"),
   912 => (x"48",x"70",x"4a",x"26"),
   913 => (x"00",x"40",x"1c",x"27"),
   914 => (x"f9",x"c8",x"58",x"00"),
   915 => (x"72",x"49",x"73",x"93"),
   916 => (x"27",x"4a",x"72",x"1e"),
   917 => (x"00",x"00",x"06",x"ae"),
   918 => (x"70",x"4a",x"26",x"0f"),
   919 => (x"40",x"20",x"27",x"48"),
   920 => (x"27",x"58",x"00",x"00"),
   921 => (x"00",x"00",x"11",x"52"),
   922 => (x"03",x"3b",x"27",x"1e"),
   923 => (x"c4",x"0f",x"00",x"00"),
   924 => (x"40",x"14",x"27",x"86"),
   925 => (x"1e",x"bf",x"00",x"00"),
   926 => (x"00",x"11",x"7f",x"27"),
   927 => (x"3b",x"27",x"1e",x"00"),
   928 => (x"0f",x"00",x"00",x"03"),
   929 => (x"84",x"27",x"86",x"c8"),
   930 => (x"1e",x"00",x"00",x"11"),
   931 => (x"00",x"03",x"3b",x"27"),
   932 => (x"86",x"c4",x"0f",x"00"),
   933 => (x"00",x"40",x"18",x"27"),
   934 => (x"27",x"1e",x"bf",x"00"),
   935 => (x"00",x"00",x"11",x"b1"),
   936 => (x"03",x"3b",x"27",x"1e"),
   937 => (x"c8",x"0f",x"00",x"00"),
   938 => (x"40",x"1c",x"27",x"86"),
   939 => (x"1e",x"bf",x"00",x"00"),
   940 => (x"00",x"11",x"b6",x"27"),
   941 => (x"3b",x"27",x"1e",x"00"),
   942 => (x"0f",x"00",x"00",x"03"),
   943 => (x"d4",x"27",x"86",x"c8"),
   944 => (x"1e",x"00",x"00",x"11"),
   945 => (x"00",x"03",x"3b",x"27"),
   946 => (x"86",x"c4",x"0f",x"00"),
   947 => (x"86",x"d0",x"48",x"c0"),
   948 => (x"4c",x"26",x"4d",x"26"),
   949 => (x"4a",x"26",x"4b",x"26"),
   950 => (x"5e",x"0e",x"4f",x"26"),
   951 => (x"5d",x"5c",x"5b",x"5a"),
   952 => (x"bf",x"66",x"d4",x"0e"),
   953 => (x"27",x"4d",x"72",x"4a"),
   954 => (x"00",x"00",x"18",x"18"),
   955 => (x"1e",x"72",x"48",x"bf"),
   956 => (x"49",x"a2",x"f0",x"c0"),
   957 => (x"a9",x"72",x"42",x"20"),
   958 => (x"26",x"87",x"f9",x"05"),
   959 => (x"4c",x"66",x"d4",x"4a"),
   960 => (x"7c",x"c5",x"84",x"cc"),
   961 => (x"83",x"cc",x"4b",x"72"),
   962 => (x"66",x"d4",x"7b",x"6c"),
   963 => (x"1e",x"72",x"7a",x"bf"),
   964 => (x"00",x"0f",x"bf",x"27"),
   965 => (x"86",x"c4",x"0f",x"00"),
   966 => (x"05",x"6a",x"82",x"c4"),
   967 => (x"75",x"87",x"f4",x"c0"),
   968 => (x"75",x"83",x"c8",x"4b"),
   969 => (x"c6",x"82",x"cc",x"4a"),
   970 => (x"d8",x"1e",x"73",x"7a"),
   971 => (x"83",x"c8",x"4b",x"66"),
   972 => (x"39",x"27",x"1e",x"6b"),
   973 => (x"0f",x"00",x"00",x"04"),
   974 => (x"18",x"27",x"86",x"c8"),
   975 => (x"bf",x"00",x"00",x"18"),
   976 => (x"1e",x"72",x"7d",x"bf"),
   977 => (x"1e",x"6a",x"1e",x"ca"),
   978 => (x"00",x"04",x"ab",x"27"),
   979 => (x"86",x"cc",x"0f",x"00"),
   980 => (x"d4",x"87",x"d7",x"c0"),
   981 => (x"d4",x"4a",x"bf",x"66"),
   982 => (x"72",x"48",x"49",x"66"),
   983 => (x"a1",x"f0",x"c0",x"1e"),
   984 => (x"71",x"41",x"20",x"4a"),
   985 => (x"87",x"f9",x"05",x"aa"),
   986 => (x"4d",x"26",x"4a",x"26"),
   987 => (x"4b",x"26",x"4c",x"26"),
   988 => (x"4f",x"26",x"4a",x"26"),
   989 => (x"5b",x"5a",x"5e",x"0e"),
   990 => (x"1e",x"0e",x"5d",x"5c"),
   991 => (x"66",x"d8",x"4d",x"6e"),
   992 => (x"ca",x"4b",x"6c",x"4c"),
   993 => (x"18",x"28",x"27",x"83"),
   994 => (x"bf",x"97",x"00",x"00"),
   995 => (x"c0",x"c0",x"c1",x"4a"),
   996 => (x"c4",x"92",x"c0",x"c0"),
   997 => (x"4a",x"92",x"b7",x"c0"),
   998 => (x"05",x"aa",x"c1",x"c1"),
   999 => (x"c1",x"87",x"cf",x"c0"),
  1000 => (x"27",x"48",x"73",x"8b"),
  1001 => (x"00",x"00",x"18",x"20"),
  1002 => (x"7c",x"70",x"88",x"bf"),
  1003 => (x"9d",x"75",x"4d",x"c0"),
  1004 => (x"87",x"d1",x"ff",x"05"),
  1005 => (x"26",x"4d",x"26",x"26"),
  1006 => (x"26",x"4b",x"26",x"4c"),
  1007 => (x"1e",x"4f",x"26",x"4a"),
  1008 => (x"18",x"27",x"1e",x"72"),
  1009 => (x"bf",x"00",x"00",x"18"),
  1010 => (x"87",x"cb",x"c0",x"02"),
  1011 => (x"27",x"49",x"66",x"c8"),
  1012 => (x"00",x"00",x"18",x"18"),
  1013 => (x"27",x"79",x"bf",x"bf"),
  1014 => (x"00",x"00",x"18",x"18"),
  1015 => (x"82",x"cc",x"4a",x"bf"),
  1016 => (x"20",x"27",x"1e",x"72"),
  1017 => (x"bf",x"00",x"00",x"18"),
  1018 => (x"27",x"1e",x"ca",x"1e"),
  1019 => (x"00",x"00",x"04",x"ab"),
  1020 => (x"26",x"86",x"cc",x"0f"),
  1021 => (x"1e",x"4f",x"26",x"4a"),
  1022 => (x"28",x"27",x"1e",x"72"),
  1023 => (x"97",x"00",x"00",x"18"),
  1024 => (x"c0",x"c1",x"4a",x"bf"),
  1025 => (x"92",x"c0",x"c0",x"c0"),
  1026 => (x"92",x"b7",x"c0",x"c4"),
  1027 => (x"aa",x"c1",x"c1",x"4a"),
  1028 => (x"87",x"c5",x"c0",x"02"),
  1029 => (x"c2",x"c0",x"4a",x"c0"),
  1030 => (x"27",x"4a",x"c1",x"87"),
  1031 => (x"00",x"00",x"18",x"24"),
  1032 => (x"b0",x"72",x"48",x"bf"),
  1033 => (x"00",x"18",x"28",x"27"),
  1034 => (x"29",x"27",x"58",x"00"),
  1035 => (x"49",x"00",x"00",x"18"),
  1036 => (x"26",x"51",x"c2",x"c1"),
  1037 => (x"1e",x"4f",x"26",x"4a"),
  1038 => (x"00",x"18",x"28",x"27"),
  1039 => (x"c1",x"c1",x"49",x"00"),
  1040 => (x"18",x"24",x"27",x"51"),
  1041 => (x"c0",x"49",x"00",x"00"),
  1042 => (x"00",x"4f",x"26",x"79"),
  1043 => (x"33",x"32",x"31",x"30"),
  1044 => (x"37",x"36",x"35",x"34"),
  1045 => (x"42",x"41",x"39",x"38"),
  1046 => (x"46",x"45",x"44",x"43"),
  1047 => (x"6f",x"72",x"50",x"00"),
  1048 => (x"6d",x"61",x"72",x"67"),
  1049 => (x"6d",x"6f",x"63",x"20"),
  1050 => (x"65",x"6c",x"69",x"70"),
  1051 => (x"69",x"77",x"20",x"64"),
  1052 => (x"27",x"20",x"68",x"74"),
  1053 => (x"69",x"67",x"65",x"72"),
  1054 => (x"72",x"65",x"74",x"73"),
  1055 => (x"74",x"61",x"20",x"27"),
  1056 => (x"62",x"69",x"72",x"74"),
  1057 => (x"0a",x"65",x"74",x"75"),
  1058 => (x"50",x"00",x"0a",x"00"),
  1059 => (x"72",x"67",x"6f",x"72"),
  1060 => (x"63",x"20",x"6d",x"61"),
  1061 => (x"69",x"70",x"6d",x"6f"),
  1062 => (x"20",x"64",x"65",x"6c"),
  1063 => (x"68",x"74",x"69",x"77"),
  1064 => (x"20",x"74",x"75",x"6f"),
  1065 => (x"67",x"65",x"72",x"27"),
  1066 => (x"65",x"74",x"73",x"69"),
  1067 => (x"61",x"20",x"27",x"72"),
  1068 => (x"69",x"72",x"74",x"74"),
  1069 => (x"65",x"74",x"75",x"62"),
  1070 => (x"00",x"0a",x"00",x"0a"),
  1071 => (x"59",x"52",x"48",x"44"),
  1072 => (x"4e",x"4f",x"54",x"53"),
  1073 => (x"52",x"50",x"20",x"45"),
  1074 => (x"41",x"52",x"47",x"4f"),
  1075 => (x"33",x"20",x"2c",x"4d"),
  1076 => (x"20",x"44",x"52",x"27"),
  1077 => (x"49",x"52",x"54",x"53"),
  1078 => (x"44",x"00",x"47",x"4e"),
  1079 => (x"53",x"59",x"52",x"48"),
  1080 => (x"45",x"4e",x"4f",x"54"),
  1081 => (x"4f",x"52",x"50",x"20"),
  1082 => (x"4d",x"41",x"52",x"47"),
  1083 => (x"27",x"32",x"20",x"2c"),
  1084 => (x"53",x"20",x"44",x"4e"),
  1085 => (x"4e",x"49",x"52",x"54"),
  1086 => (x"65",x"4d",x"00",x"47"),
  1087 => (x"72",x"75",x"73",x"61"),
  1088 => (x"74",x"20",x"64",x"65"),
  1089 => (x"20",x"65",x"6d",x"69"),
  1090 => (x"20",x"6f",x"6f",x"74"),
  1091 => (x"6c",x"61",x"6d",x"73"),
  1092 => (x"6f",x"74",x"20",x"6c"),
  1093 => (x"74",x"62",x"6f",x"20"),
  1094 => (x"20",x"6e",x"69",x"61"),
  1095 => (x"6e",x"61",x"65",x"6d"),
  1096 => (x"66",x"67",x"6e",x"69"),
  1097 => (x"72",x"20",x"6c",x"75"),
  1098 => (x"6c",x"75",x"73",x"65"),
  1099 => (x"00",x"0a",x"73",x"74"),
  1100 => (x"61",x"65",x"6c",x"50"),
  1101 => (x"69",x"20",x"65",x"73"),
  1102 => (x"65",x"72",x"63",x"6e"),
  1103 => (x"20",x"65",x"73",x"61"),
  1104 => (x"62",x"6d",x"75",x"6e"),
  1105 => (x"6f",x"20",x"72",x"65"),
  1106 => (x"75",x"72",x"20",x"66"),
  1107 => (x"00",x"0a",x"73",x"6e"),
  1108 => (x"69",x"4d",x"00",x"0a"),
  1109 => (x"73",x"6f",x"72",x"63"),
  1110 => (x"6e",x"6f",x"63",x"65"),
  1111 => (x"66",x"20",x"73",x"64"),
  1112 => (x"6f",x"20",x"72",x"6f"),
  1113 => (x"72",x"20",x"65",x"6e"),
  1114 => (x"74",x"20",x"6e",x"75"),
  1115 => (x"75",x"6f",x"72",x"68"),
  1116 => (x"44",x"20",x"68",x"67"),
  1117 => (x"73",x"79",x"72",x"68"),
  1118 => (x"65",x"6e",x"6f",x"74"),
  1119 => (x"25",x"00",x"20",x"3a"),
  1120 => (x"00",x"0a",x"20",x"64"),
  1121 => (x"79",x"72",x"68",x"44"),
  1122 => (x"6e",x"6f",x"74",x"73"),
  1123 => (x"70",x"20",x"73",x"65"),
  1124 => (x"53",x"20",x"72",x"65"),
  1125 => (x"6e",x"6f",x"63",x"65"),
  1126 => (x"20",x"20",x"3a",x"64"),
  1127 => (x"20",x"20",x"20",x"20"),
  1128 => (x"20",x"20",x"20",x"20"),
  1129 => (x"20",x"20",x"20",x"20"),
  1130 => (x"20",x"20",x"20",x"20"),
  1131 => (x"20",x"20",x"20",x"20"),
  1132 => (x"20",x"64",x"25",x"00"),
  1133 => (x"41",x"56",x"00",x"0a"),
  1134 => (x"49",x"4d",x"20",x"58"),
  1135 => (x"72",x"20",x"53",x"50"),
  1136 => (x"6e",x"69",x"74",x"61"),
  1137 => (x"20",x"2a",x"20",x"67"),
  1138 => (x"30",x"30",x"30",x"31"),
  1139 => (x"25",x"20",x"3d",x"20"),
  1140 => (x"00",x"0a",x"20",x"64"),
  1141 => (x"48",x"44",x"00",x"0a"),
  1142 => (x"54",x"53",x"59",x"52"),
  1143 => (x"20",x"45",x"4e",x"4f"),
  1144 => (x"47",x"4f",x"52",x"50"),
  1145 => (x"2c",x"4d",x"41",x"52"),
  1146 => (x"4d",x"4f",x"53",x"20"),
  1147 => (x"54",x"53",x"20",x"45"),
  1148 => (x"47",x"4e",x"49",x"52"),
  1149 => (x"52",x"48",x"44",x"00"),
  1150 => (x"4f",x"54",x"53",x"59"),
  1151 => (x"50",x"20",x"45",x"4e"),
  1152 => (x"52",x"47",x"4f",x"52"),
  1153 => (x"20",x"2c",x"4d",x"41"),
  1154 => (x"54",x"53",x"27",x"31"),
  1155 => (x"52",x"54",x"53",x"20"),
  1156 => (x"00",x"47",x"4e",x"49"),
  1157 => (x"68",x"44",x"00",x"0a"),
  1158 => (x"74",x"73",x"79",x"72"),
  1159 => (x"20",x"65",x"6e",x"6f"),
  1160 => (x"63",x"6e",x"65",x"42"),
  1161 => (x"72",x"61",x"6d",x"68"),
  1162 => (x"56",x"20",x"2c",x"6b"),
  1163 => (x"69",x"73",x"72",x"65"),
  1164 => (x"32",x"20",x"6e",x"6f"),
  1165 => (x"28",x"20",x"31",x"2e"),
  1166 => (x"67",x"6e",x"61",x"4c"),
  1167 => (x"65",x"67",x"61",x"75"),
  1168 => (x"29",x"43",x"20",x"3a"),
  1169 => (x"00",x"0a",x"00",x"0a"),
  1170 => (x"63",x"65",x"78",x"45"),
  1171 => (x"6f",x"69",x"74",x"75"),
  1172 => (x"74",x"73",x"20",x"6e"),
  1173 => (x"73",x"74",x"72",x"61"),
  1174 => (x"64",x"25",x"20",x"2c"),
  1175 => (x"6e",x"75",x"72",x"20"),
  1176 => (x"68",x"74",x"20",x"73"),
  1177 => (x"67",x"75",x"6f",x"72"),
  1178 => (x"68",x"44",x"20",x"68"),
  1179 => (x"74",x"73",x"79",x"72"),
  1180 => (x"0a",x"65",x"6e",x"6f"),
  1181 => (x"65",x"78",x"45",x"00"),
  1182 => (x"69",x"74",x"75",x"63"),
  1183 => (x"65",x"20",x"6e",x"6f"),
  1184 => (x"0a",x"73",x"64",x"6e"),
  1185 => (x"46",x"00",x"0a",x"00"),
  1186 => (x"6c",x"61",x"6e",x"69"),
  1187 => (x"6c",x"61",x"76",x"20"),
  1188 => (x"20",x"73",x"65",x"75"),
  1189 => (x"74",x"20",x"66",x"6f"),
  1190 => (x"76",x"20",x"65",x"68"),
  1191 => (x"61",x"69",x"72",x"61"),
  1192 => (x"73",x"65",x"6c",x"62"),
  1193 => (x"65",x"73",x"75",x"20"),
  1194 => (x"6e",x"69",x"20",x"64"),
  1195 => (x"65",x"68",x"74",x"20"),
  1196 => (x"6e",x"65",x"62",x"20"),
  1197 => (x"61",x"6d",x"68",x"63"),
  1198 => (x"0a",x"3a",x"6b",x"72"),
  1199 => (x"49",x"00",x"0a",x"00"),
  1200 => (x"47",x"5f",x"74",x"6e"),
  1201 => (x"3a",x"62",x"6f",x"6c"),
  1202 => (x"20",x"20",x"20",x"20"),
  1203 => (x"20",x"20",x"20",x"20"),
  1204 => (x"20",x"20",x"20",x"20"),
  1205 => (x"00",x"0a",x"64",x"25"),
  1206 => (x"20",x"20",x"20",x"20"),
  1207 => (x"20",x"20",x"20",x"20"),
  1208 => (x"75",x"6f",x"68",x"73"),
  1209 => (x"62",x"20",x"64",x"6c"),
  1210 => (x"20",x"20",x"3a",x"65"),
  1211 => (x"0a",x"64",x"25",x"20"),
  1212 => (x"6f",x"6f",x"42",x"00"),
  1213 => (x"6c",x"47",x"5f",x"6c"),
  1214 => (x"20",x"3a",x"62",x"6f"),
  1215 => (x"20",x"20",x"20",x"20"),
  1216 => (x"20",x"20",x"20",x"20"),
  1217 => (x"64",x"25",x"20",x"20"),
  1218 => (x"20",x"20",x"00",x"0a"),
  1219 => (x"20",x"20",x"20",x"20"),
  1220 => (x"68",x"73",x"20",x"20"),
  1221 => (x"64",x"6c",x"75",x"6f"),
  1222 => (x"3a",x"65",x"62",x"20"),
  1223 => (x"25",x"20",x"20",x"20"),
  1224 => (x"43",x"00",x"0a",x"64"),
  1225 => (x"5f",x"31",x"5f",x"68"),
  1226 => (x"62",x"6f",x"6c",x"47"),
  1227 => (x"20",x"20",x"20",x"3a"),
  1228 => (x"20",x"20",x"20",x"20"),
  1229 => (x"20",x"20",x"20",x"20"),
  1230 => (x"00",x"0a",x"63",x"25"),
  1231 => (x"20",x"20",x"20",x"20"),
  1232 => (x"20",x"20",x"20",x"20"),
  1233 => (x"75",x"6f",x"68",x"73"),
  1234 => (x"62",x"20",x"64",x"6c"),
  1235 => (x"20",x"20",x"3a",x"65"),
  1236 => (x"0a",x"63",x"25",x"20"),
  1237 => (x"5f",x"68",x"43",x"00"),
  1238 => (x"6c",x"47",x"5f",x"32"),
  1239 => (x"20",x"3a",x"62",x"6f"),
  1240 => (x"20",x"20",x"20",x"20"),
  1241 => (x"20",x"20",x"20",x"20"),
  1242 => (x"63",x"25",x"20",x"20"),
  1243 => (x"20",x"20",x"00",x"0a"),
  1244 => (x"20",x"20",x"20",x"20"),
  1245 => (x"68",x"73",x"20",x"20"),
  1246 => (x"64",x"6c",x"75",x"6f"),
  1247 => (x"3a",x"65",x"62",x"20"),
  1248 => (x"25",x"20",x"20",x"20"),
  1249 => (x"41",x"00",x"0a",x"63"),
  1250 => (x"31",x"5f",x"72",x"72"),
  1251 => (x"6f",x"6c",x"47",x"5f"),
  1252 => (x"5d",x"38",x"5b",x"62"),
  1253 => (x"20",x"20",x"20",x"3a"),
  1254 => (x"20",x"20",x"20",x"20"),
  1255 => (x"00",x"0a",x"64",x"25"),
  1256 => (x"20",x"20",x"20",x"20"),
  1257 => (x"20",x"20",x"20",x"20"),
  1258 => (x"75",x"6f",x"68",x"73"),
  1259 => (x"62",x"20",x"64",x"6c"),
  1260 => (x"20",x"20",x"3a",x"65"),
  1261 => (x"0a",x"64",x"25",x"20"),
  1262 => (x"72",x"72",x"41",x"00"),
  1263 => (x"47",x"5f",x"32",x"5f"),
  1264 => (x"5b",x"62",x"6f",x"6c"),
  1265 => (x"37",x"5b",x"5d",x"38"),
  1266 => (x"20",x"20",x"3a",x"5d"),
  1267 => (x"64",x"25",x"20",x"20"),
  1268 => (x"20",x"20",x"00",x"0a"),
  1269 => (x"20",x"20",x"20",x"20"),
  1270 => (x"68",x"73",x"20",x"20"),
  1271 => (x"64",x"6c",x"75",x"6f"),
  1272 => (x"3a",x"65",x"62",x"20"),
  1273 => (x"4e",x"20",x"20",x"20"),
  1274 => (x"65",x"62",x"6d",x"75"),
  1275 => (x"66",x"4f",x"5f",x"72"),
  1276 => (x"6e",x"75",x"52",x"5f"),
  1277 => (x"20",x"2b",x"20",x"73"),
  1278 => (x"00",x"0a",x"30",x"31"),
  1279 => (x"5f",x"72",x"74",x"50"),
  1280 => (x"62",x"6f",x"6c",x"47"),
  1281 => (x"00",x"0a",x"3e",x"2d"),
  1282 => (x"74",x"50",x"20",x"20"),
  1283 => (x"6f",x"43",x"5f",x"72"),
  1284 => (x"20",x"3a",x"70",x"6d"),
  1285 => (x"20",x"20",x"20",x"20"),
  1286 => (x"20",x"20",x"20",x"20"),
  1287 => (x"0a",x"64",x"25",x"20"),
  1288 => (x"20",x"20",x"20",x"00"),
  1289 => (x"20",x"20",x"20",x"20"),
  1290 => (x"6f",x"68",x"73",x"20"),
  1291 => (x"20",x"64",x"6c",x"75"),
  1292 => (x"20",x"3a",x"65",x"62"),
  1293 => (x"69",x"28",x"20",x"20"),
  1294 => (x"65",x"6c",x"70",x"6d"),
  1295 => (x"74",x"6e",x"65",x"6d"),
  1296 => (x"6f",x"69",x"74",x"61"),
  1297 => (x"65",x"64",x"2d",x"6e"),
  1298 => (x"64",x"6e",x"65",x"70"),
  1299 => (x"29",x"74",x"6e",x"65"),
  1300 => (x"20",x"20",x"00",x"0a"),
  1301 => (x"63",x"73",x"69",x"44"),
  1302 => (x"20",x"20",x"3a",x"72"),
  1303 => (x"20",x"20",x"20",x"20"),
  1304 => (x"20",x"20",x"20",x"20"),
  1305 => (x"25",x"20",x"20",x"20"),
  1306 => (x"20",x"00",x"0a",x"64"),
  1307 => (x"20",x"20",x"20",x"20"),
  1308 => (x"73",x"20",x"20",x"20"),
  1309 => (x"6c",x"75",x"6f",x"68"),
  1310 => (x"65",x"62",x"20",x"64"),
  1311 => (x"20",x"20",x"20",x"3a"),
  1312 => (x"00",x"0a",x"64",x"25"),
  1313 => (x"6e",x"45",x"20",x"20"),
  1314 => (x"43",x"5f",x"6d",x"75"),
  1315 => (x"3a",x"70",x"6d",x"6f"),
  1316 => (x"20",x"20",x"20",x"20"),
  1317 => (x"20",x"20",x"20",x"20"),
  1318 => (x"0a",x"64",x"25",x"20"),
  1319 => (x"20",x"20",x"20",x"00"),
  1320 => (x"20",x"20",x"20",x"20"),
  1321 => (x"6f",x"68",x"73",x"20"),
  1322 => (x"20",x"64",x"6c",x"75"),
  1323 => (x"20",x"3a",x"65",x"62"),
  1324 => (x"64",x"25",x"20",x"20"),
  1325 => (x"20",x"20",x"00",x"0a"),
  1326 => (x"5f",x"74",x"6e",x"49"),
  1327 => (x"70",x"6d",x"6f",x"43"),
  1328 => (x"20",x"20",x"20",x"3a"),
  1329 => (x"20",x"20",x"20",x"20"),
  1330 => (x"25",x"20",x"20",x"20"),
  1331 => (x"20",x"00",x"0a",x"64"),
  1332 => (x"20",x"20",x"20",x"20"),
  1333 => (x"73",x"20",x"20",x"20"),
  1334 => (x"6c",x"75",x"6f",x"68"),
  1335 => (x"65",x"62",x"20",x"64"),
  1336 => (x"20",x"20",x"20",x"3a"),
  1337 => (x"00",x"0a",x"64",x"25"),
  1338 => (x"74",x"53",x"20",x"20"),
  1339 => (x"6f",x"43",x"5f",x"72"),
  1340 => (x"20",x"3a",x"70",x"6d"),
  1341 => (x"20",x"20",x"20",x"20"),
  1342 => (x"20",x"20",x"20",x"20"),
  1343 => (x"0a",x"73",x"25",x"20"),
  1344 => (x"20",x"20",x"20",x"00"),
  1345 => (x"20",x"20",x"20",x"20"),
  1346 => (x"6f",x"68",x"73",x"20"),
  1347 => (x"20",x"64",x"6c",x"75"),
  1348 => (x"20",x"3a",x"65",x"62"),
  1349 => (x"48",x"44",x"20",x"20"),
  1350 => (x"54",x"53",x"59",x"52"),
  1351 => (x"20",x"45",x"4e",x"4f"),
  1352 => (x"47",x"4f",x"52",x"50"),
  1353 => (x"2c",x"4d",x"41",x"52"),
  1354 => (x"4d",x"4f",x"53",x"20"),
  1355 => (x"54",x"53",x"20",x"45"),
  1356 => (x"47",x"4e",x"49",x"52"),
  1357 => (x"65",x"4e",x"00",x"0a"),
  1358 => (x"50",x"5f",x"74",x"78"),
  1359 => (x"47",x"5f",x"72",x"74"),
  1360 => (x"2d",x"62",x"6f",x"6c"),
  1361 => (x"20",x"00",x"0a",x"3e"),
  1362 => (x"72",x"74",x"50",x"20"),
  1363 => (x"6d",x"6f",x"43",x"5f"),
  1364 => (x"20",x"20",x"3a",x"70"),
  1365 => (x"20",x"20",x"20",x"20"),
  1366 => (x"20",x"20",x"20",x"20"),
  1367 => (x"00",x"0a",x"64",x"25"),
  1368 => (x"20",x"20",x"20",x"20"),
  1369 => (x"20",x"20",x"20",x"20"),
  1370 => (x"75",x"6f",x"68",x"73"),
  1371 => (x"62",x"20",x"64",x"6c"),
  1372 => (x"20",x"20",x"3a",x"65"),
  1373 => (x"6d",x"69",x"28",x"20"),
  1374 => (x"6d",x"65",x"6c",x"70"),
  1375 => (x"61",x"74",x"6e",x"65"),
  1376 => (x"6e",x"6f",x"69",x"74"),
  1377 => (x"70",x"65",x"64",x"2d"),
  1378 => (x"65",x"64",x"6e",x"65"),
  1379 => (x"2c",x"29",x"74",x"6e"),
  1380 => (x"6d",x"61",x"73",x"20"),
  1381 => (x"73",x"61",x"20",x"65"),
  1382 => (x"6f",x"62",x"61",x"20"),
  1383 => (x"00",x"0a",x"65",x"76"),
  1384 => (x"69",x"44",x"20",x"20"),
  1385 => (x"3a",x"72",x"63",x"73"),
  1386 => (x"20",x"20",x"20",x"20"),
  1387 => (x"20",x"20",x"20",x"20"),
  1388 => (x"20",x"20",x"20",x"20"),
  1389 => (x"0a",x"64",x"25",x"20"),
  1390 => (x"20",x"20",x"20",x"00"),
  1391 => (x"20",x"20",x"20",x"20"),
  1392 => (x"6f",x"68",x"73",x"20"),
  1393 => (x"20",x"64",x"6c",x"75"),
  1394 => (x"20",x"3a",x"65",x"62"),
  1395 => (x"64",x"25",x"20",x"20"),
  1396 => (x"20",x"20",x"00",x"0a"),
  1397 => (x"6d",x"75",x"6e",x"45"),
  1398 => (x"6d",x"6f",x"43",x"5f"),
  1399 => (x"20",x"20",x"3a",x"70"),
  1400 => (x"20",x"20",x"20",x"20"),
  1401 => (x"25",x"20",x"20",x"20"),
  1402 => (x"20",x"00",x"0a",x"64"),
  1403 => (x"20",x"20",x"20",x"20"),
  1404 => (x"73",x"20",x"20",x"20"),
  1405 => (x"6c",x"75",x"6f",x"68"),
  1406 => (x"65",x"62",x"20",x"64"),
  1407 => (x"20",x"20",x"20",x"3a"),
  1408 => (x"00",x"0a",x"64",x"25"),
  1409 => (x"6e",x"49",x"20",x"20"),
  1410 => (x"6f",x"43",x"5f",x"74"),
  1411 => (x"20",x"3a",x"70",x"6d"),
  1412 => (x"20",x"20",x"20",x"20"),
  1413 => (x"20",x"20",x"20",x"20"),
  1414 => (x"0a",x"64",x"25",x"20"),
  1415 => (x"20",x"20",x"20",x"00"),
  1416 => (x"20",x"20",x"20",x"20"),
  1417 => (x"6f",x"68",x"73",x"20"),
  1418 => (x"20",x"64",x"6c",x"75"),
  1419 => (x"20",x"3a",x"65",x"62"),
  1420 => (x"64",x"25",x"20",x"20"),
  1421 => (x"20",x"20",x"00",x"0a"),
  1422 => (x"5f",x"72",x"74",x"53"),
  1423 => (x"70",x"6d",x"6f",x"43"),
  1424 => (x"20",x"20",x"20",x"3a"),
  1425 => (x"20",x"20",x"20",x"20"),
  1426 => (x"25",x"20",x"20",x"20"),
  1427 => (x"20",x"00",x"0a",x"73"),
  1428 => (x"20",x"20",x"20",x"20"),
  1429 => (x"73",x"20",x"20",x"20"),
  1430 => (x"6c",x"75",x"6f",x"68"),
  1431 => (x"65",x"62",x"20",x"64"),
  1432 => (x"20",x"20",x"20",x"3a"),
  1433 => (x"59",x"52",x"48",x"44"),
  1434 => (x"4e",x"4f",x"54",x"53"),
  1435 => (x"52",x"50",x"20",x"45"),
  1436 => (x"41",x"52",x"47",x"4f"),
  1437 => (x"53",x"20",x"2c",x"4d"),
  1438 => (x"20",x"45",x"4d",x"4f"),
  1439 => (x"49",x"52",x"54",x"53"),
  1440 => (x"00",x"0a",x"47",x"4e"),
  1441 => (x"5f",x"74",x"6e",x"49"),
  1442 => (x"6f",x"4c",x"5f",x"31"),
  1443 => (x"20",x"20",x"3a",x"63"),
  1444 => (x"20",x"20",x"20",x"20"),
  1445 => (x"20",x"20",x"20",x"20"),
  1446 => (x"0a",x"64",x"25",x"20"),
  1447 => (x"20",x"20",x"20",x"00"),
  1448 => (x"20",x"20",x"20",x"20"),
  1449 => (x"6f",x"68",x"73",x"20"),
  1450 => (x"20",x"64",x"6c",x"75"),
  1451 => (x"20",x"3a",x"65",x"62"),
  1452 => (x"64",x"25",x"20",x"20"),
  1453 => (x"6e",x"49",x"00",x"0a"),
  1454 => (x"5f",x"32",x"5f",x"74"),
  1455 => (x"3a",x"63",x"6f",x"4c"),
  1456 => (x"20",x"20",x"20",x"20"),
  1457 => (x"20",x"20",x"20",x"20"),
  1458 => (x"25",x"20",x"20",x"20"),
  1459 => (x"20",x"00",x"0a",x"64"),
  1460 => (x"20",x"20",x"20",x"20"),
  1461 => (x"73",x"20",x"20",x"20"),
  1462 => (x"6c",x"75",x"6f",x"68"),
  1463 => (x"65",x"62",x"20",x"64"),
  1464 => (x"20",x"20",x"20",x"3a"),
  1465 => (x"00",x"0a",x"64",x"25"),
  1466 => (x"5f",x"74",x"6e",x"49"),
  1467 => (x"6f",x"4c",x"5f",x"33"),
  1468 => (x"20",x"20",x"3a",x"63"),
  1469 => (x"20",x"20",x"20",x"20"),
  1470 => (x"20",x"20",x"20",x"20"),
  1471 => (x"0a",x"64",x"25",x"20"),
  1472 => (x"20",x"20",x"20",x"00"),
  1473 => (x"20",x"20",x"20",x"20"),
  1474 => (x"6f",x"68",x"73",x"20"),
  1475 => (x"20",x"64",x"6c",x"75"),
  1476 => (x"20",x"3a",x"65",x"62"),
  1477 => (x"64",x"25",x"20",x"20"),
  1478 => (x"6e",x"45",x"00",x"0a"),
  1479 => (x"4c",x"5f",x"6d",x"75"),
  1480 => (x"20",x"3a",x"63",x"6f"),
  1481 => (x"20",x"20",x"20",x"20"),
  1482 => (x"20",x"20",x"20",x"20"),
  1483 => (x"25",x"20",x"20",x"20"),
  1484 => (x"20",x"00",x"0a",x"64"),
  1485 => (x"20",x"20",x"20",x"20"),
  1486 => (x"73",x"20",x"20",x"20"),
  1487 => (x"6c",x"75",x"6f",x"68"),
  1488 => (x"65",x"62",x"20",x"64"),
  1489 => (x"20",x"20",x"20",x"3a"),
  1490 => (x"00",x"0a",x"64",x"25"),
  1491 => (x"5f",x"72",x"74",x"53"),
  1492 => (x"6f",x"4c",x"5f",x"31"),
  1493 => (x"20",x"20",x"3a",x"63"),
  1494 => (x"20",x"20",x"20",x"20"),
  1495 => (x"20",x"20",x"20",x"20"),
  1496 => (x"0a",x"73",x"25",x"20"),
  1497 => (x"20",x"20",x"20",x"00"),
  1498 => (x"20",x"20",x"20",x"20"),
  1499 => (x"6f",x"68",x"73",x"20"),
  1500 => (x"20",x"64",x"6c",x"75"),
  1501 => (x"20",x"3a",x"65",x"62"),
  1502 => (x"48",x"44",x"20",x"20"),
  1503 => (x"54",x"53",x"59",x"52"),
  1504 => (x"20",x"45",x"4e",x"4f"),
  1505 => (x"47",x"4f",x"52",x"50"),
  1506 => (x"2c",x"4d",x"41",x"52"),
  1507 => (x"53",x"27",x"31",x"20"),
  1508 => (x"54",x"53",x"20",x"54"),
  1509 => (x"47",x"4e",x"49",x"52"),
  1510 => (x"74",x"53",x"00",x"0a"),
  1511 => (x"5f",x"32",x"5f",x"72"),
  1512 => (x"3a",x"63",x"6f",x"4c"),
  1513 => (x"20",x"20",x"20",x"20"),
  1514 => (x"20",x"20",x"20",x"20"),
  1515 => (x"25",x"20",x"20",x"20"),
  1516 => (x"20",x"00",x"0a",x"73"),
  1517 => (x"20",x"20",x"20",x"20"),
  1518 => (x"73",x"20",x"20",x"20"),
  1519 => (x"6c",x"75",x"6f",x"68"),
  1520 => (x"65",x"62",x"20",x"64"),
  1521 => (x"20",x"20",x"20",x"3a"),
  1522 => (x"59",x"52",x"48",x"44"),
  1523 => (x"4e",x"4f",x"54",x"53"),
  1524 => (x"52",x"50",x"20",x"45"),
  1525 => (x"41",x"52",x"47",x"4f"),
  1526 => (x"32",x"20",x"2c",x"4d"),
  1527 => (x"20",x"44",x"4e",x"27"),
  1528 => (x"49",x"52",x"54",x"53"),
  1529 => (x"00",x"0a",x"47",x"4e"),
  1530 => (x"73",x"55",x"00",x"0a"),
  1531 => (x"74",x"20",x"72",x"65"),
  1532 => (x"3a",x"65",x"6d",x"69"),
  1533 => (x"0a",x"64",x"25",x"20"),
  1534 => (x"00",x"00",x"00",x"00"),
  1535 => (x"00",x"00",x"00",x"00"),
  1536 => (x"00",x"00",x"61",x"a8"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
